* NGSPICE file created from capbank.ext - technology: sky130B

.subckt sky130_fd_pr__res_xhigh_po_0p35_WX6KG8 a_n35_n532# a_n35_100# VSUBS
X0 a_n35_n532# a_n35_100# VSUBS sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
.ends

.subckt rf_nfet_01v8_aM02W1p65L0p15 DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=4.62e+11p pd=3.86e+06u as=9.24e+11p ps=7.72e+06u w=1.65e+06u l=150000u
X1 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_V3VADT c1_n380_n330# m3_n480_n430#
X0 c1_n380_n330# m3_n480_n430# sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
.ends

.subckt cell_unit ON V_bias OUT_P OUT_N GND
Xsky130_fd_pr__res_xhigh_po_0p35_WX6KG8_0 rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN V_bias
+ GND sky130_fd_pr__res_xhigh_po_0p35_WX6KG8
Xsky130_fd_pr__res_xhigh_po_0p35_WX6KG8_1 rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE V_bias
+ GND sky130_fd_pr__res_xhigh_po_0p35_WX6KG8
Xrf_nfet_01v8_aM02W1p65L0p15_0 rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN ON rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
+ GND rf_nfet_01v8_aM02W1p65L0p15
Xsky130_fd_pr__cap_mim_m3_1_V3VADT_0 OUT_P rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN sky130_fd_pr__cap_mim_m3_1_V3VADT
Xsky130_fd_pr__cap_mim_m3_1_V3VADT_1 OUT_N rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE sky130_fd_pr__cap_mim_m3_1_V3VADT
.ends

.subckt inv_1 ON OUT VDD GND
X0 ON OUT VDD VDD sky130_fd_pr__pfet_01v8 ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
X1 ON OUT GND GND sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=150000u
.ends

.subckt capbank OUT_P OUT_N bit0 bit1 bit2 bit3 bit4 bit5 VDD GND
Xcell_unit_29 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_18 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_19 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_0 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_1 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xinv_1_0 bit5 inv_1_0/OUT VDD GND inv_1
Xinv_1_1 bit4 inv_1_1/OUT VDD GND inv_1
Xcell_unit_3 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_2 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xinv_1_2 bit3 inv_1_2/OUT VDD GND inv_1
Xcell_unit_4 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xinv_1_3 bit2 inv_1_3/OUT VDD GND inv_1
Xcell_unit_5 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xinv_1_4 bit1 inv_1_4/OUT VDD GND inv_1
Xcell_unit_6 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xinv_1_5 bit0 inv_1_5/OUT VDD GND inv_1
Xcell_unit_7 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_8 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_9 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_60 bit1 inv_1_4/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_61 bit1 inv_1_4/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_50 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_62 bit0 inv_1_5/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_51 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_40 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_52 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_41 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_30 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_53 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_42 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_31 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_20 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_54 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_43 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_32 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_10 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_21 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_55 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_44 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_33 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_22 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_11 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_56 bit2 inv_1_3/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_45 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_34 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_23 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_12 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_58 bit2 inv_1_3/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_57 bit2 inv_1_3/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_47 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_46 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_36 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_35 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_25 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_24 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_14 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_13 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_59 bit2 inv_1_3/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_48 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_37 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_26 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_15 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_49 bit3 inv_1_2/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_38 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_27 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_16 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_39 bit4 inv_1_1/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_28 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
Xcell_unit_17 bit5 inv_1_0/OUT OUT_P OUT_N GND cell_unit
.ends

