**.subckt buffer_pex VBIAS VDD GND OUT_P OUT_N IN_P IN_N
*.iopin VBIAS
*.iopin VDD
*.iopin GND
*.opin OUT_P
*.opin OUT_N
*.ipin IN_P
*.ipin IN_N
**** begin user architecture code


* NGSPICE file created from buffer_pex.ext - technology: sky130B

.subckt buffer_pex VDD OUT_P OUT_N IN_P IN_N VBIAS GND
X0 GND.t229 GND.t226 GND.t228 GND.t227 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X1 GND GND.t221 GND GND.t222 sky130_fd_pr__nfet_01v8_lvt ad=1.01808e+14p pd=7.6752e+08u as=0p ps=0u
+ w=5.05e+06u l=150000u
X2 GND GND.t216 GND GND.t217 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X3 GND.t45 VBIAS.t8 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t47
+ GND.t44 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X4 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t46 VBIAS.t9 GND.t31
+ GND.t30 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X5 GND GND.t211 GND GND.t212 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X6 GND.t210 GND.t207 GND.t209 GND.t208 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X7 GND.t33 VBIAS.t10 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t45
+ GND.t32 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X8 GND.t206 GND.t203 GND.t205 GND.t204 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X9 GND GND.t198 GND GND.t199 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X10 GND GND.t193 GND GND.t194 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X11 GND.t192 GND.t189 GND.t191 GND.t190 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X12 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t44 VBIAS.t11
+ GND.t35 GND.t34 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X13 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t0 IN_N.t0 OUT_N.t7
+ GND.t6 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X14 GND.t43 VBIAS.t6 VBIAS.t7 GND.t42 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X15 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t43 VBIAS.t12
+ GND.t37 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X16 GND.t39 VBIAS.t13
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t42 GND.t38 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X17 VBIAS.t5 VBIAS.t4 GND.t258 GND.t257 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X18 GND GND.t184 GND GND.t185 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X19 GND GND.t179 GND GND.t180 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X20 GND.t41 VBIAS.t14
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t41 GND.t40 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X21 GND.t178 GND.t175 GND.t177 GND.t176 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X22 OUT_P.t7 IN_P.t0 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t11
+ GND.t230 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X23 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t3 IN_P.t1 OUT_P.t6
+ GND.t9 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X24 GND.t174 GND.t171 GND.t173 GND.t172 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X25 GND.t25 VBIAS.t15
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t40 GND.t24 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X26 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t39 VBIAS.t16
+ GND.t27 GND.t26 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X27 GND.t29 VBIAS.t17
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t38 GND.t28 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X28 OUT_P.t5 IN_P.t2 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t4
+ GND.t10 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X29 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t37 VBIAS.t18
+ GND.t47 GND.t46 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X30 GND.t49 VBIAS.t19
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t36 GND.t48 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X31 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t35 VBIAS.t20
+ GND.t51 GND.t50 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X32 GND.t13 VBIAS.t21
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t34 GND.t12 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X33 GND GND.t166 GND GND.t167 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X34 GND.t15 VBIAS.t22
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t33 GND.t14 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X35 GND GND.t161 GND GND.t162 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X36 OUT_P.t4 IN_P.t3 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t10
+ GND.t58 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X37 GND.t160 GND.t157 GND.t159 GND.t158 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X38 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t32 VBIAS.t23
+ GND.t17 GND.t16 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X39 GND.t19 VBIAS.t24
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t31 GND.t18 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X40 GND GND.t152 GND GND.t153 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X41 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t30 VBIAS.t25
+ GND.t21 GND.t20 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X42 GND.t23 VBIAS.t26
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t29 GND.t22 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X43 GND.t1 VBIAS.t27 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t28
+ GND.t0 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X44 GND.t255 VBIAS.t2 VBIAS.t3 GND.t254 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X45 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t2 IN_P.t4 OUT_P.t3
+ GND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X46 GND GND.t147 GND GND.t148 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X47 GND GND.t142 GND GND.t143 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X48 GND GND.t137 GND GND.t138 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X49 GND GND.t132 GND GND.t133 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X50 OUT_N.t6 IN_N.t1 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t5
+ GND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X51 OUT_P.t2 IN_P.t5 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t9
+ GND.t57 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X52 GND GND.t127 GND GND.t128 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X53 GND.t3 VBIAS.t28 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t27
+ GND.t2 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X54 GND GND.t122 GND GND.t123 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X55 OUT_N.t5 IN_N.t2 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t15
+ GND.t256 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X56 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t12 IN_N.t3 OUT_N.t4
+ GND.t231 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X57 GND GND.t117 GND GND.t118 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X58 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t6 IN_P.t6 OUT_P.t1
+ GND.t52 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X59 GND.t116 GND.t113 GND.t115 GND.t114 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X60 GND.t5 VBIAS.t29 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t26
+ GND.t4 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X61 GND GND.t108 GND GND.t109 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X62 GND GND.t103 GND GND.t104 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X63 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t25 VBIAS.t30
+ GND.t246 GND.t245 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X64 GND.t248 VBIAS.t31
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t24 GND.t247 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X65 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t23 VBIAS.t32
+ GND.t250 GND.t249 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R0 OUT_N VDD sky130_fd_pr__res_generic_po w=3.5e+06u l=3.5e+06u
X66 GND GND.t98 GND GND.t99 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X67 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t22 VBIAS.t33
+ GND.t240 GND.t239 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X68 GND GND.t93 GND GND.t94 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X69 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t13 IN_N.t4 OUT_N.t3
+ GND.t232 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R1 VDD OUT_P sky130_fd_pr__res_generic_po w=3.5e+06u l=3.5e+06u
X70 GND GND.t88 GND GND.t89 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X71 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t21 VBIAS.t34
+ GND.t242 GND.t241 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X72 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t20 VBIAS.t35
+ GND.t244 GND.t243 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X73 GND.t234 VBIAS.t36
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t19 GND.t233 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X74 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t7 IN_P.t7 OUT_P.t0
+ GND.t53 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X75 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t18 VBIAS.t37
+ GND.t236 GND.t235 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X76 VBIAS.t1 VBIAS.t0 GND.t253 GND.t252 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u
+ w=5.05e+06u l=150000u
X77 GND GND.t83 GND GND.t84 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X78 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t1 IN_N.t5 OUT_N.t2
+ GND.t7 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X79 GND GND.t78 GND GND.t79 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X80 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t17 VBIAS.t38
+ GND.t238 GND.t237 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X81 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t16 VBIAS.t39
+ GND.t55 GND.t54 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X82 GND GND.t73 GND GND.t74 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X83 GND.t72 GND.t69 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X84 OUT_N.t1 IN_N.t6 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t14
+ GND.t251 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X85 OUT_N.t0 IN_N.t7 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t8
+ GND.t56 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X86 GND GND.t64 GND GND.t65 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
X87 GND GND.t59 GND GND.t60 sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u
+ l=150000u
C0 IN_N OUT_N 3.36fF
C1 OUT_P VDD 1.41fF
C2 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE VBIAS 25.10fF
C3 IN_P m4_2257_876# 0.00fF
C4 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE IN_N 5.63fF
C5 IN_P OUT_N 0.41fF
C6 OUT_P m4_2257_876# 0.04fF
C7 IN_N VBIAS 0.20fF
C8 OUT_N VDD 0.83fF
C9 OUT_P OUT_N 7.61fF
C10 IN_P buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE 4.53fF
C11 IN_P VBIAS 0.46fF
C12 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE VDD 1.13fF
C13 OUT_N m4_2257_876# 0.21fF
C14 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE OUT_P 17.63fF
C15 IN_P IN_N 6.75fF
C16 OUT_P VBIAS 0.69fF
C17 IN_N VDD 0.31fF
C18 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE m4_2257_876# 0.40fF
C19 OUT_P IN_N 1.50fF
C20 VBIAS m4_2257_876# 0.08fF
C21 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE OUT_N 19.70fF
C22 IN_P VDD 0.11fF
C23 IN_N m4_2257_876# 0.03fF
C24 OUT_N VBIAS 0.59fF
C25 IN_P OUT_P 4.08fF
R2 GND.n14467 GND.t88 846.712
R3 GND.n15309 GND.t152 846.712
R4 GND.n15289 GND.t189 846.712
R5 GND.n14725 GND.t166 846.712
R6 GND.n15742 GND.t78 846.712
R7 GND.n15731 GND.t127 846.712
R8 GND.n15721 GND.t171 846.712
R9 GND.n15755 GND.t142 846.712
R10 GND.n2661 GND.t83 846.712
R11 GND.n4910 GND.t117 846.712
R12 GND.n1938 GND.t175 846.712
R13 GND.n2634 GND.t184 846.712
R14 GND.n7187 GND.t122 846.712
R15 GND.n7176 GND.t147 846.712
R16 GND.n7166 GND.t157 846.712
R17 GND.n6579 GND.t108 846.712
R18 GND.n10893 GND.t59 846.712
R19 GND.n10882 GND.t179 846.712
R20 GND.n12530 GND.t132 846.712
R21 GND.n10721 GND.t69 846.712
R22 GND.n13534 GND.t216 846.712
R23 GND.n13523 GND.t198 846.712
R24 GND.n13513 GND.t64 846.712
R25 GND.n11437 GND.t226 846.712
R26 GND.n6035 GND.t73 846.712
R27 GND.n6044 GND.t103 846.712
R28 GND.n6114 GND.t113 846.712
R29 GND.n6520 GND.t193 846.712
R30 GND.n9267 GND.t98 846.712
R31 GND.n9284 GND.t161 846.712
R32 GND.n9412 GND.t207 846.712
R33 GND.n8699 GND.t221 846.712
R34 GND.n3371 GND.t93 846.712
R35 GND.n3388 GND.t137 846.712
R36 GND.n1922 GND.t203 846.712
R37 GND.n3359 GND.t211 846.712
R38 GND.n14746 GND.t167 638.041
R39 GND.n15116 GND.t190 638.041
R40 GND.n3341 GND.t212 638.041
R41 GND.n4930 GND.t204 638.041
R42 GND.n3141 GND.t185 638.041
R43 GND.n4584 GND.t176 638.041
R44 GND.n10565 GND.t143 638.041
R45 GND.n15713 GND.t172 638.041
R46 GND.n7210 GND.t109 638.041
R47 GND.n7151 GND.t158 638.041
R48 GND.n6170 GND.t194 638.041
R49 GND.n7982 GND.t114 638.041
R50 GND.n13342 GND.t65 638.041
R51 GND.n11153 GND.t227 638.041
R52 GND.n12521 GND.t133 638.041
R53 GND.n13560 GND.t70 638.041
R54 GND.n11810 GND.t6 638.041
R55 GND.n12915 GND.t256 638.041
R56 GND.n12088 GND.t8 638.041
R57 GND.n13188 GND.t230 638.041
R58 GND.n7955 GND.t53 638.041
R59 GND.n12472 GND.t10 638.041
R60 GND.n7683 GND.t232 638.041
R61 GND.n12192 GND.t11 638.041
R62 GND.n5784 GND.t40 638.041
R63 GND.n8935 GND.t26 638.041
R64 GND.n1228 GND.t14 638.041
R65 GND.n9636 GND.t16 638.041
R66 GND.n1165 GND.t38 638.041
R67 GND.n15936 GND.t20 638.041
R68 GND.n882 GND.t44 638.041
R69 GND.n16224 GND.t50 638.041
R70 GND.n1520 GND.t24 638.041
R71 GND.n9924 GND.t46 638.041
R72 GND.n8713 GND.t42 638.041
R73 GND.n10144 GND.t257 638.041
R74 GND.n8414 GND.t222 638.041
R75 GND.n9970 GND.t208 638.041
R76 GND.n5501 GND.t32 638.041
R77 GND.n9223 GND.t34 638.041
R78 GND.n3664 GND.t28 638.041
R79 GND.n4242 GND.t30 638.041
R80 GND.n3946 GND.t18 638.041
R81 GND.n4531 GND.t36 638.041
R82 GND.t167 GND.t89 356.308
R83 GND.t190 GND.t153 356.308
R84 GND.t212 GND.t94 356.308
R85 GND.t204 GND.t138 356.308
R86 GND.t185 GND.t84 356.308
R87 GND.t176 GND.t118 356.308
R88 GND.t143 GND.t79 356.308
R89 GND.t172 GND.t128 356.308
R90 GND.t109 GND.t123 356.308
R91 GND.t158 GND.t148 356.308
R92 GND.t194 GND.t74 356.308
R93 GND.t114 GND.t104 356.308
R94 GND.t65 GND.t199 356.308
R95 GND.t227 GND.t217 356.308
R96 GND.t133 GND.t180 356.308
R97 GND.t70 GND.t60 356.308
R98 GND.t6 GND.t251 356.308
R99 GND.t256 GND.t231 356.308
R100 GND.t8 GND.t58 356.308
R101 GND.t230 GND.t52 356.308
R102 GND.t53 GND.t57 356.308
R103 GND.t10 GND.t9 356.308
R104 GND.t232 GND.t56 356.308
R105 GND.t11 GND.t7 356.308
R106 GND.t40 GND.t54 356.308
R107 GND.t26 GND.t4 356.308
R108 GND.t14 GND.t241 356.308
R109 GND.t16 GND.t0 356.308
R110 GND.t38 GND.t237 356.308
R111 GND.t20 GND.t22 356.308
R112 GND.t44 GND.t239 356.308
R113 GND.t50 GND.t12 356.308
R114 GND.t24 GND.t245 356.308
R115 GND.t46 GND.t48 356.308
R116 GND.t42 GND.t252 356.308
R117 GND.t257 GND.t254 356.308
R118 GND.t222 GND.t99 356.308
R119 GND.t208 GND.t162 356.308
R120 GND.t32 GND.t243 356.308
R121 GND.t34 GND.t2 356.308
R122 GND.t28 GND.t249 356.308
R123 GND.t30 GND.t247 356.308
R124 GND.t18 GND.t235 356.308
R125 GND.t36 GND.t233 356.308
R126 GND.n4163 GND.n4162 352.212
R127 GND.n2812 GND.n2811 257.615
R128 GND.n2734 GND.n2733 257.615
R129 GND.n2749 GND.n2748 251.553
R130 GND.n4068 GND.n4066 247.742
R131 GND.n2677 GND.n2676 197
R132 GND.n3956 GND.n3955 173.537
R133 GND.n4056 GND.n4055 167.905
R134 GND.n4159 GND.n4158 167.905
R135 GND.n8385 GND.n8384 158.196
R136 GND.n4151 GND.n4150 127.906
R137 GND.n11742 GND.n11741 108.689
R138 GND.n14007 GND.n14006 101.484
R139 GND.n15542 GND.n15541 101.484
R140 GND.n2811 GND.n2810 98.5
R141 GND.n12483 GND.n12482 95.515
R142 GND.n10360 GND.n10359 95.515
R143 GND.n9936 GND.n9935 95.515
R144 GND.n2802 GND.n2801 90.923
R145 GND.n4152 GND.n4149 89.545
R146 GND.n5818 GND.n5817 89.545
R147 GND.n1902 GND.n1901 89.545
R148 GND.n3961 GND.n3960 85.271
R149 GND.n4755 GND.n4754 83.575
R150 GND.n5223 GND.n5222 83.575
R151 GND.n3960 GND.n3959 79.947
R152 GND.n12118 GND.n12117 74.724
R153 GND.n12492 GND.n12491 65.666
R154 GND.n10369 GND.n10368 65.666
R155 GND.n821 GND.n820 65.666
R156 GND.n4556 GND.n4555 62.681
R157 GND.n2678 GND.n2677 60.615
R158 GND.n3962 GND.n3958 59.696
R159 GND.n8883 GND.n8882 59.696
R160 GND.n9238 GND.n9237 59.696
R161 GND.n8065 GND.n8064 55.353
R162 GND.n13424 GND.n13423 55.353
R163 GND.n12609 GND.n12608 55.353
R164 GND.n12908 GND.n12907 55.353
R165 GND.n12465 GND.n12464 55.353
R166 GND.n7074 GND.n7073 55.353
R167 GND.n957 GND.n956 55.353
R168 GND.n1400 GND.n1399 55.353
R169 GND.n5576 GND.n5575 55.353
R170 GND.n4317 GND.n4316 55.353
R171 GND.n15636 GND.n15635 55.353
R172 GND.n4659 GND.n4658 55.353
R173 GND.n5005 GND.n5004 55.353
R174 GND.n14821 GND.n14820 55.353
R175 GND.n3259 GND.n3258 54.344
R176 GND.n3916 GND.n3915 54.344
R177 GND.n3747 GND.n3746 54.344
R178 GND.n3059 GND.n3058 54.344
R179 GND.n7066 GND.n7065 54.344
R180 GND.n7075 GND.n7074 54.344
R181 GND.n8066 GND.n8065 54.344
R182 GND.n8057 GND.n8056 54.344
R183 GND.n7631 GND.n7630 54.344
R184 GND.n7926 GND.n7925 54.344
R185 GND.n13416 GND.n13415 54.344
R186 GND.n13425 GND.n13424 54.344
R187 GND.n12618 GND.n12617 54.344
R188 GND.n12610 GND.n12609 54.344
R189 GND.n13136 GND.n13135 54.344
R190 GND.n12909 GND.n12908 54.344
R191 GND.n12912 GND.n12911 54.344
R192 GND.n11781 GND.n11780 54.344
R193 GND.n12466 GND.n12465 54.344
R194 GND.n12469 GND.n12468 54.344
R195 GND.n6251 GND.n6250 54.344
R196 GND.n7616 GND.n7615 54.344
R197 GND.n11232 GND.n11231 54.344
R198 GND.n13639 GND.n13638 54.344
R199 GND.n10483 GND.n10482 54.344
R200 GND.n14830 GND.n14829 54.344
R201 GND.n14822 GND.n14821 54.344
R202 GND.n9101 GND.n9100 54.344
R203 GND.n9802 GND.n9801 54.344
R204 GND.n16102 GND.n16101 54.344
R205 GND.n1135 GND.n1134 54.344
R206 GND.n966 GND.n965 54.344
R207 GND.n958 GND.n957 54.344
R208 GND.n1198 GND.n1197 54.344
R209 GND.n1392 GND.n1391 54.344
R210 GND.n1401 GND.n1400 54.344
R211 GND.n10053 GND.n10052 54.344
R212 GND.n8792 GND.n8791 54.344
R213 GND.n5754 GND.n5753 54.344
R214 GND.n5585 GND.n5584 54.344
R215 GND.n5577 GND.n5576 54.344
R216 GND.n4326 GND.n4325 54.344
R217 GND.n4318 GND.n4317 54.344
R218 GND.n15628 GND.n15627 54.344
R219 GND.n15637 GND.n15636 54.344
R220 GND.n15190 GND.n15189 54.344
R221 GND.n4668 GND.n4667 54.344
R222 GND.n4660 GND.n4659 54.344
R223 GND.n5014 GND.n5013 54.344
R224 GND.n5006 GND.n5005 54.344
R225 GND.n4572 GND.n4571 53.727
R226 GND.n5795 GND.n5794 53.727
R227 GND.n5232 GND.n5231 53.727
R228 GND.n5446 GND.n5445 53.727
R229 GND.n2825 GND.n2824 51.523
R230 GND.n2976 GND.n2975 47.757
R231 GND.n6141 GND.n6140 47.757
R232 GND.n10337 GND.n10336 47.757
R233 GND.n9951 GND.n9950 47.757
R234 GND.n3247 GND.n3246 47.551
R235 GND.n3852 GND.n3851 47.551
R236 GND.n3647 GND.n3646 47.551
R237 GND.n3047 GND.n3046 47.551
R238 GND.n7747 GND.n7746 47.551
R239 GND.n7938 GND.n7937 47.551
R240 GND.n13072 GND.n13071 47.551
R241 GND.n11966 GND.n11965 47.551
R242 GND.n12044 GND.n12043 47.551
R243 GND.n11793 GND.n11792 47.551
R244 GND.n12259 GND.n12258 47.551
R245 GND.n12148 GND.n12147 47.551
R246 GND.n7305 GND.n7304 47.551
R247 GND.n7271 GND.n7270 47.551
R248 GND.n6263 GND.n6262 47.551
R249 GND.n11244 GND.n11243 47.551
R250 GND.n13651 GND.n13650 47.551
R251 GND.n10471 GND.n10470 47.551
R252 GND.n9001 GND.n9000 47.551
R253 GND.n8910 GND.n8909 47.551
R254 GND.n9206 GND.n9205 47.551
R255 GND.n9702 GND.n9701 47.551
R256 GND.n9611 GND.n9610 47.551
R257 GND.n9907 GND.n9906 47.551
R258 GND.n16002 GND.n16001 47.551
R259 GND.n15911 GND.n15910 47.551
R260 GND.n16207 GND.n16206 47.551
R261 GND.n1071 GND.n1070 47.551
R262 GND.n1292 GND.n1291 47.551
R263 GND.n10239 GND.n10238 47.551
R264 GND.n10205 GND.n10204 47.551
R265 GND.n10065 GND.n10064 47.551
R266 GND.n8804 GND.n8803 47.551
R267 GND.n8509 GND.n8508 47.551
R268 GND.n8475 GND.n8474 47.551
R269 GND.n5690 GND.n5689 47.551
R270 GND.n4431 GND.n4430 47.551
R271 GND.n4506 GND.n4505 47.551
R272 GND.n15178 GND.n15177 47.551
R273 GND.n3947 GND.n3913 44.155
R274 GND.n3933 GND.n3932 44.155
R275 GND.n7684 GND.n7628 44.155
R276 GND.n7661 GND.n7657 44.155
R277 GND.n13189 GND.n13133 44.155
R278 GND.n13166 GND.n13162 44.155
R279 GND.n12087 GND.n12083 44.155
R280 GND.n12191 GND.n12187 44.155
R281 GND.n7211 GND.n7209 44.155
R282 GND.n11154 GND.n11152 44.155
R283 GND.n13561 GND.n13559 44.155
R284 GND.n10413 GND.n10412 44.155
R285 GND.n10566 GND.n10564 44.155
R286 GND.n8936 GND.n8898 44.155
R287 GND.n8934 GND.n8933 44.155
R288 GND.n9637 GND.n9599 44.155
R289 GND.n9635 GND.n9634 44.155
R290 GND.n15937 GND.n15899 44.155
R291 GND.n15935 GND.n15934 44.155
R292 GND.n1166 GND.n1132 44.155
R293 GND.n1152 GND.n1151 44.155
R294 GND.n1229 GND.n1195 44.155
R295 GND.n1215 GND.n1214 44.155
R296 GND.n10303 GND.n10302 44.155
R297 GND.n10145 GND.n10143 44.155
R298 GND.n10127 GND.n10126 44.155
R299 GND.n8866 GND.n8865 44.155
R300 GND.n8714 GND.n8712 44.155
R301 GND.n8415 GND.n8413 44.155
R302 GND.n5785 GND.n5751 44.155
R303 GND.n5771 GND.n5770 44.155
R304 GND.n4532 GND.n4494 44.155
R305 GND.n4530 GND.n4529 44.155
R306 GND.n15878 GND.n15877 41.787
R307 GND.n14734 GND.n14733 41.787
R308 GND.n3235 GND.n3234 40.758
R309 GND.n3864 GND.n3863 40.758
R310 GND.n3643 GND.n3642 40.758
R311 GND.n3035 GND.n3034 40.758
R312 GND.n7041 GND.n7040 40.758
R313 GND.n7100 GND.n7099 40.758
R314 GND.n8091 GND.n8090 40.758
R315 GND.n8032 GND.n8031 40.758
R316 GND.n7730 GND.n7729 40.758
R317 GND.n7918 GND.n7917 40.758
R318 GND.n13391 GND.n13390 40.758
R319 GND.n13450 GND.n13449 40.758
R320 GND.n12643 GND.n12642 40.758
R321 GND.n12584 GND.n12583 40.758
R322 GND.n13084 GND.n13083 40.758
R323 GND.n12891 GND.n12890 40.758
R324 GND.n12965 GND.n12964 40.758
R325 GND.n11773 GND.n11772 40.758
R326 GND.n12448 GND.n12447 40.758
R327 GND.n12360 GND.n12359 40.758
R328 GND.n6275 GND.n6274 40.758
R329 GND.n11256 GND.n11255 40.758
R330 GND.n13663 GND.n13662 40.758
R331 GND.n10459 GND.n10458 40.758
R332 GND.n14855 GND.n14854 40.758
R333 GND.n14796 GND.n14795 40.758
R334 GND.n9202 GND.n9201 40.758
R335 GND.n9903 GND.n9902 40.758
R336 GND.n16203 GND.n16202 40.758
R337 GND.n1083 GND.n1082 40.758
R338 GND.n875 GND.n874 40.758
R339 GND.n932 GND.n931 40.758
R340 GND.n1275 GND.n1274 40.758
R341 GND.n1513 GND.n1512 40.758
R342 GND.n1426 GND.n1425 40.758
R343 GND.n10077 GND.n10076 40.758
R344 GND.n8816 GND.n8815 40.758
R345 GND.n5702 GND.n5701 40.758
R346 GND.n5494 GND.n5493 40.758
R347 GND.n5551 GND.n5550 40.758
R348 GND.n4235 GND.n4234 40.758
R349 GND.n4292 GND.n4291 40.758
R350 GND.n15603 GND.n15602 40.758
R351 GND.n15662 GND.n15661 40.758
R352 GND.n15166 GND.n15165 40.758
R353 GND.n4693 GND.n4692 40.758
R354 GND.n4634 GND.n4633 40.758
R355 GND.n5039 GND.n5038 40.758
R356 GND.n4980 GND.n4979 40.758
R357 GND.n3630 GND.n3629 40.459
R358 GND.n3667 GND.n3666 40.459
R359 GND.n2988 GND.n2987 40.459
R360 GND.n7983 GND.n7981 40.459
R361 GND.n7904 GND.n7903 40.459
R362 GND.n12522 GND.n12520 40.459
R363 GND.n12694 GND.n12693 40.459
R364 GND.n13501 GND.n13500 40.459
R365 GND.n13343 GND.n13341 40.459
R366 GND.n12916 GND.n12853 40.459
R367 GND.n12860 GND.n12859 40.459
R368 GND.n11759 GND.n11758 40.459
R369 GND.n11813 GND.n11812 40.459
R370 GND.n12089 GND.n12028 40.459
R371 GND.n12473 GND.n12410 40.459
R372 GND.n12417 GND.n12416 40.459
R373 GND.n12193 GND.n12132 40.459
R374 GND.n7956 GND.n7897 40.459
R375 GND.n7152 GND.n7150 40.459
R376 GND.n6992 GND.n6991 40.459
R377 GND.n8142 GND.n8141 40.459
R378 GND.n6324 GND.n6323 40.459
R379 GND.n7368 GND.n7367 40.459
R380 GND.n6171 GND.n6169 40.459
R381 GND.n13712 GND.n13711 40.459
R382 GND.n11305 GND.n11304 40.459
R383 GND.n14747 GND.n14745 40.459
R384 GND.n9189 GND.n9188 40.459
R385 GND.n9890 GND.n9889 40.459
R386 GND.n16190 GND.n16189 40.459
R387 GND.n16225 GND.n16183 40.459
R388 GND.n883 GND.n838 40.459
R389 GND.n845 GND.n844 40.459
R390 GND.n9925 GND.n9883 40.459
R391 GND.n1521 GND.n1476 40.459
R392 GND.n1483 GND.n1482 40.459
R393 GND.n9973 GND.n9972 40.459
R394 GND.n8572 GND.n8571 40.459
R395 GND.n9224 GND.n9182 40.459
R396 GND.n5502 GND.n5457 40.459
R397 GND.n5464 GND.n5463 40.459
R398 GND.n4243 GND.n4198 40.459
R399 GND.n4205 GND.n4204 40.459
R400 GND.n15714 GND.n15712 40.459
R401 GND.n15119 GND.n15118 40.459
R402 GND.n15554 GND.n15553 40.459
R403 GND.n4585 GND.n4583 40.459
R404 GND.n4931 GND.n4929 40.459
R405 GND.n4744 GND.n4743 40.459
R406 GND.n5090 GND.n5089 40.459
R407 GND.n3142 GND.n3140 40.459
R408 GND.n3189 GND.n3188 40.459
R409 GND.n3342 GND.n3340 40.459
R410 GND.n14906 GND.n14905 40.459
R411 GND.n15272 GND.n15271 40.459
R412 GND.n3330 GND.n3328 37.362
R413 GND.n3937 GND.n3936 37.362
R414 GND.n3681 GND.n3679 37.362
R415 GND.n3130 GND.n3128 37.362
R416 GND.n7006 GND.n7004 37.362
R417 GND.n7140 GND.n7138 37.362
R418 GND.n8131 GND.n8129 37.362
R419 GND.n7997 GND.n7995 37.362
R420 GND.n7668 GND.n7664 37.362
R421 GND.n13356 GND.n13354 37.362
R422 GND.n13490 GND.n13488 37.362
R423 GND.n12683 GND.n12681 37.362
R424 GND.n12549 GND.n12547 37.362
R425 GND.n13173 GND.n13169 37.362
R426 GND.n12867 GND.n12863 37.362
R427 GND.n12930 GND.n12928 37.362
R428 GND.n11826 GND.n11824 37.362
R429 GND.n12424 GND.n12420 37.362
R430 GND.n12400 GND.n12398 37.362
R431 GND.n6185 GND.n6183 37.362
R432 GND.n11166 GND.n11165 37.362
R433 GND.n13573 GND.n13572 37.362
R434 GND.n10553 GND.n10552 37.362
R435 GND.n14895 GND.n14893 37.362
R436 GND.n14761 GND.n14759 37.362
R437 GND.n9172 GND.n9170 37.362
R438 GND.n9873 GND.n9871 37.362
R439 GND.n16173 GND.n16171 37.362
R440 GND.n1156 GND.n1155 37.362
R441 GND.n852 GND.n848 37.362
R442 GND.n897 GND.n895 37.362
R443 GND.n1219 GND.n1218 37.362
R444 GND.n1490 GND.n1486 37.362
R445 GND.n1466 GND.n1464 37.362
R446 GND.n9987 GND.n9985 37.362
R447 GND.n8726 GND.n8725 37.362
R448 GND.n5775 GND.n5774 37.362
R449 GND.n5471 GND.n5467 37.362
R450 GND.n5516 GND.n5514 37.362
R451 GND.n4212 GND.n4208 37.362
R452 GND.n4257 GND.n4255 37.362
R453 GND.n15568 GND.n15566 37.362
R454 GND.n15702 GND.n15700 37.362
R455 GND.n15261 GND.n15259 37.362
R456 GND.n4733 GND.n4731 37.362
R457 GND.n4599 GND.n4597 37.362
R458 GND.n5079 GND.n5077 37.362
R459 GND.n4945 GND.n4943 37.362
R460 GND.n3200 GND.n3199 34.603
R461 GND.n3901 GND.n3900 34.603
R462 GND.n3663 GND.n3662 34.603
R463 GND.n3000 GND.n2999 34.603
R464 GND.n7695 GND.n7694 34.603
R465 GND.n7954 GND.n7953 34.603
R466 GND.n7886 GND.n7885 34.603
R467 GND.n13121 GND.n13120 34.603
R468 GND.n12080 GND.n12075 34.603
R469 GND.n11809 GND.n11808 34.603
R470 GND.n12017 GND.n12016 34.603
R471 GND.n12184 GND.n12179 34.603
R472 GND.n12205 GND.n12204 34.603
R473 GND.n7222 GND.n7221 34.603
R474 GND.n6312 GND.n6311 34.603
R475 GND.n7356 GND.n7355 34.603
R476 GND.n11293 GND.n11292 34.603
R477 GND.n13700 GND.n13699 34.603
R478 GND.n10424 GND.n10423 34.603
R479 GND.n8930 GND.n8928 34.603
R480 GND.n9222 GND.n9221 34.603
R481 GND.n9631 GND.n9629 34.603
R482 GND.n9923 GND.n9922 34.603
R483 GND.n15931 GND.n15929 34.603
R484 GND.n16223 GND.n16222 34.603
R485 GND.n15948 GND.n15947 34.603
R486 GND.n1120 GND.n1119 34.603
R487 GND.n9648 GND.n9647 34.603
R488 GND.n1240 GND.n1239 34.603
R489 GND.n10156 GND.n10155 34.603
R490 GND.n10114 GND.n10113 34.603
R491 GND.n10290 GND.n10289 34.603
R492 GND.n8853 GND.n8852 34.603
R493 GND.n8426 GND.n8425 34.603
R494 GND.n8560 GND.n8559 34.603
R495 GND.n8947 GND.n8946 34.603
R496 GND.n5739 GND.n5738 34.603
R497 GND.n4526 GND.n4524 34.603
R498 GND.n4482 GND.n4481 34.603
R499 GND.n15131 GND.n15130 34.603
R500 GND.n3223 GND.n3222 33.965
R501 GND.n3876 GND.n3875 33.965
R502 GND.n3655 GND.n3654 33.965
R503 GND.n3023 GND.n3022 33.965
R504 GND.n7718 GND.n7717 33.965
R505 GND.n7946 GND.n7945 33.965
R506 GND.n13096 GND.n13095 33.965
R507 GND.n11991 GND.n11990 33.965
R508 GND.n12060 GND.n12059 33.965
R509 GND.n11801 GND.n11800 33.965
R510 GND.n12229 GND.n12228 33.965
R511 GND.n12164 GND.n12163 33.965
R512 GND.n7330 GND.n7329 33.965
R513 GND.n7246 GND.n7245 33.965
R514 GND.n6287 GND.n6286 33.965
R515 GND.n11268 GND.n11267 33.965
R516 GND.n13675 GND.n13674 33.965
R517 GND.n10447 GND.n10446 33.965
R518 GND.n8971 GND.n8970 33.965
R519 GND.n8919 GND.n8918 33.965
R520 GND.n9214 GND.n9213 33.965
R521 GND.n9672 GND.n9671 33.965
R522 GND.n9620 GND.n9619 33.965
R523 GND.n9915 GND.n9914 33.965
R524 GND.n15972 GND.n15971 33.965
R525 GND.n15920 GND.n15919 33.965
R526 GND.n16215 GND.n16214 33.965
R527 GND.n1095 GND.n1094 33.965
R528 GND.n1263 GND.n1262 33.965
R529 GND.n10264 GND.n10263 33.965
R530 GND.n10180 GND.n10179 33.965
R531 GND.n10089 GND.n10088 33.965
R532 GND.n8828 GND.n8827 33.965
R533 GND.n8534 GND.n8533 33.965
R534 GND.n8450 GND.n8449 33.965
R535 GND.n5714 GND.n5713 33.965
R536 GND.n4456 GND.n4455 33.965
R537 GND.n4515 GND.n4514 33.965
R538 GND.n15154 GND.n15153 33.965
R539 GND.n3317 GND.n3316 30.568
R540 GND.n3929 GND.n3928 30.568
R541 GND.n3693 GND.n3692 30.568
R542 GND.n3117 GND.n3116 30.568
R543 GND.n7654 GND.n7650 30.568
R544 GND.n7875 GND.n7873 30.568
R545 GND.n13159 GND.n13155 30.568
R546 GND.n12006 GND.n12004 30.568
R547 GND.n12072 GND.n12068 30.568
R548 GND.n11839 GND.n11837 30.568
R549 GND.n12219 GND.n12217 30.568
R550 GND.n12176 GND.n12172 30.568
R551 GND.n7345 GND.n7343 30.568
R552 GND.n7236 GND.n7234 30.568
R553 GND.n6197 GND.n6196 30.568
R554 GND.n11178 GND.n11177 30.568
R555 GND.n13585 GND.n13584 30.568
R556 GND.n10541 GND.n10540 30.568
R557 GND.n8961 GND.n8959 30.568
R558 GND.n8925 GND.n8924 30.568
R559 GND.n9159 GND.n9158 30.568
R560 GND.n9662 GND.n9660 30.568
R561 GND.n9626 GND.n9625 30.568
R562 GND.n9860 GND.n9859 30.568
R563 GND.n15962 GND.n15960 30.568
R564 GND.n15926 GND.n15925 30.568
R565 GND.n16160 GND.n16159 30.568
R566 GND.n1148 GND.n1147 30.568
R567 GND.n1211 GND.n1210 30.568
R568 GND.n10279 GND.n10277 30.568
R569 GND.n10170 GND.n10168 30.568
R570 GND.n9999 GND.n9998 30.568
R571 GND.n8738 GND.n8737 30.568
R572 GND.n8549 GND.n8547 30.568
R573 GND.n8440 GND.n8438 30.568
R574 GND.n5767 GND.n5766 30.568
R575 GND.n4471 GND.n4469 30.568
R576 GND.n4521 GND.n4520 30.568
R577 GND.n15249 GND.n15247 30.568
R578 GND.n15310 GND.n15309 29.608
R579 GND.n6045 GND.n6044 29.608
R580 GND.n3212 GND.n3211 28.618
R581 GND.n3889 GND.n3888 28.618
R582 GND.n3637 GND.n3636 28.618
R583 GND.n3012 GND.n3011 28.618
R584 GND.n7126 GND.n7125 28.618
R585 GND.n8008 GND.n8007 28.618
R586 GND.n7707 GND.n7706 28.618
R587 GND.n7911 GND.n7910 28.618
R588 GND.n13476 GND.n13475 28.618
R589 GND.n12560 GND.n12559 28.618
R590 GND.n12669 GND.n12668 28.618
R591 GND.n13367 GND.n13366 28.618
R592 GND.n13109 GND.n13108 28.618
R593 GND.n12941 GND.n12940 28.618
R594 GND.n12875 GND.n12874 28.618
R595 GND.n11766 GND.n11765 28.618
R596 GND.n12386 GND.n12385 28.618
R597 GND.n12432 GND.n12431 28.618
R598 GND.n7017 GND.n7016 28.618
R599 GND.n8117 GND.n8116 28.618
R600 GND.n6300 GND.n6299 28.618
R601 GND.n11281 GND.n11280 28.618
R602 GND.n13688 GND.n13687 28.618
R603 GND.n10436 GND.n10435 28.618
R604 GND.n14772 GND.n14771 28.618
R605 GND.n9196 GND.n9195 28.618
R606 GND.n9897 GND.n9896 28.618
R607 GND.n16197 GND.n16196 28.618
R608 GND.n1108 GND.n1107 28.618
R609 GND.n908 GND.n907 28.618
R610 GND.n860 GND.n859 28.618
R611 GND.n1252 GND.n1251 28.618
R612 GND.n1452 GND.n1451 28.618
R613 GND.n1498 GND.n1497 28.618
R614 GND.n10102 GND.n10101 28.618
R615 GND.n8841 GND.n8840 28.618
R616 GND.n5727 GND.n5726 28.618
R617 GND.n5527 GND.n5526 28.618
R618 GND.n5479 GND.n5478 28.618
R619 GND.n4268 GND.n4267 28.618
R620 GND.n4220 GND.n4219 28.618
R621 GND.n15688 GND.n15687 28.618
R622 GND.n15143 GND.n15142 28.618
R623 GND.n15579 GND.n15578 28.618
R624 GND.n4610 GND.n4609 28.618
R625 GND.n4956 GND.n4955 28.618
R626 GND.n4719 GND.n4718 28.618
R627 GND.n5065 GND.n5064 28.618
R628 GND.n14881 GND.n14880 28.618
R629 GND.n3211 GND.n3210 27.172
R630 GND.n3888 GND.n3887 27.172
R631 GND.n3636 GND.n3635 27.172
R632 GND.n3011 GND.n3010 27.172
R633 GND.n7016 GND.n7015 27.172
R634 GND.n7125 GND.n7124 27.172
R635 GND.n8116 GND.n8115 27.172
R636 GND.n8007 GND.n8006 27.172
R637 GND.n7706 GND.n7705 27.172
R638 GND.n7910 GND.n7909 27.172
R639 GND.n13366 GND.n13365 27.172
R640 GND.n13475 GND.n13474 27.172
R641 GND.n12668 GND.n12667 27.172
R642 GND.n12559 GND.n12558 27.172
R643 GND.n13108 GND.n13107 27.172
R644 GND.n12874 GND.n12873 27.172
R645 GND.n12940 GND.n12939 27.172
R646 GND.n11765 GND.n11764 27.172
R647 GND.n12431 GND.n12430 27.172
R648 GND.n12385 GND.n12384 27.172
R649 GND.n6299 GND.n6298 27.172
R650 GND.n11280 GND.n11279 27.172
R651 GND.n13687 GND.n13686 27.172
R652 GND.n10435 GND.n10434 27.172
R653 GND.n14880 GND.n14879 27.172
R654 GND.n14771 GND.n14770 27.172
R655 GND.n9195 GND.n9194 27.172
R656 GND.n9896 GND.n9895 27.172
R657 GND.n16196 GND.n16195 27.172
R658 GND.n1107 GND.n1106 27.172
R659 GND.n859 GND.n858 27.172
R660 GND.n907 GND.n906 27.172
R661 GND.n1251 GND.n1250 27.172
R662 GND.n1497 GND.n1496 27.172
R663 GND.n1451 GND.n1450 27.172
R664 GND.n10101 GND.n10100 27.172
R665 GND.n8840 GND.n8839 27.172
R666 GND.n5726 GND.n5725 27.172
R667 GND.n5478 GND.n5477 27.172
R668 GND.n5526 GND.n5525 27.172
R669 GND.n4219 GND.n4218 27.172
R670 GND.n4267 GND.n4266 27.172
R671 GND.n15578 GND.n15577 27.172
R672 GND.n15687 GND.n15686 27.172
R673 GND.n15142 GND.n15141 27.172
R674 GND.n4718 GND.n4717 27.172
R675 GND.n4609 GND.n4608 27.172
R676 GND.n5064 GND.n5063 27.172
R677 GND.n4955 GND.n4954 27.172
R678 GND.n3268 GND.n3267 25.966
R679 GND.n3920 GND.n3919 25.966
R680 GND.n3740 GND.n3739 25.966
R681 GND.n3068 GND.n3067 25.966
R682 GND.n7635 GND.n7634 25.966
R683 GND.n7930 GND.n7929 25.966
R684 GND.n13140 GND.n13139 25.966
R685 GND.n13139 GND.n13138 25.966
R686 GND.n12031 GND.n12030 25.966
R687 GND.n12035 GND.n12034 25.966
R688 GND.n11785 GND.n11784 25.966
R689 GND.n12036 GND.n12035 25.966
R690 GND.n12030 GND.n12029 25.966
R691 GND.n11784 GND.n11783 25.966
R692 GND.n12135 GND.n12134 25.966
R693 GND.n12139 GND.n12138 25.966
R694 GND.n12140 GND.n12139 25.966
R695 GND.n12134 GND.n12133 25.966
R696 GND.n7634 GND.n7633 25.966
R697 GND.n7929 GND.n7928 25.966
R698 GND.n7293 GND.n7292 25.966
R699 GND.n7283 GND.n7282 25.966
R700 GND.n6244 GND.n6243 25.966
R701 GND.n7284 GND.n7283 25.966
R702 GND.n6243 GND.n6242 25.966
R703 GND.n7292 GND.n7291 25.966
R704 GND.n11225 GND.n11224 25.966
R705 GND.n13632 GND.n13631 25.966
R706 GND.n11224 GND.n11223 25.966
R707 GND.n13631 GND.n13630 25.966
R708 GND.n10492 GND.n10491 25.966
R709 GND.n8901 GND.n8900 25.966
R710 GND.n8905 GND.n8904 25.966
R711 GND.n9110 GND.n9109 25.966
R712 GND.n9602 GND.n9601 25.966
R713 GND.n9606 GND.n9605 25.966
R714 GND.n9811 GND.n9810 25.966
R715 GND.n15902 GND.n15901 25.966
R716 GND.n15906 GND.n15905 25.966
R717 GND.n16111 GND.n16110 25.966
R718 GND.n15907 GND.n15906 25.966
R719 GND.n15901 GND.n15900 25.966
R720 GND.n16110 GND.n16109 25.966
R721 GND.n1139 GND.n1138 25.966
R722 GND.n1138 GND.n1137 25.966
R723 GND.n9607 GND.n9606 25.966
R724 GND.n9601 GND.n9600 25.966
R725 GND.n9810 GND.n9809 25.966
R726 GND.n1202 GND.n1201 25.966
R727 GND.n1201 GND.n1200 25.966
R728 GND.n10227 GND.n10226 25.966
R729 GND.n10217 GND.n10216 25.966
R730 GND.n10046 GND.n10045 25.966
R731 GND.n10218 GND.n10217 25.966
R732 GND.n10226 GND.n10225 25.966
R733 GND.n10045 GND.n10044 25.966
R734 GND.n8785 GND.n8784 25.966
R735 GND.n8497 GND.n8496 25.966
R736 GND.n8487 GND.n8486 25.966
R737 GND.n8784 GND.n8783 25.966
R738 GND.n8488 GND.n8487 25.966
R739 GND.n8496 GND.n8495 25.966
R740 GND.n8906 GND.n8905 25.966
R741 GND.n8900 GND.n8899 25.966
R742 GND.n9109 GND.n9108 25.966
R743 GND.n5758 GND.n5757 25.966
R744 GND.n5757 GND.n5756 25.966
R745 GND.n4497 GND.n4496 25.966
R746 GND.n4501 GND.n4500 25.966
R747 GND.n4502 GND.n4501 25.966
R748 GND.n4496 GND.n4495 25.966
R749 GND.n15199 GND.n15198 25.966
R750 GND.n3067 GND.n3066 25.966
R751 GND.n3267 GND.n3266 25.966
R752 GND.n10491 GND.n10490 25.966
R753 GND.n15198 GND.n15197 25.966
R754 GND.n3739 GND.n3738 25.966
R755 GND.n3919 GND.n3918 25.966
R756 GND.n4541 GND.n4540 23.878
R757 GND.n5435 GND.n5434 23.878
R758 GND.n3305 GND.n3304 23.775
R759 GND.n3941 GND.n3940 23.775
R760 GND.n3705 GND.n3704 23.775
R761 GND.n3105 GND.n3104 23.775
R762 GND.n7031 GND.n7029 23.775
R763 GND.n7115 GND.n7113 23.775
R764 GND.n8106 GND.n8104 23.775
R765 GND.n8022 GND.n8020 23.775
R766 GND.n7675 GND.n7671 23.775
R767 GND.n7862 GND.n7861 23.775
R768 GND.n13381 GND.n13379 23.775
R769 GND.n13465 GND.n13463 23.775
R770 GND.n12658 GND.n12656 23.775
R771 GND.n12574 GND.n12572 23.775
R772 GND.n13180 GND.n13176 23.775
R773 GND.n12883 GND.n12878 23.775
R774 GND.n12955 GND.n12953 23.775
R775 GND.n11851 GND.n11850 23.775
R776 GND.n12440 GND.n12435 23.775
R777 GND.n12375 GND.n12373 23.775
R778 GND.n6209 GND.n6208 23.775
R779 GND.n11190 GND.n11189 23.775
R780 GND.n13597 GND.n13596 23.775
R781 GND.n10529 GND.n10528 23.775
R782 GND.n14870 GND.n14868 23.775
R783 GND.n14786 GND.n14784 23.775
R784 GND.n9147 GND.n9146 23.775
R785 GND.n9848 GND.n9847 23.775
R786 GND.n16148 GND.n16147 23.775
R787 GND.n1160 GND.n1159 23.775
R788 GND.n868 GND.n863 23.775
R789 GND.n922 GND.n920 23.775
R790 GND.n1223 GND.n1222 23.775
R791 GND.n1506 GND.n1501 23.775
R792 GND.n1441 GND.n1439 23.775
R793 GND.n10011 GND.n10010 23.775
R794 GND.n8750 GND.n8749 23.775
R795 GND.n5779 GND.n5778 23.775
R796 GND.n5487 GND.n5482 23.775
R797 GND.n5541 GND.n5539 23.775
R798 GND.n4228 GND.n4223 23.775
R799 GND.n4282 GND.n4280 23.775
R800 GND.n15593 GND.n15591 23.775
R801 GND.n15677 GND.n15675 23.775
R802 GND.n15236 GND.n15235 23.775
R803 GND.n4708 GND.n4706 23.775
R804 GND.n4624 GND.n4622 23.775
R805 GND.n5054 GND.n5052 23.775
R806 GND.n4970 GND.n4968 23.775
R807 GND.n3280 GND.n3279 22.848
R808 GND.n3944 GND.n3943 22.848
R809 GND.n3728 GND.n3727 22.848
R810 GND.n3080 GND.n3079 22.848
R811 GND.n7054 GND.n7053 22.848
R812 GND.n7087 GND.n7086 22.848
R813 GND.n8079 GND.n8078 22.848
R814 GND.n8044 GND.n8043 22.848
R815 GND.n7678 GND.n7677 22.848
R816 GND.n7837 GND.n7836 22.848
R817 GND.n13404 GND.n13403 22.848
R818 GND.n13437 GND.n13436 22.848
R819 GND.n12631 GND.n12630 22.848
R820 GND.n12596 GND.n12595 22.848
R821 GND.n12597 GND.n12596 22.848
R822 GND.n13438 GND.n13437 22.848
R823 GND.n13403 GND.n13402 22.848
R824 GND.n12630 GND.n12629 22.848
R825 GND.n13183 GND.n13182 22.848
R826 GND.n12895 GND.n12894 22.848
R827 GND.n12976 GND.n12975 22.848
R828 GND.n12977 GND.n12976 22.848
R829 GND.n12894 GND.n12893 22.848
R830 GND.n13182 GND.n13181 22.848
R831 GND.n11873 GND.n11872 22.848
R832 GND.n11872 GND.n11871 22.848
R833 GND.n12452 GND.n12451 22.848
R834 GND.n12347 GND.n12346 22.848
R835 GND.n12348 GND.n12347 22.848
R836 GND.n12451 GND.n12450 22.848
R837 GND.n7677 GND.n7676 22.848
R838 GND.n7836 GND.n7835 22.848
R839 GND.n7088 GND.n7087 22.848
R840 GND.n7053 GND.n7052 22.848
R841 GND.n8045 GND.n8044 22.848
R842 GND.n8078 GND.n8077 22.848
R843 GND.n6232 GND.n6231 22.848
R844 GND.n6231 GND.n6230 22.848
R845 GND.n11213 GND.n11212 22.848
R846 GND.n13620 GND.n13619 22.848
R847 GND.n11212 GND.n11211 22.848
R848 GND.n13619 GND.n13618 22.848
R849 GND.n10504 GND.n10503 22.848
R850 GND.n14843 GND.n14842 22.848
R851 GND.n14808 GND.n14807 22.848
R852 GND.n9122 GND.n9121 22.848
R853 GND.n9823 GND.n9822 22.848
R854 GND.n16123 GND.n16122 22.848
R855 GND.n16122 GND.n16121 22.848
R856 GND.n1163 GND.n1162 22.848
R857 GND.n879 GND.n878 22.848
R858 GND.n944 GND.n943 22.848
R859 GND.n945 GND.n944 22.848
R860 GND.n878 GND.n877 22.848
R861 GND.n1162 GND.n1161 22.848
R862 GND.n9822 GND.n9821 22.848
R863 GND.n1226 GND.n1225 22.848
R864 GND.n1517 GND.n1516 22.848
R865 GND.n1413 GND.n1412 22.848
R866 GND.n1414 GND.n1413 22.848
R867 GND.n1516 GND.n1515 22.848
R868 GND.n1225 GND.n1224 22.848
R869 GND.n10034 GND.n10033 22.848
R870 GND.n10033 GND.n10032 22.848
R871 GND.n8773 GND.n8772 22.848
R872 GND.n8772 GND.n8771 22.848
R873 GND.n9121 GND.n9120 22.848
R874 GND.n5782 GND.n5781 22.848
R875 GND.n5498 GND.n5497 22.848
R876 GND.n5563 GND.n5562 22.848
R877 GND.n5564 GND.n5563 22.848
R878 GND.n5497 GND.n5496 22.848
R879 GND.n5781 GND.n5780 22.848
R880 GND.n4239 GND.n4238 22.848
R881 GND.n4304 GND.n4303 22.848
R882 GND.n4305 GND.n4304 22.848
R883 GND.n4238 GND.n4237 22.848
R884 GND.n15616 GND.n15615 22.848
R885 GND.n15649 GND.n15648 22.848
R886 GND.n15211 GND.n15210 22.848
R887 GND.n15650 GND.n15649 22.848
R888 GND.n15615 GND.n15614 22.848
R889 GND.n4681 GND.n4680 22.848
R890 GND.n4646 GND.n4645 22.848
R891 GND.n5027 GND.n5026 22.848
R892 GND.n4992 GND.n4991 22.848
R893 GND.n4647 GND.n4646 22.848
R894 GND.n4993 GND.n4992 22.848
R895 GND.n4680 GND.n4679 22.848
R896 GND.n5026 GND.n5025 22.848
R897 GND.n3079 GND.n3078 22.848
R898 GND.n3279 GND.n3278 22.848
R899 GND.n14809 GND.n14808 22.848
R900 GND.n10503 GND.n10502 22.848
R901 GND.n14842 GND.n14841 22.848
R902 GND.n15210 GND.n15209 22.848
R903 GND.n3727 GND.n3726 22.848
R904 GND.n3943 GND.n3942 22.848
R905 GND.n3224 GND.n3223 22.503
R906 GND.n3877 GND.n3876 22.503
R907 GND.n3656 GND.n3655 22.503
R908 GND.n3024 GND.n3023 22.503
R909 GND.n7719 GND.n7718 22.503
R910 GND.n7947 GND.n7946 22.503
R911 GND.n13097 GND.n13096 22.503
R912 GND.n12065 GND.n12060 22.503
R913 GND.n11802 GND.n11801 22.503
R914 GND.n11992 GND.n11991 22.503
R915 GND.n12169 GND.n12164 22.503
R916 GND.n12230 GND.n12229 22.503
R917 GND.n7247 GND.n7246 22.503
R918 GND.n6288 GND.n6287 22.503
R919 GND.n7331 GND.n7330 22.503
R920 GND.n11269 GND.n11268 22.503
R921 GND.n13676 GND.n13675 22.503
R922 GND.n10448 GND.n10447 22.503
R923 GND.n8921 GND.n8919 22.503
R924 GND.n9215 GND.n9214 22.503
R925 GND.n9622 GND.n9620 22.503
R926 GND.n9916 GND.n9915 22.503
R927 GND.n15922 GND.n15920 22.503
R928 GND.n16216 GND.n16215 22.503
R929 GND.n15973 GND.n15972 22.503
R930 GND.n1096 GND.n1095 22.503
R931 GND.n9673 GND.n9672 22.503
R932 GND.n1264 GND.n1263 22.503
R933 GND.n10181 GND.n10180 22.503
R934 GND.n10090 GND.n10089 22.503
R935 GND.n10265 GND.n10264 22.503
R936 GND.n8829 GND.n8828 22.503
R937 GND.n8451 GND.n8450 22.503
R938 GND.n8535 GND.n8534 22.503
R939 GND.n8972 GND.n8971 22.503
R940 GND.n5715 GND.n5714 22.503
R941 GND.n4517 GND.n4515 22.503
R942 GND.n4457 GND.n4456 22.503
R943 GND.n15155 GND.n15154 22.503
R944 GND.n3199 GND.n3198 20.379
R945 GND.n3900 GND.n3899 20.379
R946 GND.n3662 GND.n3661 20.379
R947 GND.n2999 GND.n2998 20.379
R948 GND.n7694 GND.n7693 20.379
R949 GND.n7953 GND.n7952 20.379
R950 GND.n7885 GND.n7884 20.379
R951 GND.n13120 GND.n13119 20.379
R952 GND.n12016 GND.n12015 20.379
R953 GND.n12075 GND.n12074 20.379
R954 GND.n11808 GND.n11807 20.379
R955 GND.n11824 GND.n11823 20.379
R956 GND.n12204 GND.n12203 20.379
R957 GND.n12179 GND.n12178 20.379
R958 GND.n7355 GND.n7354 20.379
R959 GND.n7221 GND.n7220 20.379
R960 GND.n6311 GND.n6310 20.379
R961 GND.n7590 GND.n7589 20.379
R962 GND.n11292 GND.n11291 20.379
R963 GND.n13699 GND.n13698 20.379
R964 GND.n10423 GND.n10422 20.379
R965 GND.n8946 GND.n8945 20.379
R966 GND.n8928 GND.n8927 20.379
R967 GND.n9221 GND.n9220 20.379
R968 GND.n9647 GND.n9646 20.379
R969 GND.n9629 GND.n9628 20.379
R970 GND.n9922 GND.n9921 20.379
R971 GND.n15947 GND.n15946 20.379
R972 GND.n15929 GND.n15928 20.379
R973 GND.n16222 GND.n16221 20.379
R974 GND.n1119 GND.n1118 20.379
R975 GND.n1239 GND.n1238 20.379
R976 GND.n10289 GND.n10288 20.379
R977 GND.n10155 GND.n10154 20.379
R978 GND.n10113 GND.n10112 20.379
R979 GND.n8852 GND.n8851 20.379
R980 GND.n8559 GND.n8558 20.379
R981 GND.n8425 GND.n8424 20.379
R982 GND.n5738 GND.n5737 20.379
R983 GND.n4481 GND.n4480 20.379
R984 GND.n4524 GND.n4523 20.379
R985 GND.n15130 GND.n15129 20.379
R986 GND.n15259 GND.n15258 20.379
R987 GND.n8386 GND.n8383 19.952
R988 GND.n3292 GND.n3291 19.694
R989 GND.n3924 GND.n3923 19.694
R990 GND.n3716 GND.n3715 19.694
R991 GND.n3092 GND.n3091 19.694
R992 GND.n7643 GND.n7642 19.694
R993 GND.n7849 GND.n7848 19.694
R994 GND.n13148 GND.n13147 19.694
R995 GND.n13147 GND.n13146 19.694
R996 GND.n11979 GND.n11978 19.694
R997 GND.n12052 GND.n12051 19.694
R998 GND.n11862 GND.n11861 19.694
R999 GND.n12053 GND.n12052 19.694
R1000 GND.n11978 GND.n11977 19.694
R1001 GND.n11861 GND.n11860 19.694
R1002 GND.n12242 GND.n12241 19.694
R1003 GND.n12156 GND.n12155 19.694
R1004 GND.n12157 GND.n12156 19.694
R1005 GND.n12241 GND.n12240 19.694
R1006 GND.n7642 GND.n7641 19.694
R1007 GND.n7848 GND.n7847 19.694
R1008 GND.n7318 GND.n7317 19.694
R1009 GND.n7258 GND.n7257 19.694
R1010 GND.n6220 GND.n6219 19.694
R1011 GND.n7259 GND.n7258 19.694
R1012 GND.n6219 GND.n6218 19.694
R1013 GND.n7317 GND.n7316 19.694
R1014 GND.n11201 GND.n11200 19.694
R1015 GND.n13608 GND.n13607 19.694
R1016 GND.n11200 GND.n11199 19.694
R1017 GND.n13607 GND.n13606 19.694
R1018 GND.n10516 GND.n10515 19.694
R1019 GND.n8984 GND.n8983 19.694
R1020 GND.n8914 GND.n8913 19.694
R1021 GND.n9134 GND.n9133 19.694
R1022 GND.n9685 GND.n9684 19.694
R1023 GND.n9615 GND.n9614 19.694
R1024 GND.n9835 GND.n9834 19.694
R1025 GND.n15985 GND.n15984 19.694
R1026 GND.n15915 GND.n15914 19.694
R1027 GND.n16135 GND.n16134 19.694
R1028 GND.n15916 GND.n15915 19.694
R1029 GND.n15984 GND.n15983 19.694
R1030 GND.n16134 GND.n16133 19.694
R1031 GND.n1143 GND.n1142 19.694
R1032 GND.n1142 GND.n1141 19.694
R1033 GND.n9616 GND.n9615 19.694
R1034 GND.n9684 GND.n9683 19.694
R1035 GND.n9834 GND.n9833 19.694
R1036 GND.n1206 GND.n1205 19.694
R1037 GND.n1205 GND.n1204 19.694
R1038 GND.n10252 GND.n10251 19.694
R1039 GND.n10192 GND.n10191 19.694
R1040 GND.n10022 GND.n10021 19.694
R1041 GND.n10193 GND.n10192 19.694
R1042 GND.n10251 GND.n10250 19.694
R1043 GND.n10021 GND.n10020 19.694
R1044 GND.n8761 GND.n8760 19.694
R1045 GND.n8522 GND.n8521 19.694
R1046 GND.n8462 GND.n8461 19.694
R1047 GND.n8760 GND.n8759 19.694
R1048 GND.n8463 GND.n8462 19.694
R1049 GND.n8521 GND.n8520 19.694
R1050 GND.n8915 GND.n8914 19.694
R1051 GND.n8983 GND.n8982 19.694
R1052 GND.n9133 GND.n9132 19.694
R1053 GND.n5762 GND.n5761 19.694
R1054 GND.n5761 GND.n5760 19.694
R1055 GND.n4444 GND.n4443 19.694
R1056 GND.n4510 GND.n4509 19.694
R1057 GND.n4511 GND.n4510 19.694
R1058 GND.n4443 GND.n4442 19.694
R1059 GND.n15223 GND.n15222 19.694
R1060 GND.n3091 GND.n3090 19.694
R1061 GND.n3291 GND.n3290 19.694
R1062 GND.n10515 GND.n10514 19.694
R1063 GND.n15222 GND.n15221 19.694
R1064 GND.n3715 GND.n3714 19.694
R1065 GND.n3923 GND.n3922 19.694
R1066 GND.n7970 GND.n7969 17.909
R1067 GND.n10328 GND.n10327 17.909
R1068 GND.n9960 GND.n9959 17.909
R1069 GND.n3293 GND.n3292 16.982
R1070 GND.n3925 GND.n3924 16.982
R1071 GND.n3717 GND.n3716 16.982
R1072 GND.n3093 GND.n3092 16.982
R1073 GND.n7647 GND.n7643 16.982
R1074 GND.n7850 GND.n7849 16.982
R1075 GND.n13152 GND.n13148 16.982
R1076 GND.n11981 GND.n11979 16.982
R1077 GND.n12057 GND.n12053 16.982
R1078 GND.n11863 GND.n11862 16.982
R1079 GND.n12244 GND.n12242 16.982
R1080 GND.n12161 GND.n12157 16.982
R1081 GND.n7320 GND.n7318 16.982
R1082 GND.n7261 GND.n7259 16.982
R1083 GND.n6221 GND.n6220 16.982
R1084 GND.n11202 GND.n11201 16.982
R1085 GND.n13609 GND.n13608 16.982
R1086 GND.n10517 GND.n10516 16.982
R1087 GND.n8986 GND.n8984 16.982
R1088 GND.n8916 GND.n8915 16.982
R1089 GND.n9135 GND.n9134 16.982
R1090 GND.n9687 GND.n9685 16.982
R1091 GND.n9617 GND.n9616 16.982
R1092 GND.n9836 GND.n9835 16.982
R1093 GND.n15987 GND.n15985 16.982
R1094 GND.n15917 GND.n15916 16.982
R1095 GND.n16136 GND.n16135 16.982
R1096 GND.n1144 GND.n1143 16.982
R1097 GND.n1207 GND.n1206 16.982
R1098 GND.n10254 GND.n10252 16.982
R1099 GND.n10195 GND.n10193 16.982
R1100 GND.n10023 GND.n10022 16.982
R1101 GND.n8762 GND.n8761 16.982
R1102 GND.n8524 GND.n8522 16.982
R1103 GND.n8465 GND.n8463 16.982
R1104 GND.n5763 GND.n5762 16.982
R1105 GND.n4446 GND.n4444 16.982
R1106 GND.n4512 GND.n4511 16.982
R1107 GND.n15224 GND.n15223 16.982
R1108 GND.n3304 GND.n3303 16.504
R1109 GND.n3940 GND.n3939 16.504
R1110 GND.n3704 GND.n3703 16.504
R1111 GND.n3104 GND.n3103 16.504
R1112 GND.n7029 GND.n7028 16.504
R1113 GND.n7112 GND.n7111 16.504
R1114 GND.n8104 GND.n8103 16.504
R1115 GND.n8019 GND.n8018 16.504
R1116 GND.n7671 GND.n7670 16.504
R1117 GND.n7861 GND.n7860 16.504
R1118 GND.n13379 GND.n13378 16.504
R1119 GND.n13462 GND.n13461 16.504
R1120 GND.n12656 GND.n12655 16.504
R1121 GND.n12571 GND.n12570 16.504
R1122 GND.n12572 GND.n12571 16.504
R1123 GND.n13463 GND.n13462 16.504
R1124 GND.n13378 GND.n13377 16.504
R1125 GND.n12655 GND.n12654 16.504
R1126 GND.n13176 GND.n13175 16.504
R1127 GND.n12878 GND.n12877 16.504
R1128 GND.n12952 GND.n12951 16.504
R1129 GND.n12953 GND.n12952 16.504
R1130 GND.n12877 GND.n12876 16.504
R1131 GND.n13175 GND.n13174 16.504
R1132 GND.n11850 GND.n11849 16.504
R1133 GND.n11849 GND.n11848 16.504
R1134 GND.n12435 GND.n12434 16.504
R1135 GND.n12372 GND.n12371 16.504
R1136 GND.n12373 GND.n12372 16.504
R1137 GND.n12434 GND.n12433 16.504
R1138 GND.n7670 GND.n7669 16.504
R1139 GND.n7860 GND.n7859 16.504
R1140 GND.n7113 GND.n7112 16.504
R1141 GND.n7028 GND.n7027 16.504
R1142 GND.n8020 GND.n8019 16.504
R1143 GND.n8103 GND.n8102 16.504
R1144 GND.n6208 GND.n6207 16.504
R1145 GND.n6207 GND.n6206 16.504
R1146 GND.n11189 GND.n11188 16.504
R1147 GND.n13596 GND.n13595 16.504
R1148 GND.n11188 GND.n11187 16.504
R1149 GND.n13595 GND.n13594 16.504
R1150 GND.n10528 GND.n10527 16.504
R1151 GND.n14868 GND.n14867 16.504
R1152 GND.n14783 GND.n14782 16.504
R1153 GND.n9146 GND.n9145 16.504
R1154 GND.n9847 GND.n9846 16.504
R1155 GND.n16147 GND.n16146 16.504
R1156 GND.n16146 GND.n16145 16.504
R1157 GND.n1159 GND.n1158 16.504
R1158 GND.n863 GND.n862 16.504
R1159 GND.n919 GND.n918 16.504
R1160 GND.n920 GND.n919 16.504
R1161 GND.n862 GND.n861 16.504
R1162 GND.n1158 GND.n1157 16.504
R1163 GND.n9846 GND.n9845 16.504
R1164 GND.n1222 GND.n1221 16.504
R1165 GND.n1501 GND.n1500 16.504
R1166 GND.n1438 GND.n1437 16.504
R1167 GND.n1439 GND.n1438 16.504
R1168 GND.n1500 GND.n1499 16.504
R1169 GND.n1221 GND.n1220 16.504
R1170 GND.n10010 GND.n10009 16.504
R1171 GND.n10009 GND.n10008 16.504
R1172 GND.n8749 GND.n8748 16.504
R1173 GND.n8748 GND.n8747 16.504
R1174 GND.n9145 GND.n9144 16.504
R1175 GND.n5778 GND.n5777 16.504
R1176 GND.n5482 GND.n5481 16.504
R1177 GND.n5538 GND.n5537 16.504
R1178 GND.n5539 GND.n5538 16.504
R1179 GND.n5481 GND.n5480 16.504
R1180 GND.n5777 GND.n5776 16.504
R1181 GND.n4223 GND.n4222 16.504
R1182 GND.n4279 GND.n4278 16.504
R1183 GND.n4280 GND.n4279 16.504
R1184 GND.n4222 GND.n4221 16.504
R1185 GND.n15591 GND.n15590 16.504
R1186 GND.n15674 GND.n15673 16.504
R1187 GND.n15235 GND.n15234 16.504
R1188 GND.n15675 GND.n15674 16.504
R1189 GND.n15590 GND.n15589 16.504
R1190 GND.n4706 GND.n4705 16.504
R1191 GND.n4621 GND.n4620 16.504
R1192 GND.n5052 GND.n5051 16.504
R1193 GND.n4967 GND.n4966 16.504
R1194 GND.n4622 GND.n4621 16.504
R1195 GND.n4968 GND.n4967 16.504
R1196 GND.n4705 GND.n4704 16.504
R1197 GND.n5051 GND.n5050 16.504
R1198 GND.n3103 GND.n3102 16.504
R1199 GND.n3303 GND.n3302 16.504
R1200 GND.n14784 GND.n14783 16.504
R1201 GND.n10527 GND.n10526 16.504
R1202 GND.n14867 GND.n14866 16.504
R1203 GND.n15234 GND.n15233 16.504
R1204 GND.n3703 GND.n3702 16.504
R1205 GND.n3939 GND.n3938 16.504
R1206 GND.n3236 GND.n3235 16.252
R1207 GND.n3865 GND.n3864 16.252
R1208 GND.n3644 GND.n3643 16.252
R1209 GND.n3036 GND.n3035 16.252
R1210 GND.n7101 GND.n7100 16.252
R1211 GND.n8033 GND.n8032 16.252
R1212 GND.n7731 GND.n7730 16.252
R1213 GND.n7919 GND.n7918 16.252
R1214 GND.n13451 GND.n13450 16.252
R1215 GND.n12585 GND.n12584 16.252
R1216 GND.n12644 GND.n12643 16.252
R1217 GND.n13392 GND.n13391 16.252
R1218 GND.n13085 GND.n13084 16.252
R1219 GND.n12966 GND.n12965 16.252
R1220 GND.n12892 GND.n12891 16.252
R1221 GND.n11774 GND.n11773 16.252
R1222 GND.n12361 GND.n12360 16.252
R1223 GND.n12449 GND.n12448 16.252
R1224 GND.n7042 GND.n7041 16.252
R1225 GND.n8092 GND.n8091 16.252
R1226 GND.n6276 GND.n6275 16.252
R1227 GND.n11257 GND.n11256 16.252
R1228 GND.n13664 GND.n13663 16.252
R1229 GND.n10460 GND.n10459 16.252
R1230 GND.n14797 GND.n14796 16.252
R1231 GND.n9203 GND.n9202 16.252
R1232 GND.n9904 GND.n9903 16.252
R1233 GND.n16204 GND.n16203 16.252
R1234 GND.n1084 GND.n1083 16.252
R1235 GND.n933 GND.n932 16.252
R1236 GND.n876 GND.n875 16.252
R1237 GND.n1276 GND.n1275 16.252
R1238 GND.n1427 GND.n1426 16.252
R1239 GND.n1514 GND.n1513 16.252
R1240 GND.n10078 GND.n10077 16.252
R1241 GND.n8817 GND.n8816 16.252
R1242 GND.n5703 GND.n5702 16.252
R1243 GND.n5552 GND.n5551 16.252
R1244 GND.n5495 GND.n5494 16.252
R1245 GND.n4293 GND.n4292 16.252
R1246 GND.n4236 GND.n4235 16.252
R1247 GND.n15663 GND.n15662 16.252
R1248 GND.n15167 GND.n15166 16.252
R1249 GND.n15604 GND.n15603 16.252
R1250 GND.n4635 GND.n4634 16.252
R1251 GND.n4981 GND.n4980 16.252
R1252 GND.n4694 GND.n4693 16.252
R1253 GND.n5040 GND.n5039 16.252
R1254 GND.n14856 GND.n14855 16.252
R1255 GND.n14726 GND.n14725 15.887
R1256 GND.n15290 GND.n15289 15.887
R1257 GND.n14918 GND.n14917 15.887
R1258 GND.n15443 GND.n15442 15.887
R1259 GND.n15756 GND.n15755 15.887
R1260 GND.n15722 GND.n15721 15.887
R1261 GND.n10399 GND.n10398 15.887
R1262 GND.n15534 GND.n15533 15.887
R1263 GND.n2635 GND.n2634 15.887
R1264 GND.n1939 GND.n1938 15.887
R1265 GND.n2967 GND.n2966 15.887
R1266 GND.n4765 GND.n4764 15.887
R1267 GND.n6580 GND.n6579 15.887
R1268 GND.n7167 GND.n7166 15.887
R1269 GND.n7422 GND.n7421 15.887
R1270 GND.n6153 GND.n6152 15.887
R1271 GND.n12708 GND.n12707 15.887
R1272 GND.n11003 GND.n11002 15.887
R1273 GND.n12531 GND.n12530 15.887
R1274 GND.n10722 GND.n10721 15.887
R1275 GND.n13325 GND.n13324 15.887
R1276 GND.n11015 GND.n11014 15.887
R1277 GND.n13514 GND.n13513 15.887
R1278 GND.n11438 GND.n11437 15.887
R1279 GND.n8373 GND.n8372 15.887
R1280 GND.n6115 GND.n6114 15.887
R1281 GND.n6521 GND.n6520 15.887
R1282 GND.n8155 GND.n8154 15.887
R1283 GND.n9255 GND.n9254 15.887
R1284 GND.n9413 GND.n9412 15.887
R1285 GND.n8700 GND.n8699 15.887
R1286 GND.n1180 GND.n1179 15.887
R1287 GND.n3360 GND.n3359 15.887
R1288 GND.n1923 GND.n1922 15.887
R1289 GND.n3159 GND.n3158 15.887
R1290 GND.n1931 GND.n1930 15.887
R1291 GND.n3188 GND.n3187 13.586
R1292 GND.n3340 GND.n3339 13.586
R1293 GND.n3629 GND.n3628 13.586
R1294 GND.n3666 GND.n3665 13.586
R1295 GND.n2987 GND.n2986 13.586
R1296 GND.n3140 GND.n3139 13.586
R1297 GND.n6991 GND.n6990 13.586
R1298 GND.n7150 GND.n7149 13.586
R1299 GND.n8141 GND.n8140 13.586
R1300 GND.n7981 GND.n7980 13.586
R1301 GND.n7903 GND.n7902 13.586
R1302 GND.n7897 GND.n7896 13.586
R1303 GND.n13341 GND.n13340 13.586
R1304 GND.n13500 GND.n13499 13.586
R1305 GND.n12693 GND.n12692 13.586
R1306 GND.n12520 GND.n12519 13.586
R1307 GND.n12859 GND.n12858 13.586
R1308 GND.n12853 GND.n12852 13.586
R1309 GND.n12028 GND.n12027 13.586
R1310 GND.n11758 GND.n11757 13.586
R1311 GND.n11812 GND.n11811 13.586
R1312 GND.n12132 GND.n12131 13.586
R1313 GND.n12416 GND.n12415 13.586
R1314 GND.n12410 GND.n12409 13.586
R1315 GND.n7367 GND.n7366 13.586
R1316 GND.n6323 GND.n6322 13.586
R1317 GND.n6169 GND.n6168 13.586
R1318 GND.n13199 GND.n13198 13.586
R1319 GND.n11304 GND.n11303 13.586
R1320 GND.n13711 GND.n13710 13.586
R1321 GND.n14905 GND.n14904 13.586
R1322 GND.n14745 GND.n14744 13.586
R1323 GND.n9188 GND.n9187 13.586
R1324 GND.n9182 GND.n9181 13.586
R1325 GND.n9889 GND.n9888 13.586
R1326 GND.n9883 GND.n9882 13.586
R1327 GND.n16189 GND.n16188 13.586
R1328 GND.n16183 GND.n16182 13.586
R1329 GND.n844 GND.n843 13.586
R1330 GND.n838 GND.n837 13.586
R1331 GND.n1482 GND.n1481 13.586
R1332 GND.n1476 GND.n1475 13.586
R1333 GND.n9972 GND.n9971 13.586
R1334 GND.n8571 GND.n8570 13.586
R1335 GND.n5463 GND.n5462 13.586
R1336 GND.n5457 GND.n5456 13.586
R1337 GND.n4204 GND.n4203 13.586
R1338 GND.n4198 GND.n4197 13.586
R1339 GND.n15553 GND.n15552 13.586
R1340 GND.n15712 GND.n15711 13.586
R1341 GND.n15118 GND.n15117 13.586
R1342 GND.n15271 GND.n15270 13.586
R1343 GND.n4743 GND.n4742 13.586
R1344 GND.n4583 GND.n4582 13.586
R1345 GND.n5089 GND.n5088 13.586
R1346 GND.n4929 GND.n4928 13.586
R1347 GND.n13069 GND.n13068 13.552
R1348 GND.n12983 GND.n12982 13.552
R1349 GND.n11963 GND.n11962 13.552
R1350 GND.n11878 GND.n11877 13.552
R1351 GND.n12256 GND.n12255 13.552
R1352 GND.n12344 GND.n12343 13.552
R1353 GND.n7744 GND.n7743 13.552
R1354 GND.n7833 GND.n7832 13.552
R1355 GND.n15999 GND.n15998 13.552
R1356 GND.n814 GND.n813 13.552
R1357 GND.n16095 GND.n16094 13.552
R1358 GND.n1068 GND.n1067 13.552
R1359 GND.n817 GND.n816 13.552
R1360 GND.n975 GND.n974 13.552
R1361 GND.n9699 GND.n9698 13.552
R1362 GND.n9591 GND.n9590 13.552
R1363 GND.n9795 GND.n9794 13.552
R1364 GND.n1289 GND.n1288 13.552
R1365 GND.n1187 GND.n1186 13.552
R1366 GND.n1385 GND.n1384 13.552
R1367 GND.n8998 GND.n8997 13.552
R1368 GND.n1906 GND.n1905 13.552
R1369 GND.n9094 GND.n9093 13.552
R1370 GND.n5687 GND.n5686 13.552
R1371 GND.n1912 GND.n1911 13.552
R1372 GND.n5594 GND.n5593 13.552
R1373 GND.n4428 GND.n4427 13.552
R1374 GND.n4191 GND.n4190 13.552
R1375 GND.n4335 GND.n4334 13.552
R1376 GND.n3849 GND.n3848 13.552
R1377 GND.n3618 GND.n3617 13.552
R1378 GND.n3756 GND.n3755 13.552
R1379 GND.n3316 GND.n3315 13.278
R1380 GND.n3928 GND.n3927 13.278
R1381 GND.n3692 GND.n3691 13.278
R1382 GND.n3116 GND.n3115 13.278
R1383 GND.n7650 GND.n7649 13.278
R1384 GND.n7873 GND.n7872 13.278
R1385 GND.n13155 GND.n13154 13.278
R1386 GND.n13154 GND.n13153 13.278
R1387 GND.n12004 GND.n12003 13.278
R1388 GND.n12067 GND.n12066 13.278
R1389 GND.n11837 GND.n11836 13.278
R1390 GND.n12068 GND.n12067 13.278
R1391 GND.n12003 GND.n12002 13.278
R1392 GND.n11836 GND.n11835 13.278
R1393 GND.n12217 GND.n12216 13.278
R1394 GND.n12171 GND.n12170 13.278
R1395 GND.n12172 GND.n12171 13.278
R1396 GND.n12216 GND.n12215 13.278
R1397 GND.n7649 GND.n7648 13.278
R1398 GND.n7872 GND.n7871 13.278
R1399 GND.n7343 GND.n7342 13.278
R1400 GND.n7233 GND.n7232 13.278
R1401 GND.n6196 GND.n6195 13.278
R1402 GND.n7234 GND.n7233 13.278
R1403 GND.n6195 GND.n6194 13.278
R1404 GND.n7342 GND.n7341 13.278
R1405 GND.n11177 GND.n11176 13.278
R1406 GND.n13584 GND.n13583 13.278
R1407 GND.n11176 GND.n11175 13.278
R1408 GND.n13583 GND.n13582 13.278
R1409 GND.n10540 GND.n10539 13.278
R1410 GND.n8959 GND.n8958 13.278
R1411 GND.n8923 GND.n8922 13.278
R1412 GND.n9158 GND.n9157 13.278
R1413 GND.n9660 GND.n9659 13.278
R1414 GND.n9624 GND.n9623 13.278
R1415 GND.n9859 GND.n9858 13.278
R1416 GND.n15960 GND.n15959 13.278
R1417 GND.n15924 GND.n15923 13.278
R1418 GND.n16159 GND.n16158 13.278
R1419 GND.n15925 GND.n15924 13.278
R1420 GND.n15959 GND.n15958 13.278
R1421 GND.n16158 GND.n16157 13.278
R1422 GND.n1147 GND.n1146 13.278
R1423 GND.n1146 GND.n1145 13.278
R1424 GND.n9625 GND.n9624 13.278
R1425 GND.n9659 GND.n9658 13.278
R1426 GND.n9858 GND.n9857 13.278
R1427 GND.n1210 GND.n1209 13.278
R1428 GND.n1209 GND.n1208 13.278
R1429 GND.n10277 GND.n10276 13.278
R1430 GND.n10167 GND.n10166 13.278
R1431 GND.n9998 GND.n9997 13.278
R1432 GND.n10168 GND.n10167 13.278
R1433 GND.n10276 GND.n10275 13.278
R1434 GND.n9997 GND.n9996 13.278
R1435 GND.n8737 GND.n8736 13.278
R1436 GND.n8547 GND.n8546 13.278
R1437 GND.n8437 GND.n8436 13.278
R1438 GND.n8736 GND.n8735 13.278
R1439 GND.n8438 GND.n8437 13.278
R1440 GND.n8546 GND.n8545 13.278
R1441 GND.n8924 GND.n8923 13.278
R1442 GND.n8958 GND.n8957 13.278
R1443 GND.n9157 GND.n9156 13.278
R1444 GND.n5766 GND.n5765 13.278
R1445 GND.n5765 GND.n5764 13.278
R1446 GND.n4469 GND.n4468 13.278
R1447 GND.n4519 GND.n4518 13.278
R1448 GND.n4520 GND.n4519 13.278
R1449 GND.n4468 GND.n4467 13.278
R1450 GND.n15247 GND.n15246 13.278
R1451 GND.n3115 GND.n3114 13.278
R1452 GND.n3315 GND.n3314 13.278
R1453 GND.n10539 GND.n10538 13.278
R1454 GND.n15246 GND.n15245 13.278
R1455 GND.n3691 GND.n3690 13.278
R1456 GND.n3927 GND.n3926 13.278
R1457 GND.n15063 GND.n15062 13.176
R1458 GND.n14970 GND.n14969 13.176
R1459 GND.n14670 GND.n14669 13.176
R1460 GND.n14619 GND.n14618 13.176
R1461 GND.n15822 GND.n15821 13.176
R1462 GND.n10625 GND.n10624 13.176
R1463 GND.n15481 GND.n15480 13.176
R1464 GND.n14262 GND.n14261 13.176
R1465 GND.n14347 GND.n14346 13.176
R1466 GND.n2914 GND.n2913 13.176
R1467 GND.n3567 GND.n3566 13.176
R1468 GND.n4837 GND.n4836 13.176
R1469 GND.n5149 GND.n5148 13.176
R1470 GND.n7533 GND.n7532 13.176
R1471 GND.n12760 GND.n12759 13.176
R1472 GND.n13947 GND.n13946 13.176
R1473 GND.n10757 GND.n10756 13.176
R1474 GND.n13773 GND.n13772 13.176
R1475 GND.n13817 GND.n13816 13.176
R1476 GND.n11569 GND.n11568 13.176
R1477 GND.n11673 GND.n11672 13.176
R1478 GND.n11369 GND.n11368 13.176
R1479 GND.n11059 GND.n11058 13.176
R1480 GND.n13272 GND.n13271 13.176
R1481 GND.n8209 GND.n8208 13.176
R1482 GND.n8298 GND.n8297 13.176
R1483 GND.n6458 GND.n6457 13.176
R1484 GND.n6347 GND.n6346 13.176
R1485 GND.n5983 GND.n5982 13.176
R1486 GND.n6660 GND.n6659 13.176
R1487 GND.n6895 GND.n6894 13.176
R1488 GND.n6757 GND.n6756 13.176
R1489 GND.n7481 GND.n7480 13.176
R1490 GND.n8647 GND.n8646 13.176
R1491 GND.n9342 GND.n9341 13.176
R1492 GND.n1747 GND.n1746 13.176
R1493 GND.n9467 GND.n9466 13.176
R1494 GND.n1849 GND.n1848 13.176
R1495 GND.n2540 GND.n2539 13.176
R1496 GND.n3448 GND.n3447 13.176
R1497 GND.n2446 GND.n2445 13.176
R1498 GND.n2378 GND.n2377 13.176
R1499 GND.n2105 GND.n2104 13.176
R1500 GND.n2187 GND.n2186 13.176
R1501 GND.n15377 GND.n15376 13.176
R1502 GND.n14008 GND.n14005 12.423
R1503 GND.n15543 GND.n15540 12.423
R1504 GND.n11743 GND.n11740 12.047
R1505 GND.n12484 GND.n12481 12.047
R1506 GND.n10361 GND.n10358 12.047
R1507 GND.n9937 GND.n9934 12.047
R1508 GND.n2975 GND.n2974 11.939
R1509 GND.n12842 GND.n12841 11.939
R1510 GND.n15887 GND.n15886 11.939
R1511 GND.n810 GND.n809 11.939
R1512 GND.n5819 GND.n5816 11.294
R1513 GND.n1903 GND.n1900 11.294
R1514 GND.n4756 GND.n4753 10.541
R1515 GND.n5224 GND.n5221 10.541
R1516 GND.n14469 GND.n14468 10.328
R1517 GND.n15302 GND.n15301 10.328
R1518 GND.n14483 GND.n14482 10.328
R1519 GND.n15434 GND.n15433 10.328
R1520 GND.n15744 GND.n15743 10.328
R1521 GND.n15733 GND.n15732 10.328
R1522 GND.n14091 GND.n14090 10.328
R1523 GND.n14108 GND.n14107 10.328
R1524 GND.n2663 GND.n2662 10.328
R1525 GND.n4912 GND.n4911 10.328
R1526 GND.n1949 GND.n1948 10.328
R1527 GND.n4778 GND.n4777 10.328
R1528 GND.n7189 GND.n7188 10.328
R1529 GND.n7178 GND.n7177 10.328
R1530 GND.n7408 GND.n7407 10.328
R1531 GND.n7391 GND.n7390 10.328
R1532 GND.n10776 GND.n10775 10.328
R1533 GND.n13874 GND.n13873 10.328
R1534 GND.n10884 GND.n10883 10.328
R1535 GND.n10895 GND.n10894 10.328
R1536 GND.n11117 GND.n11116 10.328
R1537 GND.n11134 GND.n11133 10.328
R1538 GND.n13525 GND.n13524 10.328
R1539 GND.n13536 GND.n13535 10.328
R1540 GND.n6037 GND.n6036 10.328
R1541 GND.n6054 GND.n6053 10.328
R1542 GND.n8242 GND.n8241 10.328
R1543 GND.n5906 GND.n5905 10.328
R1544 GND.n9269 GND.n9268 10.328
R1545 GND.n9286 GND.n9285 10.328
R1546 GND.n1575 GND.n1574 10.328
R1547 GND.n1691 GND.n1690 10.328
R1548 GND.n3373 GND.n3372 10.328
R1549 GND.n3390 GND.n3389 10.328
R1550 GND.n3169 GND.n3168 10.328
R1551 GND.n2484 GND.n2483 10.328
R1552 GND.n3970 GND.n3967 10.24
R1553 GND.n3977 GND.n3974 10.24
R1554 GND.n3984 GND.n3981 10.24
R1555 GND.n3991 GND.n3988 10.24
R1556 GND.n4005 GND.n3995 10.24
R1557 GND.n4012 GND.n4009 10.24
R1558 GND.n4019 GND.n4016 10.24
R1559 GND.n4026 GND.n4023 10.24
R1560 GND.n4033 GND.n4030 10.24
R1561 GND.n4043 GND.n4037 10.24
R1562 GND.n4043 GND.n4040 10.24
R1563 GND.n4080 GND.n4077 10.24
R1564 GND.n4087 GND.n4084 10.24
R1565 GND.n4094 GND.n4091 10.24
R1566 GND.n4101 GND.n4098 10.24
R1567 GND.n4122 GND.n4119 10.24
R1568 GND.n4129 GND.n4126 10.24
R1569 GND.n4136 GND.n4133 10.24
R1570 GND.n4143 GND.n4140 10.24
R1571 GND.n4153 GND.n4147 10.24
R1572 GND.n2684 GND.n2682 10.24
R1573 GND.n2689 GND.n2687 10.24
R1574 GND.n2694 GND.n2692 10.24
R1575 GND.n2699 GND.n2697 10.24
R1576 GND.n2704 GND.n2702 10.24
R1577 GND.n2712 GND.n2710 10.24
R1578 GND.n2717 GND.n2715 10.24
R1579 GND.n2722 GND.n2720 10.24
R1580 GND.n2729 GND.n2725 10.24
R1581 GND.n2729 GND.n2727 10.24
R1582 GND.n2758 GND.n2756 10.24
R1583 GND.n2763 GND.n2761 10.24
R1584 GND.n2768 GND.n2766 10.24
R1585 GND.n2773 GND.n2771 10.24
R1586 GND.n2781 GND.n2779 10.24
R1587 GND.n2786 GND.n2784 10.24
R1588 GND.n2791 GND.n2789 10.24
R1589 GND.n2796 GND.n2794 10.24
R1590 GND.n2803 GND.n2799 10.24
R1591 GND.n3281 GND.n3280 10.189
R1592 GND.n3945 GND.n3944 10.189
R1593 GND.n3729 GND.n3728 10.189
R1594 GND.n3081 GND.n3080 10.189
R1595 GND.n7056 GND.n7054 10.189
R1596 GND.n7090 GND.n7088 10.189
R1597 GND.n8081 GND.n8079 10.189
R1598 GND.n8047 GND.n8045 10.189
R1599 GND.n7682 GND.n7678 10.189
R1600 GND.n7838 GND.n7837 10.189
R1601 GND.n13406 GND.n13404 10.189
R1602 GND.n13440 GND.n13438 10.189
R1603 GND.n12633 GND.n12631 10.189
R1604 GND.n12599 GND.n12597 10.189
R1605 GND.n13187 GND.n13183 10.189
R1606 GND.n12900 GND.n12895 10.189
R1607 GND.n12979 GND.n12977 10.189
R1608 GND.n11874 GND.n11873 10.189
R1609 GND.n12457 GND.n12452 10.189
R1610 GND.n12350 GND.n12348 10.189
R1611 GND.n6233 GND.n6232 10.189
R1612 GND.n11214 GND.n11213 10.189
R1613 GND.n13621 GND.n13620 10.189
R1614 GND.n10505 GND.n10504 10.189
R1615 GND.n14845 GND.n14843 10.189
R1616 GND.n14811 GND.n14809 10.189
R1617 GND.n9123 GND.n9122 10.189
R1618 GND.n9824 GND.n9823 10.189
R1619 GND.n16124 GND.n16123 10.189
R1620 GND.n1164 GND.n1163 10.189
R1621 GND.n880 GND.n879 10.189
R1622 GND.n947 GND.n945 10.189
R1623 GND.n1227 GND.n1226 10.189
R1624 GND.n1518 GND.n1517 10.189
R1625 GND.n1416 GND.n1414 10.189
R1626 GND.n10035 GND.n10034 10.189
R1627 GND.n8774 GND.n8773 10.189
R1628 GND.n5783 GND.n5782 10.189
R1629 GND.n5499 GND.n5498 10.189
R1630 GND.n5566 GND.n5564 10.189
R1631 GND.n4240 GND.n4239 10.189
R1632 GND.n4307 GND.n4305 10.189
R1633 GND.n15618 GND.n15616 10.189
R1634 GND.n15652 GND.n15650 10.189
R1635 GND.n15212 GND.n15211 10.189
R1636 GND.n4683 GND.n4681 10.189
R1637 GND.n4649 GND.n4647 10.189
R1638 GND.n5029 GND.n5027 10.189
R1639 GND.n4995 GND.n4993 10.189
R1640 GND.n3328 GND.n3327 10.016
R1641 GND.n3936 GND.n3935 10.016
R1642 GND.n3679 GND.n3678 10.016
R1643 GND.n3128 GND.n3127 10.016
R1644 GND.n7004 GND.n7003 10.016
R1645 GND.n7137 GND.n7136 10.016
R1646 GND.n8129 GND.n8128 10.016
R1647 GND.n7994 GND.n7993 10.016
R1648 GND.n7664 GND.n7663 10.016
R1649 GND.n13354 GND.n13353 10.016
R1650 GND.n13487 GND.n13486 10.016
R1651 GND.n12681 GND.n12680 10.016
R1652 GND.n12546 GND.n12545 10.016
R1653 GND.n12547 GND.n12546 10.016
R1654 GND.n13488 GND.n13487 10.016
R1655 GND.n13353 GND.n13352 10.016
R1656 GND.n12680 GND.n12679 10.016
R1657 GND.n13169 GND.n13168 10.016
R1658 GND.n12863 GND.n12862 10.016
R1659 GND.n12927 GND.n12926 10.016
R1660 GND.n12862 GND.n12861 10.016
R1661 GND.n12928 GND.n12927 10.016
R1662 GND.n13168 GND.n13167 10.016
R1663 GND.n12420 GND.n12419 10.016
R1664 GND.n12397 GND.n12396 10.016
R1665 GND.n12419 GND.n12418 10.016
R1666 GND.n12398 GND.n12397 10.016
R1667 GND.n7663 GND.n7662 10.016
R1668 GND.n7138 GND.n7137 10.016
R1669 GND.n7003 GND.n7002 10.016
R1670 GND.n8128 GND.n8127 10.016
R1671 GND.n7995 GND.n7994 10.016
R1672 GND.n6183 GND.n6182 10.016
R1673 GND.n6182 GND.n6181 10.016
R1674 GND.n11165 GND.n11164 10.016
R1675 GND.n13572 GND.n13571 10.016
R1676 GND.n11164 GND.n11163 10.016
R1677 GND.n13571 GND.n13570 10.016
R1678 GND.n10552 GND.n10551 10.016
R1679 GND.n14893 GND.n14892 10.016
R1680 GND.n14758 GND.n14757 10.016
R1681 GND.n9170 GND.n9169 10.016
R1682 GND.n9871 GND.n9870 10.016
R1683 GND.n16171 GND.n16170 10.016
R1684 GND.n16170 GND.n16169 10.016
R1685 GND.n1155 GND.n1154 10.016
R1686 GND.n848 GND.n847 10.016
R1687 GND.n894 GND.n893 10.016
R1688 GND.n895 GND.n894 10.016
R1689 GND.n847 GND.n846 10.016
R1690 GND.n1154 GND.n1153 10.016
R1691 GND.n9870 GND.n9869 10.016
R1692 GND.n1218 GND.n1217 10.016
R1693 GND.n1486 GND.n1485 10.016
R1694 GND.n1463 GND.n1462 10.016
R1695 GND.n1464 GND.n1463 10.016
R1696 GND.n1485 GND.n1484 10.016
R1697 GND.n1217 GND.n1216 10.016
R1698 GND.n9985 GND.n9984 10.016
R1699 GND.n9984 GND.n9983 10.016
R1700 GND.n8725 GND.n8724 10.016
R1701 GND.n8724 GND.n8723 10.016
R1702 GND.n9169 GND.n9168 10.016
R1703 GND.n5774 GND.n5773 10.016
R1704 GND.n5467 GND.n5466 10.016
R1705 GND.n5513 GND.n5512 10.016
R1706 GND.n5514 GND.n5513 10.016
R1707 GND.n5466 GND.n5465 10.016
R1708 GND.n5773 GND.n5772 10.016
R1709 GND.n4208 GND.n4207 10.016
R1710 GND.n4254 GND.n4253 10.016
R1711 GND.n4255 GND.n4254 10.016
R1712 GND.n4207 GND.n4206 10.016
R1713 GND.n15566 GND.n15565 10.016
R1714 GND.n15699 GND.n15698 10.016
R1715 GND.n15700 GND.n15699 10.016
R1716 GND.n15565 GND.n15564 10.016
R1717 GND.n4731 GND.n4730 10.016
R1718 GND.n4596 GND.n4595 10.016
R1719 GND.n5077 GND.n5076 10.016
R1720 GND.n4942 GND.n4941 10.016
R1721 GND.n4597 GND.n4596 10.016
R1722 GND.n4943 GND.n4942 10.016
R1723 GND.n4730 GND.n4729 10.016
R1724 GND.n5076 GND.n5075 10.016
R1725 GND.n3127 GND.n3126 10.016
R1726 GND.n3327 GND.n3326 10.016
R1727 GND.n14759 GND.n14758 10.016
R1728 GND.n10551 GND.n10550 10.016
R1729 GND.n14892 GND.n14891 10.016
R1730 GND.n3678 GND.n3677 10.016
R1731 GND.n3935 GND.n3934 10.016
R1732 GND.n3190 GND.n3189 9.944
R1733 GND.n3143 GND.n3142 9.944
R1734 GND.n13344 GND.n13343 9.944
R1735 GND.n12523 GND.n12522 9.944
R1736 GND.n3248 GND.n3247 9.861
R1737 GND.n3853 GND.n3852 9.861
R1738 GND.n3648 GND.n3647 9.861
R1739 GND.n3048 GND.n3047 9.861
R1740 GND.n7748 GND.n7747 9.861
R1741 GND.n7939 GND.n7938 9.861
R1742 GND.n13073 GND.n13072 9.861
R1743 GND.n12050 GND.n12044 9.861
R1744 GND.n11794 GND.n11793 9.861
R1745 GND.n11967 GND.n11966 9.861
R1746 GND.n12154 GND.n12148 9.861
R1747 GND.n12260 GND.n12259 9.861
R1748 GND.n7272 GND.n7271 9.861
R1749 GND.n6264 GND.n6263 9.861
R1750 GND.n7306 GND.n7305 9.861
R1751 GND.n11245 GND.n11244 9.861
R1752 GND.n13652 GND.n13651 9.861
R1753 GND.n10472 GND.n10471 9.861
R1754 GND.n8912 GND.n8910 9.861
R1755 GND.n9207 GND.n9206 9.861
R1756 GND.n9613 GND.n9611 9.861
R1757 GND.n9908 GND.n9907 9.861
R1758 GND.n15913 GND.n15911 9.861
R1759 GND.n16208 GND.n16207 9.861
R1760 GND.n16003 GND.n16002 9.861
R1761 GND.n1072 GND.n1071 9.861
R1762 GND.n9703 GND.n9702 9.861
R1763 GND.n1293 GND.n1292 9.861
R1764 GND.n10206 GND.n10205 9.861
R1765 GND.n10066 GND.n10065 9.861
R1766 GND.n10240 GND.n10239 9.861
R1767 GND.n8805 GND.n8804 9.861
R1768 GND.n8476 GND.n8475 9.861
R1769 GND.n8510 GND.n8509 9.861
R1770 GND.n9002 GND.n9001 9.861
R1771 GND.n5691 GND.n5690 9.861
R1772 GND.n4508 GND.n4506 9.861
R1773 GND.n4432 GND.n4431 9.861
R1774 GND.n15179 GND.n15178 9.861
R1775 GND.n4160 GND.n4159 9.728
R1776 GND.n2808 GND.n2807 9.728
R1777 GND.n16508 GND.n16507 9.304
R1778 GND.n16769 GND.n16768 9.304
R1779 GND.n17030 GND.n17029 9.304
R1780 GND.n17291 GND.n17290 9.304
R1781 GND.n17552 GND.n17551 9.304
R1782 GND.n683 GND.n682 9.304
R1783 GND.n729 GND.n728 9.304
R1784 GND.n425 GND.n424 9.304
R1785 GND.n471 GND.n470 9.304
R1786 GND.n167 GND.n166 9.304
R1787 GND.n213 GND.n212 9.304
R1788 GND.n17782 GND.n17781 9.304
R1789 GND.n17723 GND.n17722 9.304
R1790 GND.n14666 GND.n14665 9.3
R1791 GND.n14673 GND.n14672 9.3
R1792 GND.n14680 GND.n14679 9.3
R1793 GND.n14687 GND.n14686 9.3
R1794 GND.n14694 GND.n14693 9.3
R1795 GND.n14701 GND.n14700 9.3
R1796 GND.n14708 GND.n14707 9.3
R1797 GND.n14713 GND.n14712 9.3
R1798 GND.n14497 GND.n14496 9.3
R1799 GND.n14515 GND.n14514 9.3
R1800 GND.n14476 GND.n14475 9.3
R1801 GND.n14644 GND.n14643 9.3
R1802 GND.n14502 GND.n14501 9.3
R1803 GND.n14526 GND.n14525 9.3
R1804 GND.n14521 GND.n14520 9.3
R1805 GND.n14517 GND.n14516 9.3
R1806 GND.n14511 GND.n14510 9.3
R1807 GND.n14507 GND.n14506 9.3
R1808 GND.n14640 GND.n14639 9.3
R1809 GND.n14646 GND.n14645 9.3
R1810 GND.n14711 GND.n14710 9.3
R1811 GND.n14706 GND.n14705 9.3
R1812 GND.n14704 GND.n14703 9.3
R1813 GND.n14699 GND.n14698 9.3
R1814 GND.n14697 GND.n14696 9.3
R1815 GND.n14692 GND.n14691 9.3
R1816 GND.n14690 GND.n14689 9.3
R1817 GND.n14685 GND.n14684 9.3
R1818 GND.n14683 GND.n14682 9.3
R1819 GND.n14678 GND.n14677 9.3
R1820 GND.n14676 GND.n14675 9.3
R1821 GND.n14671 GND.n14670 9.3
R1822 GND.n14668 GND.n14667 9.3
R1823 GND.n14664 GND.n14663 9.3
R1824 GND.n14657 GND.n14656 9.3
R1825 GND.n14492 GND.n14491 9.3
R1826 GND.n14717 GND.n14716 9.3
R1827 GND.n14715 GND.n14714 9.3
R1828 GND.n14622 GND.n14621 9.3
R1829 GND.n14615 GND.n14614 9.3
R1830 GND.n14608 GND.n14607 9.3
R1831 GND.n14601 GND.n14600 9.3
R1832 GND.n14594 GND.n14593 9.3
R1833 GND.n14386 GND.n14385 9.3
R1834 GND.n14393 GND.n14392 9.3
R1835 GND.n14398 GND.n14397 9.3
R1836 GND.n14371 GND.n14370 9.3
R1837 GND.n14558 GND.n14557 9.3
R1838 GND.n14569 GND.n14568 9.3
R1839 GND.n14578 GND.n14577 9.3
R1840 GND.n14541 GND.n14540 9.3
R1841 GND.n14546 GND.n14545 9.3
R1842 GND.n14552 GND.n14551 9.3
R1843 GND.n14556 GND.n14555 9.3
R1844 GND.n14563 GND.n14562 9.3
R1845 GND.n14567 GND.n14566 9.3
R1846 GND.n14574 GND.n14573 9.3
R1847 GND.n14580 GND.n14579 9.3
R1848 GND.n14396 GND.n14395 9.3
R1849 GND.n14391 GND.n14390 9.3
R1850 GND.n14389 GND.n14388 9.3
R1851 GND.n14384 GND.n14383 9.3
R1852 GND.n14382 GND.n14381 9.3
R1853 GND.n14596 GND.n14595 9.3
R1854 GND.n14599 GND.n14598 9.3
R1855 GND.n14603 GND.n14602 9.3
R1856 GND.n14606 GND.n14605 9.3
R1857 GND.n14610 GND.n14609 9.3
R1858 GND.n14613 GND.n14612 9.3
R1859 GND.n14617 GND.n14616 9.3
R1860 GND.n14620 GND.n14619 9.3
R1861 GND.n14625 GND.n14624 9.3
R1862 GND.n14591 GND.n14590 9.3
R1863 GND.n15450 GND.n15449 9.3
R1864 GND.n14402 GND.n14401 9.3
R1865 GND.n14400 GND.n14399 9.3
R1866 GND.n10581 GND.n10580 9.3
R1867 GND.n10586 GND.n10585 9.3
R1868 GND.n10593 GND.n10592 9.3
R1869 GND.n10600 GND.n10599 9.3
R1870 GND.n10607 GND.n10606 9.3
R1871 GND.n10614 GND.n10613 9.3
R1872 GND.n10621 GND.n10620 9.3
R1873 GND.n10628 GND.n10627 9.3
R1874 GND.n10651 GND.n10650 9.3
R1875 GND.n10659 GND.n10658 9.3
R1876 GND.n10584 GND.n10583 9.3
R1877 GND.n10588 GND.n10587 9.3
R1878 GND.n10591 GND.n10590 9.3
R1879 GND.n10595 GND.n10594 9.3
R1880 GND.n10598 GND.n10597 9.3
R1881 GND.n10602 GND.n10601 9.3
R1882 GND.n10605 GND.n10604 9.3
R1883 GND.n10609 GND.n10608 9.3
R1884 GND.n10612 GND.n10611 9.3
R1885 GND.n10616 GND.n10615 9.3
R1886 GND.n10619 GND.n10618 9.3
R1887 GND.n10623 GND.n10622 9.3
R1888 GND.n10626 GND.n10625 9.3
R1889 GND.n10631 GND.n10630 9.3
R1890 GND.n10636 GND.n10635 9.3
R1891 GND.n10649 GND.n10648 9.3
R1892 GND.n10656 GND.n10655 9.3
R1893 GND.n10661 GND.n10660 9.3
R1894 GND.n10666 GND.n10665 9.3
R1895 GND.n10579 GND.n10578 9.3
R1896 GND.n10577 GND.n10576 9.3
R1897 GND.n10679 GND.n10678 9.3
R1898 GND.n10685 GND.n10684 9.3
R1899 GND.n10688 GND.n10687 9.3
R1900 GND.n10693 GND.n10692 9.3
R1901 GND.n10676 GND.n10675 9.3
R1902 GND.n10671 GND.n10670 9.3
R1903 GND.n10669 GND.n10668 9.3
R1904 GND.n15526 GND.n15525 9.3
R1905 GND.n15521 GND.n15520 9.3
R1906 GND.n15514 GND.n15513 9.3
R1907 GND.n15507 GND.n15506 9.3
R1908 GND.n15500 GND.n15499 9.3
R1909 GND.n15493 GND.n15492 9.3
R1910 GND.n15486 GND.n15485 9.3
R1911 GND.n15479 GND.n15478 9.3
R1912 GND.n14074 GND.n14073 9.3
R1913 GND.n14066 GND.n14065 9.3
R1914 GND.n15524 GND.n15523 9.3
R1915 GND.n15519 GND.n15518 9.3
R1916 GND.n15517 GND.n15516 9.3
R1917 GND.n15512 GND.n15511 9.3
R1918 GND.n15510 GND.n15509 9.3
R1919 GND.n15505 GND.n15504 9.3
R1920 GND.n15503 GND.n15502 9.3
R1921 GND.n15498 GND.n15497 9.3
R1922 GND.n15496 GND.n15495 9.3
R1923 GND.n15491 GND.n15490 9.3
R1924 GND.n15489 GND.n15488 9.3
R1925 GND.n15484 GND.n15483 9.3
R1926 GND.n15482 GND.n15481 9.3
R1927 GND.n15477 GND.n15476 9.3
R1928 GND.n15472 GND.n15471 9.3
R1929 GND.n14076 GND.n14075 9.3
R1930 GND.n14070 GND.n14069 9.3
R1931 GND.n14064 GND.n14063 9.3
R1932 GND.n14060 GND.n14059 9.3
R1933 GND.n15528 GND.n15527 9.3
R1934 GND.n15530 GND.n15529 9.3
R1935 GND.n14047 GND.n14046 9.3
R1936 GND.n14043 GND.n14042 9.3
R1937 GND.n14039 GND.n14038 9.3
R1938 GND.n14035 GND.n14034 9.3
R1939 GND.n14051 GND.n14050 9.3
R1940 GND.n14054 GND.n14053 9.3
R1941 GND.n14056 GND.n14055 9.3
R1942 GND.n14147 GND.n14146 9.3
R1943 GND.n14158 GND.n14157 9.3
R1944 GND.n14301 GND.n14300 9.3
R1945 GND.n14350 GND.n14349 9.3
R1946 GND.n14343 GND.n14342 9.3
R1947 GND.n14336 GND.n14335 9.3
R1948 GND.n14329 GND.n14328 9.3
R1949 GND.n14322 GND.n14321 9.3
R1950 GND.n10698 GND.n10697 9.3
R1951 GND.n10705 GND.n10704 9.3
R1952 GND.n10710 GND.n10709 9.3
R1953 GND.n10708 GND.n10707 9.3
R1954 GND.n10703 GND.n10702 9.3
R1955 GND.n10701 GND.n10700 9.3
R1956 GND.n10696 GND.n10695 9.3
R1957 GND.n14320 GND.n14319 9.3
R1958 GND.n14324 GND.n14323 9.3
R1959 GND.n14327 GND.n14326 9.3
R1960 GND.n14331 GND.n14330 9.3
R1961 GND.n14334 GND.n14333 9.3
R1962 GND.n14338 GND.n14337 9.3
R1963 GND.n14341 GND.n14340 9.3
R1964 GND.n14345 GND.n14344 9.3
R1965 GND.n14348 GND.n14347 9.3
R1966 GND.n14353 GND.n14352 9.3
R1967 GND.n14317 GND.n14316 9.3
R1968 GND.n14303 GND.n14302 9.3
R1969 GND.n14296 GND.n14295 9.3
R1970 GND.n14156 GND.n14155 9.3
R1971 GND.n14152 GND.n14151 9.3
R1972 GND.n14145 GND.n14144 9.3
R1973 GND.n14141 GND.n14140 9.3
R1974 GND.n14135 GND.n14134 9.3
R1975 GND.n14131 GND.n14130 9.3
R1976 GND.n14126 GND.n14125 9.3
R1977 GND.n14121 GND.n14120 9.3
R1978 GND.n10714 GND.n10713 9.3
R1979 GND.n10712 GND.n10711 9.3
R1980 GND.n14200 GND.n14199 9.3
R1981 GND.n14211 GND.n14210 9.3
R1982 GND.n14285 GND.n14284 9.3
R1983 GND.n14267 GND.n14266 9.3
R1984 GND.n14260 GND.n14259 9.3
R1985 GND.n14253 GND.n14252 9.3
R1986 GND.n14246 GND.n14245 9.3
R1987 GND.n14239 GND.n14238 9.3
R1988 GND.n14232 GND.n14231 9.3
R1989 GND.n14225 GND.n14224 9.3
R1990 GND.n14220 GND.n14219 9.3
R1991 GND.n14223 GND.n14222 9.3
R1992 GND.n14227 GND.n14226 9.3
R1993 GND.n14230 GND.n14229 9.3
R1994 GND.n14234 GND.n14233 9.3
R1995 GND.n14237 GND.n14236 9.3
R1996 GND.n14241 GND.n14240 9.3
R1997 GND.n14244 GND.n14243 9.3
R1998 GND.n14248 GND.n14247 9.3
R1999 GND.n14251 GND.n14250 9.3
R2000 GND.n14255 GND.n14254 9.3
R2001 GND.n14258 GND.n14257 9.3
R2002 GND.n14263 GND.n14262 9.3
R2003 GND.n14265 GND.n14264 9.3
R2004 GND.n14270 GND.n14269 9.3
R2005 GND.n14276 GND.n14275 9.3
R2006 GND.n14283 GND.n14282 9.3
R2007 GND.n14289 GND.n14288 9.3
R2008 GND.n14209 GND.n14208 9.3
R2009 GND.n14205 GND.n14204 9.3
R2010 GND.n14198 GND.n14197 9.3
R2011 GND.n14194 GND.n14193 9.3
R2012 GND.n14188 GND.n14187 9.3
R2013 GND.n14173 GND.n14172 9.3
R2014 GND.n14168 GND.n14167 9.3
R2015 GND.n14163 GND.n14162 9.3
R2016 GND.n10575 GND.n10574 9.3
R2017 GND.n14218 GND.n14217 9.3
R2018 GND.n3546 GND.n3545 9.3
R2019 GND.n3538 GND.n3537 9.3
R2020 GND.n3528 GND.n3527 9.3
R2021 GND.n3510 GND.n3509 9.3
R2022 GND.n3548 GND.n3547 9.3
R2023 GND.n3542 GND.n3541 9.3
R2024 GND.n3514 GND.n3513 9.3
R2025 GND.n3518 GND.n3517 9.3
R2026 GND.n3522 GND.n3521 9.3
R2027 GND.n3526 GND.n3525 9.3
R2028 GND.n3532 GND.n3531 9.3
R2029 GND.n3536 GND.n3535 9.3
R2030 GND.n3612 GND.n3611 9.3
R2031 GND.n3607 GND.n3606 9.3
R2032 GND.n3600 GND.n3599 9.3
R2033 GND.n3593 GND.n3592 9.3
R2034 GND.n3586 GND.n3585 9.3
R2035 GND.n3579 GND.n3578 9.3
R2036 GND.n3572 GND.n3571 9.3
R2037 GND.n3610 GND.n3609 9.3
R2038 GND.n3605 GND.n3604 9.3
R2039 GND.n3603 GND.n3602 9.3
R2040 GND.n3598 GND.n3597 9.3
R2041 GND.n3596 GND.n3595 9.3
R2042 GND.n3591 GND.n3590 9.3
R2043 GND.n3589 GND.n3588 9.3
R2044 GND.n3584 GND.n3583 9.3
R2045 GND.n3582 GND.n3581 9.3
R2046 GND.n3577 GND.n3576 9.3
R2047 GND.n3575 GND.n3574 9.3
R2048 GND.n3570 GND.n3569 9.3
R2049 GND.n3568 GND.n3567 9.3
R2050 GND.n3563 GND.n3562 9.3
R2051 GND.n3565 GND.n3564 9.3
R2052 GND.n3614 GND.n3613 9.3
R2053 GND.n3616 GND.n3615 9.3
R2054 GND.n3506 GND.n3505 9.3
R2055 GND.n3558 GND.n3557 9.3
R2056 GND.n4862 GND.n4861 9.3
R2057 GND.n4870 GND.n4869 9.3
R2058 GND.n4880 GND.n4879 9.3
R2059 GND.n4899 GND.n4898 9.3
R2060 GND.n4860 GND.n4859 9.3
R2061 GND.n4867 GND.n4866 9.3
R2062 GND.n4896 GND.n4895 9.3
R2063 GND.n4890 GND.n4889 9.3
R2064 GND.n4887 GND.n4886 9.3
R2065 GND.n4882 GND.n4881 9.3
R2066 GND.n4877 GND.n4876 9.3
R2067 GND.n4872 GND.n4871 9.3
R2068 GND.n4793 GND.n4792 9.3
R2069 GND.n4798 GND.n4797 9.3
R2070 GND.n4805 GND.n4804 9.3
R2071 GND.n4812 GND.n4811 9.3
R2072 GND.n4819 GND.n4818 9.3
R2073 GND.n4826 GND.n4825 9.3
R2074 GND.n4833 GND.n4832 9.3
R2075 GND.n4796 GND.n4795 9.3
R2076 GND.n4800 GND.n4799 9.3
R2077 GND.n4803 GND.n4802 9.3
R2078 GND.n4807 GND.n4806 9.3
R2079 GND.n4810 GND.n4809 9.3
R2080 GND.n4814 GND.n4813 9.3
R2081 GND.n4817 GND.n4816 9.3
R2082 GND.n4821 GND.n4820 9.3
R2083 GND.n4824 GND.n4823 9.3
R2084 GND.n4828 GND.n4827 9.3
R2085 GND.n4831 GND.n4830 9.3
R2086 GND.n4835 GND.n4834 9.3
R2087 GND.n4838 GND.n4837 9.3
R2088 GND.n4843 GND.n4842 9.3
R2089 GND.n4840 GND.n4839 9.3
R2090 GND.n4791 GND.n4790 9.3
R2091 GND.n4789 GND.n4788 9.3
R2092 GND.n4903 GND.n4902 9.3
R2093 GND.n4848 GND.n4847 9.3
R2094 GND.n10760 GND.n10759 9.3
R2095 GND.n10753 GND.n10752 9.3
R2096 GND.n10746 GND.n10745 9.3
R2097 GND.n10739 GND.n10738 9.3
R2098 GND.n10852 GND.n10851 9.3
R2099 GND.n10859 GND.n10858 9.3
R2100 GND.n10866 GND.n10865 9.3
R2101 GND.n10871 GND.n10870 9.3
R2102 GND.n10819 GND.n10818 9.3
R2103 GND.n10827 GND.n10826 9.3
R2104 GND.n10813 GND.n10812 9.3
R2105 GND.n10817 GND.n10816 9.3
R2106 GND.n10823 GND.n10822 9.3
R2107 GND.n10829 GND.n10828 9.3
R2108 GND.n10869 GND.n10868 9.3
R2109 GND.n10864 GND.n10863 9.3
R2110 GND.n10862 GND.n10861 9.3
R2111 GND.n10857 GND.n10856 9.3
R2112 GND.n10855 GND.n10854 9.3
R2113 GND.n10850 GND.n10849 9.3
R2114 GND.n10737 GND.n10736 9.3
R2115 GND.n10741 GND.n10740 9.3
R2116 GND.n10744 GND.n10743 9.3
R2117 GND.n10748 GND.n10747 9.3
R2118 GND.n10751 GND.n10750 9.3
R2119 GND.n10755 GND.n10754 9.3
R2120 GND.n10758 GND.n10757 9.3
R2121 GND.n10763 GND.n10762 9.3
R2122 GND.n10767 GND.n10766 9.3
R2123 GND.n10809 GND.n10808 9.3
R2124 GND.n10807 GND.n10806 9.3
R2125 GND.n10803 GND.n10802 9.3
R2126 GND.n10799 GND.n10798 9.3
R2127 GND.n10794 GND.n10793 9.3
R2128 GND.n10790 GND.n10789 9.3
R2129 GND.n10785 GND.n10784 9.3
R2130 GND.n10875 GND.n10874 9.3
R2131 GND.n10873 GND.n10872 9.3
R2132 GND.n13943 GND.n13942 9.3
R2133 GND.n13950 GND.n13949 9.3
R2134 GND.n13957 GND.n13956 9.3
R2135 GND.n13964 GND.n13963 9.3
R2136 GND.n13971 GND.n13970 9.3
R2137 GND.n13978 GND.n13977 9.3
R2138 GND.n13985 GND.n13984 9.3
R2139 GND.n13990 GND.n13989 9.3
R2140 GND.n13890 GND.n13889 9.3
R2141 GND.n13908 GND.n13907 9.3
R2142 GND.n13918 GND.n13917 9.3
R2143 GND.n13926 GND.n13925 9.3
R2144 GND.n13894 GND.n13893 9.3
R2145 GND.n13898 GND.n13897 9.3
R2146 GND.n13902 GND.n13901 9.3
R2147 GND.n13906 GND.n13905 9.3
R2148 GND.n13912 GND.n13911 9.3
R2149 GND.n13916 GND.n13915 9.3
R2150 GND.n13922 GND.n13921 9.3
R2151 GND.n13928 GND.n13927 9.3
R2152 GND.n13988 GND.n13987 9.3
R2153 GND.n13983 GND.n13982 9.3
R2154 GND.n13981 GND.n13980 9.3
R2155 GND.n13976 GND.n13975 9.3
R2156 GND.n13974 GND.n13973 9.3
R2157 GND.n13969 GND.n13968 9.3
R2158 GND.n13967 GND.n13966 9.3
R2159 GND.n13962 GND.n13961 9.3
R2160 GND.n13960 GND.n13959 9.3
R2161 GND.n13955 GND.n13954 9.3
R2162 GND.n13953 GND.n13952 9.3
R2163 GND.n13948 GND.n13947 9.3
R2164 GND.n13945 GND.n13944 9.3
R2165 GND.n13941 GND.n13940 9.3
R2166 GND.n13935 GND.n13934 9.3
R2167 GND.n13885 GND.n13884 9.3
R2168 GND.n13994 GND.n13993 9.3
R2169 GND.n13992 GND.n13991 9.3
R2170 GND.n13862 GND.n13861 9.3
R2171 GND.n13857 GND.n13856 9.3
R2172 GND.n13850 GND.n13849 9.3
R2173 GND.n13843 GND.n13842 9.3
R2174 GND.n13836 GND.n13835 9.3
R2175 GND.n13829 GND.n13828 9.3
R2176 GND.n13822 GND.n13821 9.3
R2177 GND.n13815 GND.n13814 9.3
R2178 GND.n10946 GND.n10945 9.3
R2179 GND.n10938 GND.n10937 9.3
R2180 GND.n13860 GND.n13859 9.3
R2181 GND.n13855 GND.n13854 9.3
R2182 GND.n13853 GND.n13852 9.3
R2183 GND.n13848 GND.n13847 9.3
R2184 GND.n13846 GND.n13845 9.3
R2185 GND.n13841 GND.n13840 9.3
R2186 GND.n13839 GND.n13838 9.3
R2187 GND.n13834 GND.n13833 9.3
R2188 GND.n13832 GND.n13831 9.3
R2189 GND.n13827 GND.n13826 9.3
R2190 GND.n13825 GND.n13824 9.3
R2191 GND.n13820 GND.n13819 9.3
R2192 GND.n13818 GND.n13817 9.3
R2193 GND.n13813 GND.n13812 9.3
R2194 GND.n13808 GND.n13807 9.3
R2195 GND.n10948 GND.n10947 9.3
R2196 GND.n10942 GND.n10941 9.3
R2197 GND.n10936 GND.n10935 9.3
R2198 GND.n10932 GND.n10931 9.3
R2199 GND.n13864 GND.n13863 9.3
R2200 GND.n13866 GND.n13865 9.3
R2201 GND.n10919 GND.n10918 9.3
R2202 GND.n10915 GND.n10914 9.3
R2203 GND.n10911 GND.n10910 9.3
R2204 GND.n10907 GND.n10906 9.3
R2205 GND.n10923 GND.n10922 9.3
R2206 GND.n10926 GND.n10925 9.3
R2207 GND.n10928 GND.n10927 9.3
R2208 GND.n13729 GND.n13728 9.3
R2209 GND.n13734 GND.n13733 9.3
R2210 GND.n13741 GND.n13740 9.3
R2211 GND.n13748 GND.n13747 9.3
R2212 GND.n13755 GND.n13754 9.3
R2213 GND.n13762 GND.n13761 9.3
R2214 GND.n13769 GND.n13768 9.3
R2215 GND.n13776 GND.n13775 9.3
R2216 GND.n10995 GND.n10994 9.3
R2217 GND.n10987 GND.n10986 9.3
R2218 GND.n13732 GND.n13731 9.3
R2219 GND.n13736 GND.n13735 9.3
R2220 GND.n13739 GND.n13738 9.3
R2221 GND.n13743 GND.n13742 9.3
R2222 GND.n13746 GND.n13745 9.3
R2223 GND.n13750 GND.n13749 9.3
R2224 GND.n13753 GND.n13752 9.3
R2225 GND.n13757 GND.n13756 9.3
R2226 GND.n13760 GND.n13759 9.3
R2227 GND.n13764 GND.n13763 9.3
R2228 GND.n13767 GND.n13766 9.3
R2229 GND.n13771 GND.n13770 9.3
R2230 GND.n13774 GND.n13773 9.3
R2231 GND.n13779 GND.n13778 9.3
R2232 GND.n13783 GND.n13782 9.3
R2233 GND.n10997 GND.n10996 9.3
R2234 GND.n10991 GND.n10990 9.3
R2235 GND.n10985 GND.n10984 9.3
R2236 GND.n10981 GND.n10980 9.3
R2237 GND.n13727 GND.n13726 9.3
R2238 GND.n13725 GND.n13724 9.3
R2239 GND.n10968 GND.n10967 9.3
R2240 GND.n10964 GND.n10963 9.3
R2241 GND.n10960 GND.n10959 9.3
R2242 GND.n10956 GND.n10955 9.3
R2243 GND.n10972 GND.n10971 9.3
R2244 GND.n10975 GND.n10974 9.3
R2245 GND.n10977 GND.n10976 9.3
R2246 GND.n11312 GND.n11311 9.3
R2247 GND.n11286 GND.n11285 9.3
R2248 GND.n11274 GND.n11273 9.3
R2249 GND.n11262 GND.n11261 9.3
R2250 GND.n11250 GND.n11249 9.3
R2251 GND.n11238 GND.n11237 9.3
R2252 GND.n11220 GND.n11219 9.3
R2253 GND.n11208 GND.n11207 9.3
R2254 GND.n11196 GND.n11195 9.3
R2255 GND.n11184 GND.n11183 9.3
R2256 GND.n11172 GND.n11171 9.3
R2257 GND.n11160 GND.n11159 9.3
R2258 GND.n11147 GND.n11146 9.3
R2259 GND.n11310 GND.n11309 9.3
R2260 GND.n11288 GND.n11287 9.3
R2261 GND.n11276 GND.n11275 9.3
R2262 GND.n11264 GND.n11263 9.3
R2263 GND.n11252 GND.n11251 9.3
R2264 GND.n11240 GND.n11239 9.3
R2265 GND.n11218 GND.n11217 9.3
R2266 GND.n11206 GND.n11205 9.3
R2267 GND.n11194 GND.n11193 9.3
R2268 GND.n11182 GND.n11181 9.3
R2269 GND.n11170 GND.n11169 9.3
R2270 GND.n11158 GND.n11157 9.3
R2271 GND.n11006 GND.n11005 9.3
R2272 GND.n11298 GND.n11297 9.3
R2273 GND.n11300 GND.n11299 9.3
R2274 GND.n13554 GND.n13553 9.3
R2275 GND.n13567 GND.n13566 9.3
R2276 GND.n13579 GND.n13578 9.3
R2277 GND.n13591 GND.n13590 9.3
R2278 GND.n13603 GND.n13602 9.3
R2279 GND.n13615 GND.n13614 9.3
R2280 GND.n13627 GND.n13626 9.3
R2281 GND.n13645 GND.n13644 9.3
R2282 GND.n13657 GND.n13656 9.3
R2283 GND.n13669 GND.n13668 9.3
R2284 GND.n13681 GND.n13680 9.3
R2285 GND.n13693 GND.n13692 9.3
R2286 GND.n13705 GND.n13704 9.3
R2287 GND.n13717 GND.n13716 9.3
R2288 GND.n10717 GND.n10716 9.3
R2289 GND.n13565 GND.n13564 9.3
R2290 GND.n13577 GND.n13576 9.3
R2291 GND.n13589 GND.n13588 9.3
R2292 GND.n13601 GND.n13600 9.3
R2293 GND.n13613 GND.n13612 9.3
R2294 GND.n13625 GND.n13624 9.3
R2295 GND.n13647 GND.n13646 9.3
R2296 GND.n13659 GND.n13658 9.3
R2297 GND.n13671 GND.n13670 9.3
R2298 GND.n13683 GND.n13682 9.3
R2299 GND.n13695 GND.n13694 9.3
R2300 GND.n13707 GND.n13706 9.3
R2301 GND.n13719 GND.n13718 9.3
R2302 GND.n10724 GND.n10723 9.3
R2303 GND.n10879 GND.n10878 9.3
R2304 GND.n10877 GND.n10876 9.3
R2305 GND.n10887 GND.n10886 9.3
R2306 GND.n10886 GND.n10885 9.3
R2307 GND.n10898 GND.n10897 9.3
R2308 GND.n10897 GND.n10896 9.3
R2309 GND.n13996 GND.n13995 9.3
R2310 GND.n12714 GND.n12713 9.3
R2311 GND.n12721 GND.n12720 9.3
R2312 GND.n12728 GND.n12727 9.3
R2313 GND.n12735 GND.n12734 9.3
R2314 GND.n12742 GND.n12741 9.3
R2315 GND.n12749 GND.n12748 9.3
R2316 GND.n12756 GND.n12755 9.3
R2317 GND.n12763 GND.n12762 9.3
R2318 GND.n12785 GND.n12784 9.3
R2319 GND.n12793 GND.n12792 9.3
R2320 GND.n12783 GND.n12782 9.3
R2321 GND.n12790 GND.n12789 9.3
R2322 GND.n12795 GND.n12794 9.3
R2323 GND.n12800 GND.n12799 9.3
R2324 GND.n12771 GND.n12770 9.3
R2325 GND.n12766 GND.n12765 9.3
R2326 GND.n12761 GND.n12760 9.3
R2327 GND.n12758 GND.n12757 9.3
R2328 GND.n12754 GND.n12753 9.3
R2329 GND.n12751 GND.n12750 9.3
R2330 GND.n12747 GND.n12746 9.3
R2331 GND.n12744 GND.n12743 9.3
R2332 GND.n12740 GND.n12739 9.3
R2333 GND.n12737 GND.n12736 9.3
R2334 GND.n12733 GND.n12732 9.3
R2335 GND.n12730 GND.n12729 9.3
R2336 GND.n12726 GND.n12725 9.3
R2337 GND.n12723 GND.n12722 9.3
R2338 GND.n12719 GND.n12718 9.3
R2339 GND.n12716 GND.n12715 9.3
R2340 GND.n12712 GND.n12711 9.3
R2341 GND.n12813 GND.n12812 9.3
R2342 GND.n12819 GND.n12818 9.3
R2343 GND.n12822 GND.n12821 9.3
R2344 GND.n12827 GND.n12826 9.3
R2345 GND.n12810 GND.n12809 9.3
R2346 GND.n12805 GND.n12804 9.3
R2347 GND.n12803 GND.n12802 9.3
R2348 GND.n13879 GND.n13878 9.3
R2349 GND.n10781 GND.n10780 9.3
R2350 GND.n10771 GND.n10770 9.3
R2351 GND.n10779 GND.n10778 9.3
R2352 GND.n10778 GND.n10777 9.3
R2353 GND.n13877 GND.n13876 9.3
R2354 GND.n13876 GND.n13875 9.3
R2355 GND.n13881 GND.n13880 9.3
R2356 GND.n12699 GND.n12698 9.3
R2357 GND.n12687 GND.n12686 9.3
R2358 GND.n12674 GND.n12673 9.3
R2359 GND.n12662 GND.n12661 9.3
R2360 GND.n12649 GND.n12648 9.3
R2361 GND.n12637 GND.n12636 9.3
R2362 GND.n12624 GND.n12623 9.3
R2363 GND.n12605 GND.n12604 9.3
R2364 GND.n12592 GND.n12591 9.3
R2365 GND.n12580 GND.n12579 9.3
R2366 GND.n12567 GND.n12566 9.3
R2367 GND.n12555 GND.n12554 9.3
R2368 GND.n12542 GND.n12541 9.3
R2369 GND.n12540 GND.n12539 9.3
R2370 GND.n12551 GND.n12550 9.3
R2371 GND.n12550 GND.n12549 9.3
R2372 GND.n12553 GND.n12552 9.3
R2373 GND.n12563 GND.n12562 9.3
R2374 GND.n12562 GND.n12561 9.3
R2375 GND.n12565 GND.n12564 9.3
R2376 GND.n12576 GND.n12575 9.3
R2377 GND.n12575 GND.n12574 9.3
R2378 GND.n12578 GND.n12577 9.3
R2379 GND.n12588 GND.n12587 9.3
R2380 GND.n12587 GND.n12586 9.3
R2381 GND.n12590 GND.n12589 9.3
R2382 GND.n12601 GND.n12600 9.3
R2383 GND.n12600 GND.n12599 9.3
R2384 GND.n12603 GND.n12602 9.3
R2385 GND.n12614 GND.n12613 9.3
R2386 GND.n12613 GND.n12612 9.3
R2387 GND.n12622 GND.n12621 9.3
R2388 GND.n12621 GND.n12620 9.3
R2389 GND.n12626 GND.n12625 9.3
R2390 GND.n12635 GND.n12634 9.3
R2391 GND.n12634 GND.n12633 9.3
R2392 GND.n12639 GND.n12638 9.3
R2393 GND.n12647 GND.n12646 9.3
R2394 GND.n12646 GND.n12645 9.3
R2395 GND.n12651 GND.n12650 9.3
R2396 GND.n12660 GND.n12659 9.3
R2397 GND.n12659 GND.n12658 9.3
R2398 GND.n12664 GND.n12663 9.3
R2399 GND.n12672 GND.n12671 9.3
R2400 GND.n12671 GND.n12670 9.3
R2401 GND.n12676 GND.n12675 9.3
R2402 GND.n12685 GND.n12684 9.3
R2403 GND.n12684 GND.n12683 9.3
R2404 GND.n12689 GND.n12688 9.3
R2405 GND.n12697 GND.n12696 9.3
R2406 GND.n12696 GND.n12695 9.3
R2407 GND.n12701 GND.n12700 9.3
R2408 GND.n11669 GND.n11668 9.3
R2409 GND.n11676 GND.n11675 9.3
R2410 GND.n11683 GND.n11682 9.3
R2411 GND.n11690 GND.n11689 9.3
R2412 GND.n11697 GND.n11696 9.3
R2413 GND.n11704 GND.n11703 9.3
R2414 GND.n11711 GND.n11710 9.3
R2415 GND.n11716 GND.n11715 9.3
R2416 GND.n11480 GND.n11479 9.3
R2417 GND.n11488 GND.n11487 9.3
R2418 GND.n11474 GND.n11473 9.3
R2419 GND.n11478 GND.n11477 9.3
R2420 GND.n11484 GND.n11483 9.3
R2421 GND.n11490 GND.n11489 9.3
R2422 GND.n11714 GND.n11713 9.3
R2423 GND.n11709 GND.n11708 9.3
R2424 GND.n11707 GND.n11706 9.3
R2425 GND.n11702 GND.n11701 9.3
R2426 GND.n11700 GND.n11699 9.3
R2427 GND.n11695 GND.n11694 9.3
R2428 GND.n11693 GND.n11692 9.3
R2429 GND.n11688 GND.n11687 9.3
R2430 GND.n11686 GND.n11685 9.3
R2431 GND.n11681 GND.n11680 9.3
R2432 GND.n11679 GND.n11678 9.3
R2433 GND.n11674 GND.n11673 9.3
R2434 GND.n11671 GND.n11670 9.3
R2435 GND.n11667 GND.n11666 9.3
R2436 GND.n11661 GND.n11660 9.3
R2437 GND.n11470 GND.n11469 9.3
R2438 GND.n11468 GND.n11467 9.3
R2439 GND.n11464 GND.n11463 9.3
R2440 GND.n11460 GND.n11459 9.3
R2441 GND.n11455 GND.n11454 9.3
R2442 GND.n11451 GND.n11450 9.3
R2443 GND.n11446 GND.n11445 9.3
R2444 GND.n11720 GND.n11719 9.3
R2445 GND.n11718 GND.n11717 9.3
R2446 GND.n11565 GND.n11564 9.3
R2447 GND.n11572 GND.n11571 9.3
R2448 GND.n11579 GND.n11578 9.3
R2449 GND.n11586 GND.n11585 9.3
R2450 GND.n11593 GND.n11592 9.3
R2451 GND.n11600 GND.n11599 9.3
R2452 GND.n11607 GND.n11606 9.3
R2453 GND.n11612 GND.n11611 9.3
R2454 GND.n11512 GND.n11511 9.3
R2455 GND.n11530 GND.n11529 9.3
R2456 GND.n11540 GND.n11539 9.3
R2457 GND.n11548 GND.n11547 9.3
R2458 GND.n11516 GND.n11515 9.3
R2459 GND.n11520 GND.n11519 9.3
R2460 GND.n11524 GND.n11523 9.3
R2461 GND.n11528 GND.n11527 9.3
R2462 GND.n11534 GND.n11533 9.3
R2463 GND.n11538 GND.n11537 9.3
R2464 GND.n11544 GND.n11543 9.3
R2465 GND.n11550 GND.n11549 9.3
R2466 GND.n11610 GND.n11609 9.3
R2467 GND.n11605 GND.n11604 9.3
R2468 GND.n11603 GND.n11602 9.3
R2469 GND.n11598 GND.n11597 9.3
R2470 GND.n11596 GND.n11595 9.3
R2471 GND.n11591 GND.n11590 9.3
R2472 GND.n11589 GND.n11588 9.3
R2473 GND.n11584 GND.n11583 9.3
R2474 GND.n11582 GND.n11581 9.3
R2475 GND.n11577 GND.n11576 9.3
R2476 GND.n11575 GND.n11574 9.3
R2477 GND.n11570 GND.n11569 9.3
R2478 GND.n11567 GND.n11566 9.3
R2479 GND.n11563 GND.n11562 9.3
R2480 GND.n11557 GND.n11556 9.3
R2481 GND.n11507 GND.n11506 9.3
R2482 GND.n11616 GND.n11615 9.3
R2483 GND.n11614 GND.n11613 9.3
R2484 GND.n11104 GND.n11103 9.3
R2485 GND.n11099 GND.n11098 9.3
R2486 GND.n11092 GND.n11091 9.3
R2487 GND.n11085 GND.n11084 9.3
R2488 GND.n11078 GND.n11077 9.3
R2489 GND.n11071 GND.n11070 9.3
R2490 GND.n11064 GND.n11063 9.3
R2491 GND.n11057 GND.n11056 9.3
R2492 GND.n11025 GND.n11024 9.3
R2493 GND.n11618 GND.n11617 9.3
R2494 GND.n11102 GND.n11101 9.3
R2495 GND.n11097 GND.n11096 9.3
R2496 GND.n11095 GND.n11094 9.3
R2497 GND.n11090 GND.n11089 9.3
R2498 GND.n11088 GND.n11087 9.3
R2499 GND.n11083 GND.n11082 9.3
R2500 GND.n11081 GND.n11080 9.3
R2501 GND.n11076 GND.n11075 9.3
R2502 GND.n11074 GND.n11073 9.3
R2503 GND.n11069 GND.n11068 9.3
R2504 GND.n11067 GND.n11066 9.3
R2505 GND.n11062 GND.n11061 9.3
R2506 GND.n11060 GND.n11059 9.3
R2507 GND.n11055 GND.n11054 9.3
R2508 GND.n11050 GND.n11049 9.3
R2509 GND.n11027 GND.n11026 9.3
R2510 GND.n11021 GND.n11020 9.3
R2511 GND.n11620 GND.n11619 9.3
R2512 GND.n11625 GND.n11624 9.3
R2513 GND.n11106 GND.n11105 9.3
R2514 GND.n11108 GND.n11107 9.3
R2515 GND.n11638 GND.n11637 9.3
R2516 GND.n11644 GND.n11643 9.3
R2517 GND.n11647 GND.n11646 9.3
R2518 GND.n11652 GND.n11651 9.3
R2519 GND.n11635 GND.n11634 9.3
R2520 GND.n11630 GND.n11629 9.3
R2521 GND.n11628 GND.n11627 9.3
R2522 GND.n13319 GND.n13318 9.3
R2523 GND.n13312 GND.n13311 9.3
R2524 GND.n13305 GND.n13304 9.3
R2525 GND.n13298 GND.n13297 9.3
R2526 GND.n13291 GND.n13290 9.3
R2527 GND.n13284 GND.n13283 9.3
R2528 GND.n13277 GND.n13276 9.3
R2529 GND.n13270 GND.n13269 9.3
R2530 GND.n13250 GND.n13249 9.3
R2531 GND.n13242 GND.n13241 9.3
R2532 GND.n13252 GND.n13251 9.3
R2533 GND.n13246 GND.n13245 9.3
R2534 GND.n13240 GND.n13239 9.3
R2535 GND.n13236 GND.n13235 9.3
R2536 GND.n13263 GND.n13262 9.3
R2537 GND.n13268 GND.n13267 9.3
R2538 GND.n13273 GND.n13272 9.3
R2539 GND.n13275 GND.n13274 9.3
R2540 GND.n13280 GND.n13279 9.3
R2541 GND.n13282 GND.n13281 9.3
R2542 GND.n13287 GND.n13286 9.3
R2543 GND.n13289 GND.n13288 9.3
R2544 GND.n13294 GND.n13293 9.3
R2545 GND.n13296 GND.n13295 9.3
R2546 GND.n13301 GND.n13300 9.3
R2547 GND.n13303 GND.n13302 9.3
R2548 GND.n13308 GND.n13307 9.3
R2549 GND.n13310 GND.n13309 9.3
R2550 GND.n13315 GND.n13314 9.3
R2551 GND.n13317 GND.n13316 9.3
R2552 GND.n13321 GND.n13320 9.3
R2553 GND.n13223 GND.n13222 9.3
R2554 GND.n13219 GND.n13218 9.3
R2555 GND.n13215 GND.n13214 9.3
R2556 GND.n13211 GND.n13210 9.3
R2557 GND.n13227 GND.n13226 9.3
R2558 GND.n13230 GND.n13229 9.3
R2559 GND.n13232 GND.n13231 9.3
R2560 GND.n11325 GND.n11324 9.3
R2561 GND.n11330 GND.n11329 9.3
R2562 GND.n11337 GND.n11336 9.3
R2563 GND.n11344 GND.n11343 9.3
R2564 GND.n11351 GND.n11350 9.3
R2565 GND.n11358 GND.n11357 9.3
R2566 GND.n11365 GND.n11364 9.3
R2567 GND.n11372 GND.n11371 9.3
R2568 GND.n11392 GND.n11391 9.3
R2569 GND.n11400 GND.n11399 9.3
R2570 GND.n11328 GND.n11327 9.3
R2571 GND.n11332 GND.n11331 9.3
R2572 GND.n11335 GND.n11334 9.3
R2573 GND.n11339 GND.n11338 9.3
R2574 GND.n11342 GND.n11341 9.3
R2575 GND.n11346 GND.n11345 9.3
R2576 GND.n11349 GND.n11348 9.3
R2577 GND.n11353 GND.n11352 9.3
R2578 GND.n11356 GND.n11355 9.3
R2579 GND.n11360 GND.n11359 9.3
R2580 GND.n11363 GND.n11362 9.3
R2581 GND.n11367 GND.n11366 9.3
R2582 GND.n11370 GND.n11369 9.3
R2583 GND.n11375 GND.n11374 9.3
R2584 GND.n11379 GND.n11378 9.3
R2585 GND.n11390 GND.n11389 9.3
R2586 GND.n11397 GND.n11396 9.3
R2587 GND.n11402 GND.n11401 9.3
R2588 GND.n11407 GND.n11406 9.3
R2589 GND.n11323 GND.n11322 9.3
R2590 GND.n11321 GND.n11320 9.3
R2591 GND.n11420 GND.n11419 9.3
R2592 GND.n11426 GND.n11425 9.3
R2593 GND.n11429 GND.n11428 9.3
R2594 GND.n11433 GND.n11432 9.3
R2595 GND.n11417 GND.n11416 9.3
R2596 GND.n11412 GND.n11411 9.3
R2597 GND.n11410 GND.n11409 9.3
R2598 GND.n13541 GND.n13540 9.3
R2599 GND.n13520 GND.n13519 9.3
R2600 GND.n13544 GND.n13543 9.3
R2601 GND.n13539 GND.n13538 9.3
R2602 GND.n13538 GND.n13537 9.3
R2603 GND.n13528 GND.n13527 9.3
R2604 GND.n13527 GND.n13526 9.3
R2605 GND.n13517 GND.n13516 9.3
R2606 GND.n13358 GND.n13357 9.3
R2607 GND.n13357 GND.n13356 9.3
R2608 GND.n13362 GND.n13361 9.3
R2609 GND.n13374 GND.n13373 9.3
R2610 GND.n13387 GND.n13386 9.3
R2611 GND.n13399 GND.n13398 9.3
R2612 GND.n13412 GND.n13411 9.3
R2613 GND.n13431 GND.n13430 9.3
R2614 GND.n13444 GND.n13443 9.3
R2615 GND.n13456 GND.n13455 9.3
R2616 GND.n13469 GND.n13468 9.3
R2617 GND.n13481 GND.n13480 9.3
R2618 GND.n13494 GND.n13493 9.3
R2619 GND.n13360 GND.n13359 9.3
R2620 GND.n13370 GND.n13369 9.3
R2621 GND.n13369 GND.n13368 9.3
R2622 GND.n13372 GND.n13371 9.3
R2623 GND.n13383 GND.n13382 9.3
R2624 GND.n13382 GND.n13381 9.3
R2625 GND.n13385 GND.n13384 9.3
R2626 GND.n13395 GND.n13394 9.3
R2627 GND.n13394 GND.n13393 9.3
R2628 GND.n13397 GND.n13396 9.3
R2629 GND.n13408 GND.n13407 9.3
R2630 GND.n13407 GND.n13406 9.3
R2631 GND.n13410 GND.n13409 9.3
R2632 GND.n13420 GND.n13419 9.3
R2633 GND.n13419 GND.n13418 9.3
R2634 GND.n13429 GND.n13428 9.3
R2635 GND.n13428 GND.n13427 9.3
R2636 GND.n13433 GND.n13432 9.3
R2637 GND.n13442 GND.n13441 9.3
R2638 GND.n13441 GND.n13440 9.3
R2639 GND.n13446 GND.n13445 9.3
R2640 GND.n13454 GND.n13453 9.3
R2641 GND.n13453 GND.n13452 9.3
R2642 GND.n13458 GND.n13457 9.3
R2643 GND.n13467 GND.n13466 9.3
R2644 GND.n13466 GND.n13465 9.3
R2645 GND.n13471 GND.n13470 9.3
R2646 GND.n13479 GND.n13478 9.3
R2647 GND.n13478 GND.n13477 9.3
R2648 GND.n13483 GND.n13482 9.3
R2649 GND.n13492 GND.n13491 9.3
R2650 GND.n13491 GND.n13490 9.3
R2651 GND.n13496 GND.n13495 9.3
R2652 GND.n13504 GND.n13503 9.3
R2653 GND.n13503 GND.n13502 9.3
R2654 GND.n13508 GND.n13507 9.3
R2655 GND.n13506 GND.n13505 9.3
R2656 GND.n13349 GND.n13348 9.3
R2657 GND.n13347 GND.n13346 9.3
R2658 GND.n11112 GND.n11111 9.3
R2659 GND.n11139 GND.n11138 9.3
R2660 GND.n11110 GND.n11109 9.3
R2661 GND.n11120 GND.n11119 9.3
R2662 GND.n11119 GND.n11118 9.3
R2663 GND.n11137 GND.n11136 9.3
R2664 GND.n11136 GND.n11135 9.3
R2665 GND.n11141 GND.n11140 9.3
R2666 GND.n11816 GND.n11815 9.3
R2667 GND.n11815 GND.n11814 9.3
R2668 GND.n11820 GND.n11819 9.3
R2669 GND.n11832 GND.n11831 9.3
R2670 GND.n11845 GND.n11844 9.3
R2671 GND.n11857 GND.n11856 9.3
R2672 GND.n11869 GND.n11868 9.3
R2673 GND.n11900 GND.n11899 9.3
R2674 GND.n11905 GND.n11904 9.3
R2675 GND.n11910 GND.n11909 9.3
R2676 GND.n11925 GND.n11924 9.3
R2677 GND.n11930 GND.n11929 9.3
R2678 GND.n11935 GND.n11934 9.3
R2679 GND.n11940 GND.n11939 9.3
R2680 GND.n11945 GND.n11944 9.3
R2681 GND.n11972 GND.n11971 9.3
R2682 GND.n11985 GND.n11984 9.3
R2683 GND.n11997 GND.n11996 9.3
R2684 GND.n12010 GND.n12009 9.3
R2685 GND.n12022 GND.n12021 9.3
R2686 GND.n12096 GND.n12095 9.3
R2687 GND.n12024 GND.n12023 9.3
R2688 GND.n12020 GND.n12019 9.3
R2689 GND.n12019 GND.n12018 9.3
R2690 GND.n12012 GND.n12011 9.3
R2691 GND.n12008 GND.n12007 9.3
R2692 GND.n12007 GND.n12006 9.3
R2693 GND.n11999 GND.n11998 9.3
R2694 GND.n11995 GND.n11994 9.3
R2695 GND.n11994 GND.n11993 9.3
R2696 GND.n11987 GND.n11986 9.3
R2697 GND.n11983 GND.n11982 9.3
R2698 GND.n11982 GND.n11981 9.3
R2699 GND.n11974 GND.n11973 9.3
R2700 GND.n11970 GND.n11969 9.3
R2701 GND.n11969 GND.n11968 9.3
R2702 GND.n12041 GND.n12040 9.3
R2703 GND.n11952 GND.n11951 9.3
R2704 GND.n12049 GND.n12048 9.3
R2705 GND.n11948 GND.n11947 9.3
R2706 GND.n12057 GND.n12056 9.3
R2707 GND.n11943 GND.n11942 9.3
R2708 GND.n12064 GND.n12063 9.3
R2709 GND.n11938 GND.n11937 9.3
R2710 GND.n12072 GND.n12071 9.3
R2711 GND.n11933 GND.n11932 9.3
R2712 GND.n12079 GND.n12078 9.3
R2713 GND.n11928 GND.n11927 9.3
R2714 GND.n12087 GND.n12086 9.3
R2715 GND.n12088 GND.n12087 9.3
R2716 GND.n11923 GND.n11922 9.3
R2717 GND.n11912 GND.n11911 9.3
R2718 GND.n11756 GND.n11755 9.3
R2719 GND.n11907 GND.n11906 9.3
R2720 GND.n11806 GND.n11805 9.3
R2721 GND.n11902 GND.n11901 9.3
R2722 GND.n11763 GND.n11762 9.3
R2723 GND.n11897 GND.n11896 9.3
R2724 GND.n11799 GND.n11798 9.3
R2725 GND.n11893 GND.n11892 9.3
R2726 GND.n11771 GND.n11770 9.3
R2727 GND.n11889 GND.n11888 9.3
R2728 GND.n11791 GND.n11790 9.3
R2729 GND.n11885 GND.n11884 9.3
R2730 GND.n11779 GND.n11778 9.3
R2731 GND.n11810 GND.n11786 9.3
R2732 GND.n11879 GND.n11878 9.3
R2733 GND.n11875 GND.n11870 9.3
R2734 GND.n11875 GND.n11874 9.3
R2735 GND.n11867 GND.n11866 9.3
R2736 GND.n11865 GND.n11864 9.3
R2737 GND.n11864 GND.n11863 9.3
R2738 GND.n11855 GND.n11854 9.3
R2739 GND.n11853 GND.n11852 9.3
R2740 GND.n11852 GND.n11851 9.3
R2741 GND.n11843 GND.n11842 9.3
R2742 GND.n11841 GND.n11840 9.3
R2743 GND.n11840 GND.n11839 9.3
R2744 GND.n11830 GND.n11829 9.3
R2745 GND.n11818 GND.n11817 9.3
R2746 GND.n11828 GND.n11827 9.3
R2747 GND.n11827 GND.n11826 9.3
R2748 GND.n12092 GND.n12091 9.3
R2749 GND.n12091 GND.n12090 9.3
R2750 GND.n12094 GND.n12093 9.3
R2751 GND.n11750 GND.n11749 9.3
R2752 GND.n11735 GND.n11734 9.3
R2753 GND.n12476 GND.n12475 9.3
R2754 GND.n12475 GND.n12474 9.3
R2755 GND.n12404 GND.n12403 9.3
R2756 GND.n12391 GND.n12390 9.3
R2757 GND.n12379 GND.n12378 9.3
R2758 GND.n12366 GND.n12365 9.3
R2759 GND.n12354 GND.n12353 9.3
R2760 GND.n12322 GND.n12321 9.3
R2761 GND.n12317 GND.n12316 9.3
R2762 GND.n12312 GND.n12311 9.3
R2763 GND.n12297 GND.n12296 9.3
R2764 GND.n12292 GND.n12291 9.3
R2765 GND.n12287 GND.n12286 9.3
R2766 GND.n12282 GND.n12281 9.3
R2767 GND.n12277 GND.n12276 9.3
R2768 GND.n12250 GND.n12249 9.3
R2769 GND.n12237 GND.n12236 9.3
R2770 GND.n12225 GND.n12224 9.3
R2771 GND.n12212 GND.n12211 9.3
R2772 GND.n12200 GND.n12199 9.3
R2773 GND.n12126 GND.n12125 9.3
R2774 GND.n12198 GND.n12197 9.3
R2775 GND.n12208 GND.n12207 9.3
R2776 GND.n12207 GND.n12206 9.3
R2777 GND.n12210 GND.n12209 9.3
R2778 GND.n12221 GND.n12220 9.3
R2779 GND.n12220 GND.n12219 9.3
R2780 GND.n12223 GND.n12222 9.3
R2781 GND.n12233 GND.n12232 9.3
R2782 GND.n12232 GND.n12231 9.3
R2783 GND.n12235 GND.n12234 9.3
R2784 GND.n12246 GND.n12245 9.3
R2785 GND.n12245 GND.n12244 9.3
R2786 GND.n12248 GND.n12247 9.3
R2787 GND.n12263 GND.n12262 9.3
R2788 GND.n12262 GND.n12261 9.3
R2789 GND.n12145 GND.n12144 9.3
R2790 GND.n12270 GND.n12269 9.3
R2791 GND.n12153 GND.n12152 9.3
R2792 GND.n12274 GND.n12273 9.3
R2793 GND.n12161 GND.n12160 9.3
R2794 GND.n12279 GND.n12278 9.3
R2795 GND.n12168 GND.n12167 9.3
R2796 GND.n12284 GND.n12283 9.3
R2797 GND.n12176 GND.n12175 9.3
R2798 GND.n12289 GND.n12288 9.3
R2799 GND.n12183 GND.n12182 9.3
R2800 GND.n12294 GND.n12293 9.3
R2801 GND.n12191 GND.n12190 9.3
R2802 GND.n12192 GND.n12191 9.3
R2803 GND.n12299 GND.n12298 9.3
R2804 GND.n12310 GND.n12309 9.3
R2805 GND.n12414 GND.n12413 9.3
R2806 GND.n12315 GND.n12314 9.3
R2807 GND.n12424 GND.n12423 9.3
R2808 GND.n12320 GND.n12319 9.3
R2809 GND.n12429 GND.n12428 9.3
R2810 GND.n12325 GND.n12324 9.3
R2811 GND.n12440 GND.n12439 9.3
R2812 GND.n12329 GND.n12328 9.3
R2813 GND.n12446 GND.n12445 9.3
R2814 GND.n12333 GND.n12332 9.3
R2815 GND.n12457 GND.n12456 9.3
R2816 GND.n12337 GND.n12336 9.3
R2817 GND.n12463 GND.n12462 9.3
R2818 GND.n12343 GND.n12342 9.3
R2819 GND.n12352 GND.n12351 9.3
R2820 GND.n12351 GND.n12350 9.3
R2821 GND.n12356 GND.n12355 9.3
R2822 GND.n12364 GND.n12363 9.3
R2823 GND.n12363 GND.n12362 9.3
R2824 GND.n12368 GND.n12367 9.3
R2825 GND.n12377 GND.n12376 9.3
R2826 GND.n12376 GND.n12375 9.3
R2827 GND.n12381 GND.n12380 9.3
R2828 GND.n12389 GND.n12388 9.3
R2829 GND.n12388 GND.n12387 9.3
R2830 GND.n12393 GND.n12392 9.3
R2831 GND.n12406 GND.n12405 9.3
R2832 GND.n12402 GND.n12401 9.3
R2833 GND.n12401 GND.n12400 9.3
R2834 GND.n12196 GND.n12195 9.3
R2835 GND.n12195 GND.n12194 9.3
R2836 GND.n12128 GND.n12127 9.3
R2837 GND.n12478 GND.n12477 9.3
R2838 GND.n12480 GND.n12479 9.3
R2839 GND.n12919 GND.n12918 9.3
R2840 GND.n12918 GND.n12917 9.3
R2841 GND.n12923 GND.n12922 9.3
R2842 GND.n12936 GND.n12935 9.3
R2843 GND.n12948 GND.n12947 9.3
R2844 GND.n12961 GND.n12960 9.3
R2845 GND.n12973 GND.n12972 9.3
R2846 GND.n13005 GND.n13004 9.3
R2847 GND.n13010 GND.n13009 9.3
R2848 GND.n13015 GND.n13014 9.3
R2849 GND.n13030 GND.n13029 9.3
R2850 GND.n13035 GND.n13034 9.3
R2851 GND.n13040 GND.n13039 9.3
R2852 GND.n13045 GND.n13044 9.3
R2853 GND.n13050 GND.n13049 9.3
R2854 GND.n13055 GND.n13054 9.3
R2855 GND.n13078 GND.n13077 9.3
R2856 GND.n13090 GND.n13089 9.3
R2857 GND.n13102 GND.n13101 9.3
R2858 GND.n13114 GND.n13113 9.3
R2859 GND.n13126 GND.n13125 9.3
R2860 GND.n13195 GND.n13194 9.3
R2861 GND.n13128 GND.n13127 9.3
R2862 GND.n13124 GND.n13123 9.3
R2863 GND.n13123 GND.n13122 9.3
R2864 GND.n13116 GND.n13115 9.3
R2865 GND.n13112 GND.n13111 9.3
R2866 GND.n13111 GND.n13110 9.3
R2867 GND.n13104 GND.n13103 9.3
R2868 GND.n13100 GND.n13099 9.3
R2869 GND.n13099 GND.n13098 9.3
R2870 GND.n13092 GND.n13091 9.3
R2871 GND.n13088 GND.n13087 9.3
R2872 GND.n13087 GND.n13086 9.3
R2873 GND.n13080 GND.n13079 9.3
R2874 GND.n13076 GND.n13075 9.3
R2875 GND.n13075 GND.n13074 9.3
R2876 GND.n13145 GND.n13144 9.3
R2877 GND.n13188 GND.n13145 9.3
R2878 GND.n13058 GND.n13057 9.3
R2879 GND.n13187 GND.n13186 9.3
R2880 GND.n13188 GND.n13187 9.3
R2881 GND.n13053 GND.n13052 9.3
R2882 GND.n13152 GND.n13151 9.3
R2883 GND.n13188 GND.n13152 9.3
R2884 GND.n13048 GND.n13047 9.3
R2885 GND.n13180 GND.n13179 9.3
R2886 GND.n13188 GND.n13180 9.3
R2887 GND.n13043 GND.n13042 9.3
R2888 GND.n13159 GND.n13158 9.3
R2889 GND.n13188 GND.n13159 9.3
R2890 GND.n13038 GND.n13037 9.3
R2891 GND.n13173 GND.n13172 9.3
R2892 GND.n13188 GND.n13173 9.3
R2893 GND.n13033 GND.n13032 9.3
R2894 GND.n13166 GND.n13165 9.3
R2895 GND.n13188 GND.n13166 9.3
R2896 GND.n13028 GND.n13027 9.3
R2897 GND.n13017 GND.n13016 9.3
R2898 GND.n12857 GND.n12856 9.3
R2899 GND.n13012 GND.n13011 9.3
R2900 GND.n12867 GND.n12866 9.3
R2901 GND.n13007 GND.n13006 9.3
R2902 GND.n12872 GND.n12871 9.3
R2903 GND.n13002 GND.n13001 9.3
R2904 GND.n12883 GND.n12882 9.3
R2905 GND.n12998 GND.n12997 9.3
R2906 GND.n12889 GND.n12888 9.3
R2907 GND.n12994 GND.n12993 9.3
R2908 GND.n12900 GND.n12899 9.3
R2909 GND.n12990 GND.n12989 9.3
R2910 GND.n12906 GND.n12905 9.3
R2911 GND.n12984 GND.n12983 9.3
R2912 GND.n12980 GND.n12974 9.3
R2913 GND.n12980 GND.n12979 9.3
R2914 GND.n12971 GND.n12970 9.3
R2915 GND.n12969 GND.n12968 9.3
R2916 GND.n12968 GND.n12967 9.3
R2917 GND.n12959 GND.n12958 9.3
R2918 GND.n12957 GND.n12956 9.3
R2919 GND.n12956 GND.n12955 9.3
R2920 GND.n12946 GND.n12945 9.3
R2921 GND.n12944 GND.n12943 9.3
R2922 GND.n12943 GND.n12942 9.3
R2923 GND.n12934 GND.n12933 9.3
R2924 GND.n12921 GND.n12920 9.3
R2925 GND.n12932 GND.n12931 9.3
R2926 GND.n12931 GND.n12930 9.3
R2927 GND.n13191 GND.n13190 9.3
R2928 GND.n13190 GND.n13189 9.3
R2929 GND.n13189 GND.n13188 9.3
R2930 GND.n13193 GND.n13192 9.3
R2931 GND.n12849 GND.n12848 9.3
R2932 GND.n12847 GND.n12846 9.3
R2933 GND.n7959 GND.n7958 9.3
R2934 GND.n7958 GND.n7957 9.3
R2935 GND.n7891 GND.n7890 9.3
R2936 GND.n7879 GND.n7878 9.3
R2937 GND.n7866 GND.n7865 9.3
R2938 GND.n7854 GND.n7853 9.3
R2939 GND.n7842 GND.n7841 9.3
R2940 GND.n7811 GND.n7810 9.3
R2941 GND.n7806 GND.n7805 9.3
R2942 GND.n7801 GND.n7800 9.3
R2943 GND.n7786 GND.n7785 9.3
R2944 GND.n7781 GND.n7780 9.3
R2945 GND.n7776 GND.n7775 9.3
R2946 GND.n7771 GND.n7770 9.3
R2947 GND.n7766 GND.n7765 9.3
R2948 GND.n7761 GND.n7760 9.3
R2949 GND.n7738 GND.n7737 9.3
R2950 GND.n7726 GND.n7725 9.3
R2951 GND.n7714 GND.n7713 9.3
R2952 GND.n7702 GND.n7701 9.3
R2953 GND.n7690 GND.n7689 9.3
R2954 GND.n7621 GND.n7620 9.3
R2955 GND.n7688 GND.n7687 9.3
R2956 GND.n7698 GND.n7697 9.3
R2957 GND.n7697 GND.n7696 9.3
R2958 GND.n7700 GND.n7699 9.3
R2959 GND.n7710 GND.n7709 9.3
R2960 GND.n7709 GND.n7708 9.3
R2961 GND.n7712 GND.n7711 9.3
R2962 GND.n7722 GND.n7721 9.3
R2963 GND.n7721 GND.n7720 9.3
R2964 GND.n7724 GND.n7723 9.3
R2965 GND.n7734 GND.n7733 9.3
R2966 GND.n7733 GND.n7732 9.3
R2967 GND.n7736 GND.n7735 9.3
R2968 GND.n7751 GND.n7750 9.3
R2969 GND.n7750 GND.n7749 9.3
R2970 GND.n7640 GND.n7639 9.3
R2971 GND.n7683 GND.n7640 9.3
R2972 GND.n7758 GND.n7757 9.3
R2973 GND.n7682 GND.n7681 9.3
R2974 GND.n7683 GND.n7682 9.3
R2975 GND.n7763 GND.n7762 9.3
R2976 GND.n7647 GND.n7646 9.3
R2977 GND.n7683 GND.n7647 9.3
R2978 GND.n7768 GND.n7767 9.3
R2979 GND.n7675 GND.n7674 9.3
R2980 GND.n7683 GND.n7675 9.3
R2981 GND.n7773 GND.n7772 9.3
R2982 GND.n7654 GND.n7653 9.3
R2983 GND.n7683 GND.n7654 9.3
R2984 GND.n7778 GND.n7777 9.3
R2985 GND.n7668 GND.n7667 9.3
R2986 GND.n7683 GND.n7668 9.3
R2987 GND.n7783 GND.n7782 9.3
R2988 GND.n7661 GND.n7660 9.3
R2989 GND.n7683 GND.n7661 9.3
R2990 GND.n7788 GND.n7787 9.3
R2991 GND.n7799 GND.n7798 9.3
R2992 GND.n7901 GND.n7900 9.3
R2993 GND.n7804 GND.n7803 9.3
R2994 GND.n7951 GND.n7950 9.3
R2995 GND.n7809 GND.n7808 9.3
R2996 GND.n7908 GND.n7907 9.3
R2997 GND.n7814 GND.n7813 9.3
R2998 GND.n7944 GND.n7943 9.3
R2999 GND.n7818 GND.n7817 9.3
R3000 GND.n7916 GND.n7915 9.3
R3001 GND.n7822 GND.n7821 9.3
R3002 GND.n7936 GND.n7935 9.3
R3003 GND.n7826 GND.n7825 9.3
R3004 GND.n7924 GND.n7923 9.3
R3005 GND.n7955 GND.n7931 9.3
R3006 GND.n7832 GND.n7831 9.3
R3007 GND.n7840 GND.n7839 9.3
R3008 GND.n7839 GND.n7838 9.3
R3009 GND.n7844 GND.n7843 9.3
R3010 GND.n7852 GND.n7851 9.3
R3011 GND.n7851 GND.n7850 9.3
R3012 GND.n7856 GND.n7855 9.3
R3013 GND.n7864 GND.n7863 9.3
R3014 GND.n7863 GND.n7862 9.3
R3015 GND.n7868 GND.n7867 9.3
R3016 GND.n7877 GND.n7876 9.3
R3017 GND.n7876 GND.n7875 9.3
R3018 GND.n7881 GND.n7880 9.3
R3019 GND.n7893 GND.n7892 9.3
R3020 GND.n7889 GND.n7888 9.3
R3021 GND.n7888 GND.n7887 9.3
R3022 GND.n7686 GND.n7685 9.3
R3023 GND.n7685 GND.n7684 9.3
R3024 GND.n7684 GND.n7683 9.3
R3025 GND.n7623 GND.n7622 9.3
R3026 GND.n7961 GND.n7960 9.3
R3027 GND.n7963 GND.n7962 9.3
R3028 GND.n6329 GND.n6328 9.3
R3029 GND.n6317 GND.n6316 9.3
R3030 GND.n6305 GND.n6304 9.3
R3031 GND.n6293 GND.n6292 9.3
R3032 GND.n6281 GND.n6280 9.3
R3033 GND.n6269 GND.n6268 9.3
R3034 GND.n6257 GND.n6256 9.3
R3035 GND.n6239 GND.n6238 9.3
R3036 GND.n6227 GND.n6226 9.3
R3037 GND.n6215 GND.n6214 9.3
R3038 GND.n6203 GND.n6202 9.3
R3039 GND.n6191 GND.n6190 9.3
R3040 GND.n6178 GND.n6177 9.3
R3041 GND.n6165 GND.n6164 9.3
R3042 GND.n6176 GND.n6175 9.3
R3043 GND.n6189 GND.n6188 9.3
R3044 GND.n6201 GND.n6200 9.3
R3045 GND.n6213 GND.n6212 9.3
R3046 GND.n6225 GND.n6224 9.3
R3047 GND.n6237 GND.n6236 9.3
R3048 GND.n6259 GND.n6258 9.3
R3049 GND.n6271 GND.n6270 9.3
R3050 GND.n6283 GND.n6282 9.3
R3051 GND.n6295 GND.n6294 9.3
R3052 GND.n6307 GND.n6306 9.3
R3053 GND.n6319 GND.n6318 9.3
R3054 GND.n6331 GND.n6330 9.3
R3055 GND.n5822 GND.n5821 9.3
R3056 GND.n8165 GND.n8164 9.3
R3057 GND.n8170 GND.n8169 9.3
R3058 GND.n8177 GND.n8176 9.3
R3059 GND.n8184 GND.n8183 9.3
R3060 GND.n8191 GND.n8190 9.3
R3061 GND.n8198 GND.n8197 9.3
R3062 GND.n8205 GND.n8204 9.3
R3063 GND.n8212 GND.n8211 9.3
R3064 GND.n6063 GND.n6062 9.3
R3065 GND.n6071 GND.n6070 9.3
R3066 GND.n8168 GND.n8167 9.3
R3067 GND.n8172 GND.n8171 9.3
R3068 GND.n8175 GND.n8174 9.3
R3069 GND.n8179 GND.n8178 9.3
R3070 GND.n8182 GND.n8181 9.3
R3071 GND.n8186 GND.n8185 9.3
R3072 GND.n8189 GND.n8188 9.3
R3073 GND.n8193 GND.n8192 9.3
R3074 GND.n8196 GND.n8195 9.3
R3075 GND.n8200 GND.n8199 9.3
R3076 GND.n8203 GND.n8202 9.3
R3077 GND.n8207 GND.n8206 9.3
R3078 GND.n8210 GND.n8209 9.3
R3079 GND.n8215 GND.n8214 9.3
R3080 GND.n8220 GND.n8219 9.3
R3081 GND.n6061 GND.n6060 9.3
R3082 GND.n6068 GND.n6067 9.3
R3083 GND.n6073 GND.n6072 9.3
R3084 GND.n6078 GND.n6077 9.3
R3085 GND.n8163 GND.n8162 9.3
R3086 GND.n8161 GND.n8160 9.3
R3087 GND.n6091 GND.n6090 9.3
R3088 GND.n6097 GND.n6096 9.3
R3089 GND.n6100 GND.n6099 9.3
R3090 GND.n6105 GND.n6104 9.3
R3091 GND.n6088 GND.n6087 9.3
R3092 GND.n6083 GND.n6082 9.3
R3093 GND.n6081 GND.n6080 9.3
R3094 GND.n8252 GND.n8251 9.3
R3095 GND.n8259 GND.n8258 9.3
R3096 GND.n8266 GND.n8265 9.3
R3097 GND.n8273 GND.n8272 9.3
R3098 GND.n8280 GND.n8279 9.3
R3099 GND.n8287 GND.n8286 9.3
R3100 GND.n8294 GND.n8293 9.3
R3101 GND.n8301 GND.n8300 9.3
R3102 GND.n8324 GND.n8323 9.3
R3103 GND.n8332 GND.n8331 9.3
R3104 GND.n8322 GND.n8321 9.3
R3105 GND.n8329 GND.n8328 9.3
R3106 GND.n8334 GND.n8333 9.3
R3107 GND.n8339 GND.n8338 9.3
R3108 GND.n8309 GND.n8308 9.3
R3109 GND.n8304 GND.n8303 9.3
R3110 GND.n8299 GND.n8298 9.3
R3111 GND.n8296 GND.n8295 9.3
R3112 GND.n8292 GND.n8291 9.3
R3113 GND.n8289 GND.n8288 9.3
R3114 GND.n8285 GND.n8284 9.3
R3115 GND.n8282 GND.n8281 9.3
R3116 GND.n8278 GND.n8277 9.3
R3117 GND.n8275 GND.n8274 9.3
R3118 GND.n8271 GND.n8270 9.3
R3119 GND.n8268 GND.n8267 9.3
R3120 GND.n8264 GND.n8263 9.3
R3121 GND.n8261 GND.n8260 9.3
R3122 GND.n8257 GND.n8256 9.3
R3123 GND.n8254 GND.n8253 9.3
R3124 GND.n8250 GND.n8249 9.3
R3125 GND.n8352 GND.n8351 9.3
R3126 GND.n8358 GND.n8357 9.3
R3127 GND.n8361 GND.n8360 9.3
R3128 GND.n8366 GND.n8365 9.3
R3129 GND.n8349 GND.n8348 9.3
R3130 GND.n8344 GND.n8343 9.3
R3131 GND.n8342 GND.n8341 9.3
R3132 GND.n6392 GND.n6391 9.3
R3133 GND.n6370 GND.n6369 9.3
R3134 GND.n6378 GND.n6377 9.3
R3135 GND.n6350 GND.n6349 9.3
R3136 GND.n5857 GND.n5856 9.3
R3137 GND.n5864 GND.n5863 9.3
R3138 GND.n5871 GND.n5870 9.3
R3139 GND.n5878 GND.n5877 9.3
R3140 GND.n5885 GND.n5884 9.3
R3141 GND.n5892 GND.n5891 9.3
R3142 GND.n5897 GND.n5896 9.3
R3143 GND.n5895 GND.n5894 9.3
R3144 GND.n5890 GND.n5889 9.3
R3145 GND.n5888 GND.n5887 9.3
R3146 GND.n5883 GND.n5882 9.3
R3147 GND.n5881 GND.n5880 9.3
R3148 GND.n5876 GND.n5875 9.3
R3149 GND.n5874 GND.n5873 9.3
R3150 GND.n5869 GND.n5868 9.3
R3151 GND.n5867 GND.n5866 9.3
R3152 GND.n5862 GND.n5861 9.3
R3153 GND.n5860 GND.n5859 9.3
R3154 GND.n5855 GND.n5854 9.3
R3155 GND.n6348 GND.n6347 9.3
R3156 GND.n6353 GND.n6352 9.3
R3157 GND.n6356 GND.n6355 9.3
R3158 GND.n6380 GND.n6379 9.3
R3159 GND.n6374 GND.n6373 9.3
R3160 GND.n6368 GND.n6367 9.3
R3161 GND.n6389 GND.n6388 9.3
R3162 GND.n6394 GND.n6393 9.3
R3163 GND.n6398 GND.n6397 9.3
R3164 GND.n6400 GND.n6399 9.3
R3165 GND.n5840 GND.n5839 9.3
R3166 GND.n5843 GND.n5842 9.3
R3167 GND.n5847 GND.n5846 9.3
R3168 GND.n5901 GND.n5900 9.3
R3169 GND.n5899 GND.n5898 9.3
R3170 GND.n5979 GND.n5978 9.3
R3171 GND.n5986 GND.n5985 9.3
R3172 GND.n5993 GND.n5992 9.3
R3173 GND.n6000 GND.n5999 9.3
R3174 GND.n6007 GND.n6006 9.3
R3175 GND.n6014 GND.n6013 9.3
R3176 GND.n6021 GND.n6020 9.3
R3177 GND.n6026 GND.n6025 9.3
R3178 GND.n5920 GND.n5919 9.3
R3179 GND.n5939 GND.n5938 9.3
R3180 GND.n5949 GND.n5948 9.3
R3181 GND.n5957 GND.n5956 9.3
R3182 GND.n5924 GND.n5923 9.3
R3183 GND.n5929 GND.n5928 9.3
R3184 GND.n5933 GND.n5932 9.3
R3185 GND.n5937 GND.n5936 9.3
R3186 GND.n5943 GND.n5942 9.3
R3187 GND.n5947 GND.n5946 9.3
R3188 GND.n5953 GND.n5952 9.3
R3189 GND.n5959 GND.n5958 9.3
R3190 GND.n6024 GND.n6023 9.3
R3191 GND.n6019 GND.n6018 9.3
R3192 GND.n6017 GND.n6016 9.3
R3193 GND.n6012 GND.n6011 9.3
R3194 GND.n6010 GND.n6009 9.3
R3195 GND.n6005 GND.n6004 9.3
R3196 GND.n6003 GND.n6002 9.3
R3197 GND.n5998 GND.n5997 9.3
R3198 GND.n5996 GND.n5995 9.3
R3199 GND.n5991 GND.n5990 9.3
R3200 GND.n5989 GND.n5988 9.3
R3201 GND.n5984 GND.n5983 9.3
R3202 GND.n5981 GND.n5980 9.3
R3203 GND.n5977 GND.n5976 9.3
R3204 GND.n5971 GND.n5970 9.3
R3205 GND.n5915 GND.n5914 9.3
R3206 GND.n6030 GND.n6029 9.3
R3207 GND.n6028 GND.n6027 9.3
R3208 GND.n6463 GND.n6462 9.3
R3209 GND.n6456 GND.n6455 9.3
R3210 GND.n6449 GND.n6448 9.3
R3211 GND.n6442 GND.n6441 9.3
R3212 GND.n6435 GND.n6434 9.3
R3213 GND.n6428 GND.n6427 9.3
R3214 GND.n6421 GND.n6420 9.3
R3215 GND.n6416 GND.n6415 9.3
R3216 GND.n6486 GND.n6485 9.3
R3217 GND.n6479 GND.n6478 9.3
R3218 GND.n6492 GND.n6491 9.3
R3219 GND.n6488 GND.n6487 9.3
R3220 GND.n6483 GND.n6482 9.3
R3221 GND.n6477 GND.n6476 9.3
R3222 GND.n6419 GND.n6418 9.3
R3223 GND.n6423 GND.n6422 9.3
R3224 GND.n6426 GND.n6425 9.3
R3225 GND.n6430 GND.n6429 9.3
R3226 GND.n6433 GND.n6432 9.3
R3227 GND.n6437 GND.n6436 9.3
R3228 GND.n6440 GND.n6439 9.3
R3229 GND.n6444 GND.n6443 9.3
R3230 GND.n6447 GND.n6446 9.3
R3231 GND.n6451 GND.n6450 9.3
R3232 GND.n6454 GND.n6453 9.3
R3233 GND.n6459 GND.n6458 9.3
R3234 GND.n6461 GND.n6460 9.3
R3235 GND.n6466 GND.n6465 9.3
R3236 GND.n6470 GND.n6469 9.3
R3237 GND.n6495 GND.n6494 9.3
R3238 GND.n6497 GND.n6496 9.3
R3239 GND.n6501 GND.n6500 9.3
R3240 GND.n6504 GND.n6503 9.3
R3241 GND.n6509 GND.n6508 9.3
R3242 GND.n6512 GND.n6511 9.3
R3243 GND.n6516 GND.n6515 9.3
R3244 GND.n5824 GND.n5823 9.3
R3245 GND.n6414 GND.n6413 9.3
R3246 GND.n5833 GND.n5832 9.3
R3247 GND.n8247 GND.n8246 9.3
R3248 GND.n8237 GND.n8236 9.3
R3249 GND.n8245 GND.n8244 9.3
R3250 GND.n8244 GND.n8243 9.3
R3251 GND.n5909 GND.n5908 9.3
R3252 GND.n5908 GND.n5907 9.3
R3253 GND.n8158 GND.n8157 9.3
R3254 GND.n6059 GND.n6058 9.3
R3255 GND.n6032 GND.n6031 9.3
R3256 GND.n8377 GND.n8376 9.3
R3257 GND.n6108 GND.n6107 9.3
R3258 GND.n6057 GND.n6056 9.3
R3259 GND.n6056 GND.n6055 9.3
R3260 GND.n6040 GND.n6039 9.3
R3261 GND.n6039 GND.n6038 9.3
R3262 GND.n8369 GND.n8368 9.3
R3263 GND.n8375 GND.n8374 9.3
R3264 GND.n7986 GND.n7985 9.3
R3265 GND.n7985 GND.n7984 9.3
R3266 GND.n7990 GND.n7989 9.3
R3267 GND.n8003 GND.n8002 9.3
R3268 GND.n8015 GND.n8014 9.3
R3269 GND.n8028 GND.n8027 9.3
R3270 GND.n8040 GND.n8039 9.3
R3271 GND.n8053 GND.n8052 9.3
R3272 GND.n8072 GND.n8071 9.3
R3273 GND.n8085 GND.n8084 9.3
R3274 GND.n8097 GND.n8096 9.3
R3275 GND.n8110 GND.n8109 9.3
R3276 GND.n8122 GND.n8121 9.3
R3277 GND.n8135 GND.n8134 9.3
R3278 GND.n8147 GND.n8146 9.3
R3279 GND.n8149 GND.n8148 9.3
R3280 GND.n8145 GND.n8144 9.3
R3281 GND.n8144 GND.n8143 9.3
R3282 GND.n8137 GND.n8136 9.3
R3283 GND.n8133 GND.n8132 9.3
R3284 GND.n8132 GND.n8131 9.3
R3285 GND.n8124 GND.n8123 9.3
R3286 GND.n8120 GND.n8119 9.3
R3287 GND.n8119 GND.n8118 9.3
R3288 GND.n8112 GND.n8111 9.3
R3289 GND.n8108 GND.n8107 9.3
R3290 GND.n8107 GND.n8106 9.3
R3291 GND.n8099 GND.n8098 9.3
R3292 GND.n8095 GND.n8094 9.3
R3293 GND.n8094 GND.n8093 9.3
R3294 GND.n8087 GND.n8086 9.3
R3295 GND.n8083 GND.n8082 9.3
R3296 GND.n8082 GND.n8081 9.3
R3297 GND.n8074 GND.n8073 9.3
R3298 GND.n8070 GND.n8069 9.3
R3299 GND.n8069 GND.n8068 9.3
R3300 GND.n8061 GND.n8060 9.3
R3301 GND.n8060 GND.n8059 9.3
R3302 GND.n8051 GND.n8050 9.3
R3303 GND.n8049 GND.n8048 9.3
R3304 GND.n8048 GND.n8047 9.3
R3305 GND.n8038 GND.n8037 9.3
R3306 GND.n8036 GND.n8035 9.3
R3307 GND.n8035 GND.n8034 9.3
R3308 GND.n8026 GND.n8025 9.3
R3309 GND.n8024 GND.n8023 9.3
R3310 GND.n8023 GND.n8022 9.3
R3311 GND.n8013 GND.n8012 9.3
R3312 GND.n8011 GND.n8010 9.3
R3313 GND.n8010 GND.n8009 9.3
R3314 GND.n8001 GND.n8000 9.3
R3315 GND.n7988 GND.n7987 9.3
R3316 GND.n7999 GND.n7998 9.3
R3317 GND.n7998 GND.n7997 9.3
R3318 GND.n7977 GND.n7976 9.3
R3319 GND.n7975 GND.n7974 9.3
R3320 GND.n6149 GND.n6148 9.3
R3321 GND.n6995 GND.n6994 9.3
R3322 GND.n6994 GND.n6993 9.3
R3323 GND.n7008 GND.n7007 9.3
R3324 GND.n7007 GND.n7006 9.3
R3325 GND.n6987 GND.n6986 9.3
R3326 GND.n7012 GND.n7011 9.3
R3327 GND.n7024 GND.n7023 9.3
R3328 GND.n7037 GND.n7036 9.3
R3329 GND.n7049 GND.n7048 9.3
R3330 GND.n7062 GND.n7061 9.3
R3331 GND.n7081 GND.n7080 9.3
R3332 GND.n7094 GND.n7093 9.3
R3333 GND.n7106 GND.n7105 9.3
R3334 GND.n7119 GND.n7118 9.3
R3335 GND.n7131 GND.n7130 9.3
R3336 GND.n7144 GND.n7143 9.3
R3337 GND.n7010 GND.n7009 9.3
R3338 GND.n7020 GND.n7019 9.3
R3339 GND.n7019 GND.n7018 9.3
R3340 GND.n7022 GND.n7021 9.3
R3341 GND.n7033 GND.n7032 9.3
R3342 GND.n7032 GND.n7031 9.3
R3343 GND.n7035 GND.n7034 9.3
R3344 GND.n7045 GND.n7044 9.3
R3345 GND.n7044 GND.n7043 9.3
R3346 GND.n7047 GND.n7046 9.3
R3347 GND.n7058 GND.n7057 9.3
R3348 GND.n7057 GND.n7056 9.3
R3349 GND.n7060 GND.n7059 9.3
R3350 GND.n7070 GND.n7069 9.3
R3351 GND.n7069 GND.n7068 9.3
R3352 GND.n7079 GND.n7078 9.3
R3353 GND.n7078 GND.n7077 9.3
R3354 GND.n7083 GND.n7082 9.3
R3355 GND.n7092 GND.n7091 9.3
R3356 GND.n7091 GND.n7090 9.3
R3357 GND.n7096 GND.n7095 9.3
R3358 GND.n7104 GND.n7103 9.3
R3359 GND.n7103 GND.n7102 9.3
R3360 GND.n7108 GND.n7107 9.3
R3361 GND.n7117 GND.n7116 9.3
R3362 GND.n7116 GND.n7115 9.3
R3363 GND.n7121 GND.n7120 9.3
R3364 GND.n7129 GND.n7128 9.3
R3365 GND.n7128 GND.n7127 9.3
R3366 GND.n7133 GND.n7132 9.3
R3367 GND.n7142 GND.n7141 9.3
R3368 GND.n7141 GND.n7140 9.3
R3369 GND.n7146 GND.n7145 9.3
R3370 GND.n7155 GND.n7154 9.3
R3371 GND.n7154 GND.n7153 9.3
R3372 GND.n7159 GND.n7158 9.3
R3373 GND.n7157 GND.n7156 9.3
R3374 GND.n6999 GND.n6998 9.3
R3375 GND.n6997 GND.n6996 9.3
R3376 GND.n6891 GND.n6890 9.3
R3377 GND.n6898 GND.n6897 9.3
R3378 GND.n6905 GND.n6904 9.3
R3379 GND.n6912 GND.n6911 9.3
R3380 GND.n6919 GND.n6918 9.3
R3381 GND.n6926 GND.n6925 9.3
R3382 GND.n6933 GND.n6932 9.3
R3383 GND.n6938 GND.n6937 9.3
R3384 GND.n6833 GND.n6832 9.3
R3385 GND.n6852 GND.n6851 9.3
R3386 GND.n6862 GND.n6861 9.3
R3387 GND.n6870 GND.n6869 9.3
R3388 GND.n6837 GND.n6836 9.3
R3389 GND.n6842 GND.n6841 9.3
R3390 GND.n6846 GND.n6845 9.3
R3391 GND.n6850 GND.n6849 9.3
R3392 GND.n6856 GND.n6855 9.3
R3393 GND.n6860 GND.n6859 9.3
R3394 GND.n6866 GND.n6865 9.3
R3395 GND.n6872 GND.n6871 9.3
R3396 GND.n6936 GND.n6935 9.3
R3397 GND.n6931 GND.n6930 9.3
R3398 GND.n6929 GND.n6928 9.3
R3399 GND.n6924 GND.n6923 9.3
R3400 GND.n6922 GND.n6921 9.3
R3401 GND.n6917 GND.n6916 9.3
R3402 GND.n6915 GND.n6914 9.3
R3403 GND.n6910 GND.n6909 9.3
R3404 GND.n6908 GND.n6907 9.3
R3405 GND.n6903 GND.n6902 9.3
R3406 GND.n6901 GND.n6900 9.3
R3407 GND.n6896 GND.n6895 9.3
R3408 GND.n6893 GND.n6892 9.3
R3409 GND.n6889 GND.n6888 9.3
R3410 GND.n6883 GND.n6882 9.3
R3411 GND.n6828 GND.n6827 9.3
R3412 GND.n6942 GND.n6941 9.3
R3413 GND.n6940 GND.n6939 9.3
R3414 GND.n6656 GND.n6655 9.3
R3415 GND.n6663 GND.n6662 9.3
R3416 GND.n6670 GND.n6669 9.3
R3417 GND.n6677 GND.n6676 9.3
R3418 GND.n6684 GND.n6683 9.3
R3419 GND.n6691 GND.n6690 9.3
R3420 GND.n6698 GND.n6697 9.3
R3421 GND.n6703 GND.n6702 9.3
R3422 GND.n6627 GND.n6626 9.3
R3423 GND.n6635 GND.n6634 9.3
R3424 GND.n6621 GND.n6620 9.3
R3425 GND.n6625 GND.n6624 9.3
R3426 GND.n6631 GND.n6630 9.3
R3427 GND.n6637 GND.n6636 9.3
R3428 GND.n6701 GND.n6700 9.3
R3429 GND.n6696 GND.n6695 9.3
R3430 GND.n6694 GND.n6693 9.3
R3431 GND.n6689 GND.n6688 9.3
R3432 GND.n6687 GND.n6686 9.3
R3433 GND.n6682 GND.n6681 9.3
R3434 GND.n6680 GND.n6679 9.3
R3435 GND.n6675 GND.n6674 9.3
R3436 GND.n6673 GND.n6672 9.3
R3437 GND.n6668 GND.n6667 9.3
R3438 GND.n6666 GND.n6665 9.3
R3439 GND.n6661 GND.n6660 9.3
R3440 GND.n6658 GND.n6657 9.3
R3441 GND.n6654 GND.n6653 9.3
R3442 GND.n6648 GND.n6647 9.3
R3443 GND.n6617 GND.n6616 9.3
R3444 GND.n6615 GND.n6614 9.3
R3445 GND.n6611 GND.n6610 9.3
R3446 GND.n6607 GND.n6606 9.3
R3447 GND.n6602 GND.n6601 9.3
R3448 GND.n6598 GND.n6597 9.3
R3449 GND.n6593 GND.n6592 9.3
R3450 GND.n6707 GND.n6706 9.3
R3451 GND.n6705 GND.n6704 9.3
R3452 GND.n6713 GND.n6712 9.3
R3453 GND.n6718 GND.n6717 9.3
R3454 GND.n6725 GND.n6724 9.3
R3455 GND.n6732 GND.n6731 9.3
R3456 GND.n6739 GND.n6738 9.3
R3457 GND.n6746 GND.n6745 9.3
R3458 GND.n6753 GND.n6752 9.3
R3459 GND.n6760 GND.n6759 9.3
R3460 GND.n6783 GND.n6782 9.3
R3461 GND.n6791 GND.n6790 9.3
R3462 GND.n6716 GND.n6715 9.3
R3463 GND.n6720 GND.n6719 9.3
R3464 GND.n6723 GND.n6722 9.3
R3465 GND.n6727 GND.n6726 9.3
R3466 GND.n6730 GND.n6729 9.3
R3467 GND.n6734 GND.n6733 9.3
R3468 GND.n6737 GND.n6736 9.3
R3469 GND.n6741 GND.n6740 9.3
R3470 GND.n6744 GND.n6743 9.3
R3471 GND.n6748 GND.n6747 9.3
R3472 GND.n6751 GND.n6750 9.3
R3473 GND.n6755 GND.n6754 9.3
R3474 GND.n6758 GND.n6757 9.3
R3475 GND.n6763 GND.n6762 9.3
R3476 GND.n6768 GND.n6767 9.3
R3477 GND.n6781 GND.n6780 9.3
R3478 GND.n6788 GND.n6787 9.3
R3479 GND.n6793 GND.n6792 9.3
R3480 GND.n6798 GND.n6797 9.3
R3481 GND.n6711 GND.n6710 9.3
R3482 GND.n6709 GND.n6708 9.3
R3483 GND.n6811 GND.n6810 9.3
R3484 GND.n6817 GND.n6816 9.3
R3485 GND.n6820 GND.n6819 9.3
R3486 GND.n6825 GND.n6824 9.3
R3487 GND.n6808 GND.n6807 9.3
R3488 GND.n6803 GND.n6802 9.3
R3489 GND.n6801 GND.n6800 9.3
R3490 GND.n7435 GND.n7434 9.3
R3491 GND.n7442 GND.n7441 9.3
R3492 GND.n7449 GND.n7448 9.3
R3493 GND.n7456 GND.n7455 9.3
R3494 GND.n7463 GND.n7462 9.3
R3495 GND.n7470 GND.n7469 9.3
R3496 GND.n7477 GND.n7476 9.3
R3497 GND.n7484 GND.n7483 9.3
R3498 GND.n6533 GND.n6532 9.3
R3499 GND.n6541 GND.n6540 9.3
R3500 GND.n6531 GND.n6530 9.3
R3501 GND.n6538 GND.n6537 9.3
R3502 GND.n6543 GND.n6542 9.3
R3503 GND.n6548 GND.n6547 9.3
R3504 GND.n7492 GND.n7491 9.3
R3505 GND.n7487 GND.n7486 9.3
R3506 GND.n7482 GND.n7481 9.3
R3507 GND.n7479 GND.n7478 9.3
R3508 GND.n7475 GND.n7474 9.3
R3509 GND.n7472 GND.n7471 9.3
R3510 GND.n7468 GND.n7467 9.3
R3511 GND.n7465 GND.n7464 9.3
R3512 GND.n7461 GND.n7460 9.3
R3513 GND.n7458 GND.n7457 9.3
R3514 GND.n7454 GND.n7453 9.3
R3515 GND.n7451 GND.n7450 9.3
R3516 GND.n7447 GND.n7446 9.3
R3517 GND.n7444 GND.n7443 9.3
R3518 GND.n7440 GND.n7439 9.3
R3519 GND.n7437 GND.n7436 9.3
R3520 GND.n7433 GND.n7432 9.3
R3521 GND.n6561 GND.n6560 9.3
R3522 GND.n6567 GND.n6566 9.3
R3523 GND.n6570 GND.n6569 9.3
R3524 GND.n6575 GND.n6574 9.3
R3525 GND.n6558 GND.n6557 9.3
R3526 GND.n6553 GND.n6552 9.3
R3527 GND.n6551 GND.n6550 9.3
R3528 GND.n7426 GND.n7425 9.3
R3529 GND.n7413 GND.n7412 9.3
R3530 GND.n7386 GND.n7385 9.3
R3531 GND.n7424 GND.n7423 9.3
R3532 GND.n7418 GND.n7417 9.3
R3533 GND.n7411 GND.n7410 9.3
R3534 GND.n7410 GND.n7409 9.3
R3535 GND.n7394 GND.n7393 9.3
R3536 GND.n7393 GND.n7392 9.3
R3537 GND.n7384 GND.n7383 9.3
R3538 GND.n7578 GND.n7577 9.3
R3539 GND.n7573 GND.n7572 9.3
R3540 GND.n7566 GND.n7565 9.3
R3541 GND.n7559 GND.n7558 9.3
R3542 GND.n7552 GND.n7551 9.3
R3543 GND.n7545 GND.n7544 9.3
R3544 GND.n7538 GND.n7537 9.3
R3545 GND.n7531 GND.n7530 9.3
R3546 GND.n7516 GND.n7515 9.3
R3547 GND.n6950 GND.n6949 9.3
R3548 GND.n7576 GND.n7575 9.3
R3549 GND.n7571 GND.n7570 9.3
R3550 GND.n7569 GND.n7568 9.3
R3551 GND.n7564 GND.n7563 9.3
R3552 GND.n7562 GND.n7561 9.3
R3553 GND.n7557 GND.n7556 9.3
R3554 GND.n7555 GND.n7554 9.3
R3555 GND.n7550 GND.n7549 9.3
R3556 GND.n7548 GND.n7547 9.3
R3557 GND.n7543 GND.n7542 9.3
R3558 GND.n7541 GND.n7540 9.3
R3559 GND.n7536 GND.n7535 9.3
R3560 GND.n7534 GND.n7533 9.3
R3561 GND.n7529 GND.n7528 9.3
R3562 GND.n7524 GND.n7523 9.3
R3563 GND.n7518 GND.n7517 9.3
R3564 GND.n6947 GND.n6946 9.3
R3565 GND.n6952 GND.n6951 9.3
R3566 GND.n6957 GND.n6956 9.3
R3567 GND.n7580 GND.n7579 9.3
R3568 GND.n7582 GND.n7581 9.3
R3569 GND.n6970 GND.n6969 9.3
R3570 GND.n6976 GND.n6975 9.3
R3571 GND.n6979 GND.n6978 9.3
R3572 GND.n6984 GND.n6983 9.3
R3573 GND.n6967 GND.n6966 9.3
R3574 GND.n6962 GND.n6961 9.3
R3575 GND.n6960 GND.n6959 9.3
R3576 GND.n7173 GND.n7172 9.3
R3577 GND.n7194 GND.n7193 9.3
R3578 GND.n7170 GND.n7169 9.3
R3579 GND.n7181 GND.n7180 9.3
R3580 GND.n7180 GND.n7179 9.3
R3581 GND.n7192 GND.n7191 9.3
R3582 GND.n7191 GND.n7190 9.3
R3583 GND.n7197 GND.n7196 9.3
R3584 GND.n7361 GND.n7360 9.3
R3585 GND.n7349 GND.n7348 9.3
R3586 GND.n7336 GND.n7335 9.3
R3587 GND.n7324 GND.n7323 9.3
R3588 GND.n7311 GND.n7310 9.3
R3589 GND.n7299 GND.n7298 9.3
R3590 GND.n7279 GND.n7278 9.3
R3591 GND.n7267 GND.n7266 9.3
R3592 GND.n7254 GND.n7253 9.3
R3593 GND.n7242 GND.n7241 9.3
R3594 GND.n7229 GND.n7228 9.3
R3595 GND.n7217 GND.n7216 9.3
R3596 GND.n7204 GND.n7203 9.3
R3597 GND.n7202 GND.n7201 9.3
R3598 GND.n7215 GND.n7214 9.3
R3599 GND.n7227 GND.n7226 9.3
R3600 GND.n7240 GND.n7239 9.3
R3601 GND.n7252 GND.n7251 9.3
R3602 GND.n7265 GND.n7264 9.3
R3603 GND.n7277 GND.n7276 9.3
R3604 GND.n7301 GND.n7300 9.3
R3605 GND.n7313 GND.n7312 9.3
R3606 GND.n7326 GND.n7325 9.3
R3607 GND.n7338 GND.n7337 9.3
R3608 GND.n7351 GND.n7350 9.3
R3609 GND.n7363 GND.n7362 9.3
R3610 GND.n7373 GND.n7372 9.3
R3611 GND.n7375 GND.n7374 9.3
R3612 GND.n7371 GND.n7370 9.3
R3613 GND.n7370 GND.n7369 9.3
R3614 GND.n6187 GND.n6186 9.3
R3615 GND.n6186 GND.n6185 9.3
R3616 GND.n6199 GND.n6198 9.3
R3617 GND.n6198 GND.n6197 9.3
R3618 GND.n6211 GND.n6210 9.3
R3619 GND.n6210 GND.n6209 9.3
R3620 GND.n6223 GND.n6222 9.3
R3621 GND.n6222 GND.n6221 9.3
R3622 GND.n6235 GND.n6234 9.3
R3623 GND.n6234 GND.n6233 9.3
R3624 GND.n6247 GND.n6246 9.3
R3625 GND.n6246 GND.n6245 9.3
R3626 GND.n6255 GND.n6254 9.3
R3627 GND.n6254 GND.n6253 9.3
R3628 GND.n6267 GND.n6266 9.3
R3629 GND.n6266 GND.n6265 9.3
R3630 GND.n6279 GND.n6278 9.3
R3631 GND.n6278 GND.n6277 9.3
R3632 GND.n6291 GND.n6290 9.3
R3633 GND.n6290 GND.n6289 9.3
R3634 GND.n6303 GND.n6302 9.3
R3635 GND.n6302 GND.n6301 9.3
R3636 GND.n6315 GND.n6314 9.3
R3637 GND.n6314 GND.n6313 9.3
R3638 GND.n6327 GND.n6326 9.3
R3639 GND.n6326 GND.n6325 9.3
R3640 GND.n7213 GND.n7212 9.3
R3641 GND.n7212 GND.n7211 9.3
R3642 GND.n7211 GND.n7210 9.3
R3643 GND.n7225 GND.n7224 9.3
R3644 GND.n7224 GND.n7223 9.3
R3645 GND.n7238 GND.n7237 9.3
R3646 GND.n7237 GND.n7236 9.3
R3647 GND.n7250 GND.n7249 9.3
R3648 GND.n7249 GND.n7248 9.3
R3649 GND.n7263 GND.n7262 9.3
R3650 GND.n7262 GND.n7261 9.3
R3651 GND.n7275 GND.n7274 9.3
R3652 GND.n7274 GND.n7273 9.3
R3653 GND.n7288 GND.n7287 9.3
R3654 GND.n7287 GND.n7286 9.3
R3655 GND.n7297 GND.n7296 9.3
R3656 GND.n7296 GND.n7295 9.3
R3657 GND.n7309 GND.n7308 9.3
R3658 GND.n7308 GND.n7307 9.3
R3659 GND.n7322 GND.n7321 9.3
R3660 GND.n7321 GND.n7320 9.3
R3661 GND.n7334 GND.n7333 9.3
R3662 GND.n7333 GND.n7332 9.3
R3663 GND.n7347 GND.n7346 9.3
R3664 GND.n7346 GND.n7345 9.3
R3665 GND.n7359 GND.n7358 9.3
R3666 GND.n7358 GND.n7357 9.3
R3667 GND.n6174 GND.n6173 9.3
R3668 GND.n6173 GND.n6172 9.3
R3669 GND.n11308 GND.n11307 9.3
R3670 GND.n11307 GND.n11306 9.3
R3671 GND.n11296 GND.n11295 9.3
R3672 GND.n11295 GND.n11294 9.3
R3673 GND.n11284 GND.n11283 9.3
R3674 GND.n11283 GND.n11282 9.3
R3675 GND.n11272 GND.n11271 9.3
R3676 GND.n11271 GND.n11270 9.3
R3677 GND.n11260 GND.n11259 9.3
R3678 GND.n11259 GND.n11258 9.3
R3679 GND.n11248 GND.n11247 9.3
R3680 GND.n11247 GND.n11246 9.3
R3681 GND.n11236 GND.n11235 9.3
R3682 GND.n11235 GND.n11234 9.3
R3683 GND.n11228 GND.n11227 9.3
R3684 GND.n11227 GND.n11226 9.3
R3685 GND.n11216 GND.n11215 9.3
R3686 GND.n11215 GND.n11214 9.3
R3687 GND.n11204 GND.n11203 9.3
R3688 GND.n11203 GND.n11202 9.3
R3689 GND.n11192 GND.n11191 9.3
R3690 GND.n11191 GND.n11190 9.3
R3691 GND.n11180 GND.n11179 9.3
R3692 GND.n11179 GND.n11178 9.3
R3693 GND.n11168 GND.n11167 9.3
R3694 GND.n11167 GND.n11166 9.3
R3695 GND.n11156 GND.n11155 9.3
R3696 GND.n11155 GND.n11154 9.3
R3697 GND.n11154 GND.n11153 9.3
R3698 GND.n13563 GND.n13562 9.3
R3699 GND.n13562 GND.n13561 9.3
R3700 GND.n13561 GND.n13560 9.3
R3701 GND.n13575 GND.n13574 9.3
R3702 GND.n13574 GND.n13573 9.3
R3703 GND.n13587 GND.n13586 9.3
R3704 GND.n13586 GND.n13585 9.3
R3705 GND.n13599 GND.n13598 9.3
R3706 GND.n13598 GND.n13597 9.3
R3707 GND.n13611 GND.n13610 9.3
R3708 GND.n13610 GND.n13609 9.3
R3709 GND.n13623 GND.n13622 9.3
R3710 GND.n13622 GND.n13621 9.3
R3711 GND.n13635 GND.n13634 9.3
R3712 GND.n13634 GND.n13633 9.3
R3713 GND.n13643 GND.n13642 9.3
R3714 GND.n13642 GND.n13641 9.3
R3715 GND.n13655 GND.n13654 9.3
R3716 GND.n13654 GND.n13653 9.3
R3717 GND.n13667 GND.n13666 9.3
R3718 GND.n13666 GND.n13665 9.3
R3719 GND.n13679 GND.n13678 9.3
R3720 GND.n13678 GND.n13677 9.3
R3721 GND.n13691 GND.n13690 9.3
R3722 GND.n13690 GND.n13689 9.3
R3723 GND.n13703 GND.n13702 9.3
R3724 GND.n13702 GND.n13701 9.3
R3725 GND.n13715 GND.n13714 9.3
R3726 GND.n13714 GND.n13713 9.3
R3727 GND.n15939 GND.n15938 9.3
R3728 GND.n15938 GND.n15937 9.3
R3729 GND.n15937 GND.n15936 9.3
R3730 GND.n15943 GND.n15942 9.3
R3731 GND.n15955 GND.n15954 9.3
R3732 GND.n15968 GND.n15967 9.3
R3733 GND.n15980 GND.n15979 9.3
R3734 GND.n15993 GND.n15992 9.3
R3735 GND.n16015 GND.n16014 9.3
R3736 GND.n16023 GND.n16022 9.3
R3737 GND.n16031 GND.n16030 9.3
R3738 GND.n16039 GND.n16038 9.3
R3739 GND.n16047 GND.n16046 9.3
R3740 GND.n16055 GND.n16054 9.3
R3741 GND.n16063 GND.n16062 9.3
R3742 GND.n16069 GND.n16068 9.3
R3743 GND.n16074 GND.n16073 9.3
R3744 GND.n16079 GND.n16078 9.3
R3745 GND.n16098 GND.n16097 9.3
R3746 GND.n16116 GND.n16115 9.3
R3747 GND.n16128 GND.n16127 9.3
R3748 GND.n16140 GND.n16139 9.3
R3749 GND.n16152 GND.n16151 9.3
R3750 GND.n16164 GND.n16163 9.3
R3751 GND.n16177 GND.n16176 9.3
R3752 GND.n16179 GND.n16178 9.3
R3753 GND.n16166 GND.n16165 9.3
R3754 GND.n16154 GND.n16153 9.3
R3755 GND.n16142 GND.n16141 9.3
R3756 GND.n16130 GND.n16129 9.3
R3757 GND.n16118 GND.n16117 9.3
R3758 GND.n16096 GND.n16095 9.3
R3759 GND.n16086 GND.n16085 9.3
R3760 GND.n16082 GND.n16081 9.3
R3761 GND.n16077 GND.n16076 9.3
R3762 GND.n16072 GND.n16071 9.3
R3763 GND.n16067 GND.n16066 9.3
R3764 GND.n16065 GND.n16064 9.3
R3765 GND.n16061 GND.n16060 9.3
R3766 GND.n15936 GND.n15935 9.3
R3767 GND.n16057 GND.n16056 9.3
R3768 GND.n16053 GND.n16052 9.3
R3769 GND.n16049 GND.n16048 9.3
R3770 GND.n16045 GND.n16044 9.3
R3771 GND.n16041 GND.n16040 9.3
R3772 GND.n16037 GND.n16036 9.3
R3773 GND.n16033 GND.n16032 9.3
R3774 GND.n16029 GND.n16028 9.3
R3775 GND.n16025 GND.n16024 9.3
R3776 GND.n16021 GND.n16020 9.3
R3777 GND.n16017 GND.n16016 9.3
R3778 GND.n16013 GND.n16012 9.3
R3779 GND.n16006 GND.n16005 9.3
R3780 GND.n16005 GND.n16004 9.3
R3781 GND.n15991 GND.n15990 9.3
R3782 GND.n15989 GND.n15988 9.3
R3783 GND.n15988 GND.n15987 9.3
R3784 GND.n15978 GND.n15977 9.3
R3785 GND.n15976 GND.n15975 9.3
R3786 GND.n15975 GND.n15974 9.3
R3787 GND.n15966 GND.n15965 9.3
R3788 GND.n15964 GND.n15963 9.3
R3789 GND.n15963 GND.n15962 9.3
R3790 GND.n15953 GND.n15952 9.3
R3791 GND.n15951 GND.n15950 9.3
R3792 GND.n15950 GND.n15949 9.3
R3793 GND.n15941 GND.n15940 9.3
R3794 GND.n16232 GND.n16231 9.3
R3795 GND.n16230 GND.n16229 9.3
R3796 GND.n15894 GND.n15893 9.3
R3797 GND.n15892 GND.n15891 9.3
R3798 GND.n16175 GND.n16174 9.3
R3799 GND.n16174 GND.n16173 9.3
R3800 GND.n16162 GND.n16161 9.3
R3801 GND.n16161 GND.n16160 9.3
R3802 GND.n16150 GND.n16149 9.3
R3803 GND.n16149 GND.n16148 9.3
R3804 GND.n16138 GND.n16137 9.3
R3805 GND.n16137 GND.n16136 9.3
R3806 GND.n16126 GND.n16125 9.3
R3807 GND.n16125 GND.n16124 9.3
R3808 GND.n16114 GND.n16113 9.3
R3809 GND.n16113 GND.n16112 9.3
R3810 GND.n16106 GND.n16105 9.3
R3811 GND.n16105 GND.n16104 9.3
R3812 GND.n16092 GND.n16091 9.3
R3813 GND.n16201 GND.n16200 9.3
R3814 GND.n16213 GND.n16212 9.3
R3815 GND.n16194 GND.n16193 9.3
R3816 GND.n16220 GND.n16219 9.3
R3817 GND.n16187 GND.n16186 9.3
R3818 GND.n16228 GND.n16227 9.3
R3819 GND.n16227 GND.n16226 9.3
R3820 GND.n1168 GND.n1167 9.3
R3821 GND.n1167 GND.n1166 9.3
R3822 GND.n1166 GND.n1165 9.3
R3823 GND.n1125 GND.n1124 9.3
R3824 GND.n1113 GND.n1112 9.3
R3825 GND.n1101 GND.n1100 9.3
R3826 GND.n1089 GND.n1088 9.3
R3827 GND.n1077 GND.n1076 9.3
R3828 GND.n1055 GND.n1054 9.3
R3829 GND.n1047 GND.n1046 9.3
R3830 GND.n1039 GND.n1038 9.3
R3831 GND.n1031 GND.n1030 9.3
R3832 GND.n1023 GND.n1022 9.3
R3833 GND.n1015 GND.n1014 9.3
R3834 GND.n1007 GND.n1006 9.3
R3835 GND.n1001 GND.n1000 9.3
R3836 GND.n996 GND.n995 9.3
R3837 GND.n991 GND.n990 9.3
R3838 GND.n972 GND.n971 9.3
R3839 GND.n953 GND.n952 9.3
R3840 GND.n940 GND.n939 9.3
R3841 GND.n928 GND.n927 9.3
R3842 GND.n915 GND.n914 9.3
R3843 GND.n903 GND.n902 9.3
R3844 GND.n890 GND.n889 9.3
R3845 GND.n888 GND.n887 9.3
R3846 GND.n899 GND.n898 9.3
R3847 GND.n898 GND.n897 9.3
R3848 GND.n901 GND.n900 9.3
R3849 GND.n911 GND.n910 9.3
R3850 GND.n910 GND.n909 9.3
R3851 GND.n913 GND.n912 9.3
R3852 GND.n924 GND.n923 9.3
R3853 GND.n923 GND.n922 9.3
R3854 GND.n926 GND.n925 9.3
R3855 GND.n936 GND.n935 9.3
R3856 GND.n935 GND.n934 9.3
R3857 GND.n938 GND.n937 9.3
R3858 GND.n949 GND.n948 9.3
R3859 GND.n948 GND.n947 9.3
R3860 GND.n951 GND.n950 9.3
R3861 GND.n962 GND.n961 9.3
R3862 GND.n961 GND.n960 9.3
R3863 GND.n970 GND.n969 9.3
R3864 GND.n969 GND.n968 9.3
R3865 GND.n974 GND.n973 9.3
R3866 GND.n978 GND.n977 9.3
R3867 GND.n873 GND.n872 9.3
R3868 GND.n984 GND.n983 9.3
R3869 GND.n868 GND.n867 9.3
R3870 GND.n988 GND.n987 9.3
R3871 GND.n857 GND.n856 9.3
R3872 GND.n993 GND.n992 9.3
R3873 GND.n852 GND.n851 9.3
R3874 GND.n998 GND.n997 9.3
R3875 GND.n842 GND.n841 9.3
R3876 GND.n1003 GND.n1002 9.3
R3877 GND.n1005 GND.n1004 9.3
R3878 GND.n1011 GND.n1010 9.3
R3879 GND.n1165 GND.n1152 9.3
R3880 GND.n1013 GND.n1012 9.3
R3881 GND.n1019 GND.n1018 9.3
R3882 GND.n1165 GND.n1156 9.3
R3883 GND.n1021 GND.n1020 9.3
R3884 GND.n1027 GND.n1026 9.3
R3885 GND.n1165 GND.n1148 9.3
R3886 GND.n1029 GND.n1028 9.3
R3887 GND.n1035 GND.n1034 9.3
R3888 GND.n1165 GND.n1160 9.3
R3889 GND.n1037 GND.n1036 9.3
R3890 GND.n1043 GND.n1042 9.3
R3891 GND.n1165 GND.n1144 9.3
R3892 GND.n1045 GND.n1044 9.3
R3893 GND.n1051 GND.n1050 9.3
R3894 GND.n1165 GND.n1164 9.3
R3895 GND.n1053 GND.n1052 9.3
R3896 GND.n1059 GND.n1058 9.3
R3897 GND.n1165 GND.n1140 9.3
R3898 GND.n1075 GND.n1074 9.3
R3899 GND.n1074 GND.n1073 9.3
R3900 GND.n1079 GND.n1078 9.3
R3901 GND.n1087 GND.n1086 9.3
R3902 GND.n1086 GND.n1085 9.3
R3903 GND.n1091 GND.n1090 9.3
R3904 GND.n1099 GND.n1098 9.3
R3905 GND.n1098 GND.n1097 9.3
R3906 GND.n1103 GND.n1102 9.3
R3907 GND.n1111 GND.n1110 9.3
R3908 GND.n1110 GND.n1109 9.3
R3909 GND.n1115 GND.n1114 9.3
R3910 GND.n1123 GND.n1122 9.3
R3911 GND.n1122 GND.n1121 9.3
R3912 GND.n1127 GND.n1126 9.3
R3913 GND.n886 GND.n885 9.3
R3914 GND.n885 GND.n884 9.3
R3915 GND.n832 GND.n831 9.3
R3916 GND.n834 GND.n833 9.3
R3917 GND.n1170 GND.n1169 9.3
R3918 GND.n1172 GND.n1171 9.3
R3919 GND.n9639 GND.n9638 9.3
R3920 GND.n9638 GND.n9637 9.3
R3921 GND.n9637 GND.n9636 9.3
R3922 GND.n9643 GND.n9642 9.3
R3923 GND.n9655 GND.n9654 9.3
R3924 GND.n9668 GND.n9667 9.3
R3925 GND.n9680 GND.n9679 9.3
R3926 GND.n9693 GND.n9692 9.3
R3927 GND.n9715 GND.n9714 9.3
R3928 GND.n9723 GND.n9722 9.3
R3929 GND.n9731 GND.n9730 9.3
R3930 GND.n9739 GND.n9738 9.3
R3931 GND.n9747 GND.n9746 9.3
R3932 GND.n9755 GND.n9754 9.3
R3933 GND.n9763 GND.n9762 9.3
R3934 GND.n9769 GND.n9768 9.3
R3935 GND.n9774 GND.n9773 9.3
R3936 GND.n9779 GND.n9778 9.3
R3937 GND.n9798 GND.n9797 9.3
R3938 GND.n9816 GND.n9815 9.3
R3939 GND.n9828 GND.n9827 9.3
R3940 GND.n9840 GND.n9839 9.3
R3941 GND.n9852 GND.n9851 9.3
R3942 GND.n9864 GND.n9863 9.3
R3943 GND.n9877 GND.n9876 9.3
R3944 GND.n9879 GND.n9878 9.3
R3945 GND.n9866 GND.n9865 9.3
R3946 GND.n9854 GND.n9853 9.3
R3947 GND.n9842 GND.n9841 9.3
R3948 GND.n9830 GND.n9829 9.3
R3949 GND.n9818 GND.n9817 9.3
R3950 GND.n9796 GND.n9795 9.3
R3951 GND.n9786 GND.n9785 9.3
R3952 GND.n9782 GND.n9781 9.3
R3953 GND.n9777 GND.n9776 9.3
R3954 GND.n9772 GND.n9771 9.3
R3955 GND.n9767 GND.n9766 9.3
R3956 GND.n9765 GND.n9764 9.3
R3957 GND.n9761 GND.n9760 9.3
R3958 GND.n9636 GND.n9635 9.3
R3959 GND.n9757 GND.n9756 9.3
R3960 GND.n9753 GND.n9752 9.3
R3961 GND.n9749 GND.n9748 9.3
R3962 GND.n9745 GND.n9744 9.3
R3963 GND.n9741 GND.n9740 9.3
R3964 GND.n9737 GND.n9736 9.3
R3965 GND.n9733 GND.n9732 9.3
R3966 GND.n9729 GND.n9728 9.3
R3967 GND.n9725 GND.n9724 9.3
R3968 GND.n9721 GND.n9720 9.3
R3969 GND.n9717 GND.n9716 9.3
R3970 GND.n9713 GND.n9712 9.3
R3971 GND.n9706 GND.n9705 9.3
R3972 GND.n9705 GND.n9704 9.3
R3973 GND.n9691 GND.n9690 9.3
R3974 GND.n9689 GND.n9688 9.3
R3975 GND.n9688 GND.n9687 9.3
R3976 GND.n9678 GND.n9677 9.3
R3977 GND.n9676 GND.n9675 9.3
R3978 GND.n9675 GND.n9674 9.3
R3979 GND.n9666 GND.n9665 9.3
R3980 GND.n9664 GND.n9663 9.3
R3981 GND.n9663 GND.n9662 9.3
R3982 GND.n9653 GND.n9652 9.3
R3983 GND.n9651 GND.n9650 9.3
R3984 GND.n9650 GND.n9649 9.3
R3985 GND.n9641 GND.n9640 9.3
R3986 GND.n9932 GND.n9931 9.3
R3987 GND.n9930 GND.n9929 9.3
R3988 GND.n9594 GND.n9593 9.3
R3989 GND.n1174 GND.n1173 9.3
R3990 GND.n9875 GND.n9874 9.3
R3991 GND.n9874 GND.n9873 9.3
R3992 GND.n9862 GND.n9861 9.3
R3993 GND.n9861 GND.n9860 9.3
R3994 GND.n9850 GND.n9849 9.3
R3995 GND.n9849 GND.n9848 9.3
R3996 GND.n9838 GND.n9837 9.3
R3997 GND.n9837 GND.n9836 9.3
R3998 GND.n9826 GND.n9825 9.3
R3999 GND.n9825 GND.n9824 9.3
R4000 GND.n9814 GND.n9813 9.3
R4001 GND.n9813 GND.n9812 9.3
R4002 GND.n9806 GND.n9805 9.3
R4003 GND.n9805 GND.n9804 9.3
R4004 GND.n9792 GND.n9791 9.3
R4005 GND.n9901 GND.n9900 9.3
R4006 GND.n9913 GND.n9912 9.3
R4007 GND.n9894 GND.n9893 9.3
R4008 GND.n9920 GND.n9919 9.3
R4009 GND.n9887 GND.n9886 9.3
R4010 GND.n9928 GND.n9927 9.3
R4011 GND.n9927 GND.n9926 9.3
R4012 GND.n1231 GND.n1230 9.3
R4013 GND.n1230 GND.n1229 9.3
R4014 GND.n1229 GND.n1228 9.3
R4015 GND.n1235 GND.n1234 9.3
R4016 GND.n1247 GND.n1246 9.3
R4017 GND.n1259 GND.n1258 9.3
R4018 GND.n1271 GND.n1270 9.3
R4019 GND.n1283 GND.n1282 9.3
R4020 GND.n1305 GND.n1304 9.3
R4021 GND.n1313 GND.n1312 9.3
R4022 GND.n1321 GND.n1320 9.3
R4023 GND.n1329 GND.n1328 9.3
R4024 GND.n1337 GND.n1336 9.3
R4025 GND.n1345 GND.n1344 9.3
R4026 GND.n1353 GND.n1352 9.3
R4027 GND.n1359 GND.n1358 9.3
R4028 GND.n1364 GND.n1363 9.3
R4029 GND.n1369 GND.n1368 9.3
R4030 GND.n1388 GND.n1387 9.3
R4031 GND.n1407 GND.n1406 9.3
R4032 GND.n1420 GND.n1419 9.3
R4033 GND.n1432 GND.n1431 9.3
R4034 GND.n1445 GND.n1444 9.3
R4035 GND.n1457 GND.n1456 9.3
R4036 GND.n1470 GND.n1469 9.3
R4037 GND.n1472 GND.n1471 9.3
R4038 GND.n1468 GND.n1467 9.3
R4039 GND.n1467 GND.n1466 9.3
R4040 GND.n1459 GND.n1458 9.3
R4041 GND.n1455 GND.n1454 9.3
R4042 GND.n1454 GND.n1453 9.3
R4043 GND.n1447 GND.n1446 9.3
R4044 GND.n1443 GND.n1442 9.3
R4045 GND.n1442 GND.n1441 9.3
R4046 GND.n1434 GND.n1433 9.3
R4047 GND.n1430 GND.n1429 9.3
R4048 GND.n1429 GND.n1428 9.3
R4049 GND.n1422 GND.n1421 9.3
R4050 GND.n1418 GND.n1417 9.3
R4051 GND.n1417 GND.n1416 9.3
R4052 GND.n1409 GND.n1408 9.3
R4053 GND.n1405 GND.n1404 9.3
R4054 GND.n1404 GND.n1403 9.3
R4055 GND.n1396 GND.n1395 9.3
R4056 GND.n1395 GND.n1394 9.3
R4057 GND.n1386 GND.n1385 9.3
R4058 GND.n1382 GND.n1381 9.3
R4059 GND.n1511 GND.n1510 9.3
R4060 GND.n1376 GND.n1375 9.3
R4061 GND.n1506 GND.n1505 9.3
R4062 GND.n1372 GND.n1371 9.3
R4063 GND.n1495 GND.n1494 9.3
R4064 GND.n1367 GND.n1366 9.3
R4065 GND.n1490 GND.n1489 9.3
R4066 GND.n1362 GND.n1361 9.3
R4067 GND.n1480 GND.n1479 9.3
R4068 GND.n1357 GND.n1356 9.3
R4069 GND.n1355 GND.n1354 9.3
R4070 GND.n1351 GND.n1350 9.3
R4071 GND.n1228 GND.n1215 9.3
R4072 GND.n1347 GND.n1346 9.3
R4073 GND.n1343 GND.n1342 9.3
R4074 GND.n1228 GND.n1219 9.3
R4075 GND.n1339 GND.n1338 9.3
R4076 GND.n1335 GND.n1334 9.3
R4077 GND.n1228 GND.n1211 9.3
R4078 GND.n1331 GND.n1330 9.3
R4079 GND.n1327 GND.n1326 9.3
R4080 GND.n1228 GND.n1223 9.3
R4081 GND.n1323 GND.n1322 9.3
R4082 GND.n1319 GND.n1318 9.3
R4083 GND.n1228 GND.n1207 9.3
R4084 GND.n1315 GND.n1314 9.3
R4085 GND.n1311 GND.n1310 9.3
R4086 GND.n1228 GND.n1227 9.3
R4087 GND.n1307 GND.n1306 9.3
R4088 GND.n1303 GND.n1302 9.3
R4089 GND.n1228 GND.n1203 9.3
R4090 GND.n1296 GND.n1295 9.3
R4091 GND.n1295 GND.n1294 9.3
R4092 GND.n1281 GND.n1280 9.3
R4093 GND.n1279 GND.n1278 9.3
R4094 GND.n1278 GND.n1277 9.3
R4095 GND.n1269 GND.n1268 9.3
R4096 GND.n1267 GND.n1266 9.3
R4097 GND.n1266 GND.n1265 9.3
R4098 GND.n1257 GND.n1256 9.3
R4099 GND.n1255 GND.n1254 9.3
R4100 GND.n1254 GND.n1253 9.3
R4101 GND.n1245 GND.n1244 9.3
R4102 GND.n1243 GND.n1242 9.3
R4103 GND.n1242 GND.n1241 9.3
R4104 GND.n1233 GND.n1232 9.3
R4105 GND.n1524 GND.n1523 9.3
R4106 GND.n1523 GND.n1522 9.3
R4107 GND.n1528 GND.n1527 9.3
R4108 GND.n1526 GND.n1525 9.3
R4109 GND.n1190 GND.n1189 9.3
R4110 GND.n1176 GND.n1175 9.3
R4111 GND.n10305 GND.n10304 9.3
R4112 GND.n10304 GND.n10303 9.3
R4113 GND.n10295 GND.n10294 9.3
R4114 GND.n10283 GND.n10282 9.3
R4115 GND.n10270 GND.n10269 9.3
R4116 GND.n10258 GND.n10257 9.3
R4117 GND.n10245 GND.n10244 9.3
R4118 GND.n10233 GND.n10232 9.3
R4119 GND.n10213 GND.n10212 9.3
R4120 GND.n10201 GND.n10200 9.3
R4121 GND.n10188 GND.n10187 9.3
R4122 GND.n10176 GND.n10175 9.3
R4123 GND.n10163 GND.n10162 9.3
R4124 GND.n10151 GND.n10150 9.3
R4125 GND.n10147 GND.n10146 9.3
R4126 GND.n10146 GND.n10145 9.3
R4127 GND.n10145 GND.n10144 9.3
R4128 GND.n10149 GND.n10148 9.3
R4129 GND.n10159 GND.n10158 9.3
R4130 GND.n10158 GND.n10157 9.3
R4131 GND.n10161 GND.n10160 9.3
R4132 GND.n10172 GND.n10171 9.3
R4133 GND.n10171 GND.n10170 9.3
R4134 GND.n10174 GND.n10173 9.3
R4135 GND.n10184 GND.n10183 9.3
R4136 GND.n10183 GND.n10182 9.3
R4137 GND.n10186 GND.n10185 9.3
R4138 GND.n10197 GND.n10196 9.3
R4139 GND.n10196 GND.n10195 9.3
R4140 GND.n10199 GND.n10198 9.3
R4141 GND.n10209 GND.n10208 9.3
R4142 GND.n10208 GND.n10207 9.3
R4143 GND.n10211 GND.n10210 9.3
R4144 GND.n10222 GND.n10221 9.3
R4145 GND.n10221 GND.n10220 9.3
R4146 GND.n10231 GND.n10230 9.3
R4147 GND.n10230 GND.n10229 9.3
R4148 GND.n10235 GND.n10234 9.3
R4149 GND.n10243 GND.n10242 9.3
R4150 GND.n10242 GND.n10241 9.3
R4151 GND.n10247 GND.n10246 9.3
R4152 GND.n10256 GND.n10255 9.3
R4153 GND.n10255 GND.n10254 9.3
R4154 GND.n10260 GND.n10259 9.3
R4155 GND.n10268 GND.n10267 9.3
R4156 GND.n10267 GND.n10266 9.3
R4157 GND.n10272 GND.n10271 9.3
R4158 GND.n10281 GND.n10280 9.3
R4159 GND.n10280 GND.n10279 9.3
R4160 GND.n10285 GND.n10284 9.3
R4161 GND.n10293 GND.n10292 9.3
R4162 GND.n10292 GND.n10291 9.3
R4163 GND.n10297 GND.n10296 9.3
R4164 GND.n10136 GND.n10135 9.3
R4165 GND.n10138 GND.n10137 9.3
R4166 GND.n10307 GND.n10306 9.3
R4167 GND.n10309 GND.n10308 9.3
R4168 GND.n8868 GND.n8867 9.3
R4169 GND.n8867 GND.n8866 9.3
R4170 GND.n8858 GND.n8857 9.3
R4171 GND.n8846 GND.n8845 9.3
R4172 GND.n8834 GND.n8833 9.3
R4173 GND.n8822 GND.n8821 9.3
R4174 GND.n8810 GND.n8809 9.3
R4175 GND.n8798 GND.n8797 9.3
R4176 GND.n8780 GND.n8779 9.3
R4177 GND.n8768 GND.n8767 9.3
R4178 GND.n8756 GND.n8755 9.3
R4179 GND.n8744 GND.n8743 9.3
R4180 GND.n8732 GND.n8731 9.3
R4181 GND.n8720 GND.n8719 9.3
R4182 GND.n8716 GND.n8715 9.3
R4183 GND.n8715 GND.n8714 9.3
R4184 GND.n8714 GND.n8713 9.3
R4185 GND.n8718 GND.n8717 9.3
R4186 GND.n8728 GND.n8727 9.3
R4187 GND.n8727 GND.n8726 9.3
R4188 GND.n8730 GND.n8729 9.3
R4189 GND.n8740 GND.n8739 9.3
R4190 GND.n8739 GND.n8738 9.3
R4191 GND.n8742 GND.n8741 9.3
R4192 GND.n8752 GND.n8751 9.3
R4193 GND.n8751 GND.n8750 9.3
R4194 GND.n8754 GND.n8753 9.3
R4195 GND.n8764 GND.n8763 9.3
R4196 GND.n8763 GND.n8762 9.3
R4197 GND.n8766 GND.n8765 9.3
R4198 GND.n8776 GND.n8775 9.3
R4199 GND.n8775 GND.n8774 9.3
R4200 GND.n8778 GND.n8777 9.3
R4201 GND.n8788 GND.n8787 9.3
R4202 GND.n8787 GND.n8786 9.3
R4203 GND.n8796 GND.n8795 9.3
R4204 GND.n8795 GND.n8794 9.3
R4205 GND.n8800 GND.n8799 9.3
R4206 GND.n8808 GND.n8807 9.3
R4207 GND.n8807 GND.n8806 9.3
R4208 GND.n8812 GND.n8811 9.3
R4209 GND.n8820 GND.n8819 9.3
R4210 GND.n8819 GND.n8818 9.3
R4211 GND.n8824 GND.n8823 9.3
R4212 GND.n8832 GND.n8831 9.3
R4213 GND.n8831 GND.n8830 9.3
R4214 GND.n8836 GND.n8835 9.3
R4215 GND.n8844 GND.n8843 9.3
R4216 GND.n8843 GND.n8842 9.3
R4217 GND.n8848 GND.n8847 9.3
R4218 GND.n8856 GND.n8855 9.3
R4219 GND.n8855 GND.n8854 9.3
R4220 GND.n8860 GND.n8859 9.3
R4221 GND.n8705 GND.n8704 9.3
R4222 GND.n8707 GND.n8706 9.3
R4223 GND.n8870 GND.n8869 9.3
R4224 GND.n8872 GND.n8871 9.3
R4225 GND.n8577 GND.n8576 9.3
R4226 GND.n8565 GND.n8564 9.3
R4227 GND.n8553 GND.n8552 9.3
R4228 GND.n8540 GND.n8539 9.3
R4229 GND.n8528 GND.n8527 9.3
R4230 GND.n8515 GND.n8514 9.3
R4231 GND.n8503 GND.n8502 9.3
R4232 GND.n8483 GND.n8482 9.3
R4233 GND.n8471 GND.n8470 9.3
R4234 GND.n8458 GND.n8457 9.3
R4235 GND.n8446 GND.n8445 9.3
R4236 GND.n8433 GND.n8432 9.3
R4237 GND.n8421 GND.n8420 9.3
R4238 GND.n8417 GND.n8416 9.3
R4239 GND.n8416 GND.n8415 9.3
R4240 GND.n8415 GND.n8414 9.3
R4241 GND.n8567 GND.n8566 9.3
R4242 GND.n8563 GND.n8562 9.3
R4243 GND.n8562 GND.n8561 9.3
R4244 GND.n8555 GND.n8554 9.3
R4245 GND.n8551 GND.n8550 9.3
R4246 GND.n8550 GND.n8549 9.3
R4247 GND.n8542 GND.n8541 9.3
R4248 GND.n8538 GND.n8537 9.3
R4249 GND.n8537 GND.n8536 9.3
R4250 GND.n8530 GND.n8529 9.3
R4251 GND.n8526 GND.n8525 9.3
R4252 GND.n8525 GND.n8524 9.3
R4253 GND.n8517 GND.n8516 9.3
R4254 GND.n8513 GND.n8512 9.3
R4255 GND.n8512 GND.n8511 9.3
R4256 GND.n8505 GND.n8504 9.3
R4257 GND.n8501 GND.n8500 9.3
R4258 GND.n8500 GND.n8499 9.3
R4259 GND.n8492 GND.n8491 9.3
R4260 GND.n8491 GND.n8490 9.3
R4261 GND.n8481 GND.n8480 9.3
R4262 GND.n8479 GND.n8478 9.3
R4263 GND.n8478 GND.n8477 9.3
R4264 GND.n8469 GND.n8468 9.3
R4265 GND.n8467 GND.n8466 9.3
R4266 GND.n8466 GND.n8465 9.3
R4267 GND.n8456 GND.n8455 9.3
R4268 GND.n8454 GND.n8453 9.3
R4269 GND.n8453 GND.n8452 9.3
R4270 GND.n8444 GND.n8443 9.3
R4271 GND.n8442 GND.n8441 9.3
R4272 GND.n8441 GND.n8440 9.3
R4273 GND.n8431 GND.n8430 9.3
R4274 GND.n8419 GND.n8418 9.3
R4275 GND.n8429 GND.n8428 9.3
R4276 GND.n8428 GND.n8427 9.3
R4277 GND.n8575 GND.n8574 9.3
R4278 GND.n8574 GND.n8573 9.3
R4279 GND.n8579 GND.n8578 9.3
R4280 GND.n1899 GND.n1898 9.3
R4281 GND.n8408 GND.n8407 9.3
R4282 GND.n9296 GND.n9295 9.3
R4283 GND.n9303 GND.n9302 9.3
R4284 GND.n9310 GND.n9309 9.3
R4285 GND.n9317 GND.n9316 9.3
R4286 GND.n9324 GND.n9323 9.3
R4287 GND.n9331 GND.n9330 9.3
R4288 GND.n9338 GND.n9337 9.3
R4289 GND.n9345 GND.n9344 9.3
R4290 GND.n9366 GND.n9365 9.3
R4291 GND.n9374 GND.n9373 9.3
R4292 GND.n9384 GND.n9383 9.3
R4293 GND.n9403 GND.n9402 9.3
R4294 GND.n9400 GND.n9399 9.3
R4295 GND.n9394 GND.n9393 9.3
R4296 GND.n9391 GND.n9390 9.3
R4297 GND.n9386 GND.n9385 9.3
R4298 GND.n9381 GND.n9380 9.3
R4299 GND.n9376 GND.n9375 9.3
R4300 GND.n9371 GND.n9370 9.3
R4301 GND.n9364 GND.n9363 9.3
R4302 GND.n9353 GND.n9352 9.3
R4303 GND.n9348 GND.n9347 9.3
R4304 GND.n9343 GND.n9342 9.3
R4305 GND.n9340 GND.n9339 9.3
R4306 GND.n9336 GND.n9335 9.3
R4307 GND.n9333 GND.n9332 9.3
R4308 GND.n9329 GND.n9328 9.3
R4309 GND.n9326 GND.n9325 9.3
R4310 GND.n9322 GND.n9321 9.3
R4311 GND.n9319 GND.n9318 9.3
R4312 GND.n9315 GND.n9314 9.3
R4313 GND.n9312 GND.n9311 9.3
R4314 GND.n9308 GND.n9307 9.3
R4315 GND.n9305 GND.n9304 9.3
R4316 GND.n9301 GND.n9300 9.3
R4317 GND.n9298 GND.n9297 9.3
R4318 GND.n9294 GND.n9293 9.3
R4319 GND.n9407 GND.n9406 9.3
R4320 GND.n1701 GND.n1700 9.3
R4321 GND.n1708 GND.n1707 9.3
R4322 GND.n1715 GND.n1714 9.3
R4323 GND.n1722 GND.n1721 9.3
R4324 GND.n1729 GND.n1728 9.3
R4325 GND.n1736 GND.n1735 9.3
R4326 GND.n1743 GND.n1742 9.3
R4327 GND.n1750 GND.n1749 9.3
R4328 GND.n1773 GND.n1772 9.3
R4329 GND.n1781 GND.n1780 9.3
R4330 GND.n1791 GND.n1790 9.3
R4331 GND.n1810 GND.n1809 9.3
R4332 GND.n1807 GND.n1806 9.3
R4333 GND.n1801 GND.n1800 9.3
R4334 GND.n1798 GND.n1797 9.3
R4335 GND.n1793 GND.n1792 9.3
R4336 GND.n1788 GND.n1787 9.3
R4337 GND.n1783 GND.n1782 9.3
R4338 GND.n1778 GND.n1777 9.3
R4339 GND.n1771 GND.n1770 9.3
R4340 GND.n1758 GND.n1757 9.3
R4341 GND.n1753 GND.n1752 9.3
R4342 GND.n1748 GND.n1747 9.3
R4343 GND.n1745 GND.n1744 9.3
R4344 GND.n1741 GND.n1740 9.3
R4345 GND.n1738 GND.n1737 9.3
R4346 GND.n1734 GND.n1733 9.3
R4347 GND.n1731 GND.n1730 9.3
R4348 GND.n1727 GND.n1726 9.3
R4349 GND.n1724 GND.n1723 9.3
R4350 GND.n1720 GND.n1719 9.3
R4351 GND.n1717 GND.n1716 9.3
R4352 GND.n1713 GND.n1712 9.3
R4353 GND.n1710 GND.n1709 9.3
R4354 GND.n1706 GND.n1705 9.3
R4355 GND.n1703 GND.n1702 9.3
R4356 GND.n1699 GND.n1698 9.3
R4357 GND.n1814 GND.n1813 9.3
R4358 GND.n1656 GND.n1655 9.3
R4359 GND.n1636 GND.n1635 9.3
R4360 GND.n9490 GND.n9489 9.3
R4361 GND.n9472 GND.n9471 9.3
R4362 GND.n9465 GND.n9464 9.3
R4363 GND.n9458 GND.n9457 9.3
R4364 GND.n9451 GND.n9450 9.3
R4365 GND.n9444 GND.n9443 9.3
R4366 GND.n9437 GND.n9436 9.3
R4367 GND.n9430 GND.n9429 9.3
R4368 GND.n9425 GND.n9424 9.3
R4369 GND.n9428 GND.n9427 9.3
R4370 GND.n9432 GND.n9431 9.3
R4371 GND.n9435 GND.n9434 9.3
R4372 GND.n9439 GND.n9438 9.3
R4373 GND.n9442 GND.n9441 9.3
R4374 GND.n9446 GND.n9445 9.3
R4375 GND.n9449 GND.n9448 9.3
R4376 GND.n9453 GND.n9452 9.3
R4377 GND.n9456 GND.n9455 9.3
R4378 GND.n9460 GND.n9459 9.3
R4379 GND.n9463 GND.n9462 9.3
R4380 GND.n9468 GND.n9467 9.3
R4381 GND.n9470 GND.n9469 9.3
R4382 GND.n9475 GND.n9474 9.3
R4383 GND.n9481 GND.n9480 9.3
R4384 GND.n9488 GND.n9487 9.3
R4385 GND.n9494 GND.n9493 9.3
R4386 GND.n1648 GND.n1647 9.3
R4387 GND.n1652 GND.n1651 9.3
R4388 GND.n1658 GND.n1657 9.3
R4389 GND.n1662 GND.n1661 9.3
R4390 GND.n1667 GND.n1666 9.3
R4391 GND.n1672 GND.n1671 9.3
R4392 GND.n1676 GND.n1675 9.3
R4393 GND.n1680 GND.n1679 9.3
R4394 GND.n9421 GND.n9420 9.3
R4395 GND.n9423 GND.n9422 9.3
R4396 GND.n1622 GND.n1621 9.3
R4397 GND.n1633 GND.n1632 9.3
R4398 GND.n1823 GND.n1822 9.3
R4399 GND.n1845 GND.n1844 9.3
R4400 GND.n1852 GND.n1851 9.3
R4401 GND.n1859 GND.n1858 9.3
R4402 GND.n1866 GND.n1865 9.3
R4403 GND.n1873 GND.n1872 9.3
R4404 GND.n1880 GND.n1879 9.3
R4405 GND.n1887 GND.n1886 9.3
R4406 GND.n1892 GND.n1891 9.3
R4407 GND.n1890 GND.n1889 9.3
R4408 GND.n1885 GND.n1884 9.3
R4409 GND.n1883 GND.n1882 9.3
R4410 GND.n1878 GND.n1877 9.3
R4411 GND.n1876 GND.n1875 9.3
R4412 GND.n1871 GND.n1870 9.3
R4413 GND.n1869 GND.n1868 9.3
R4414 GND.n1864 GND.n1863 9.3
R4415 GND.n1862 GND.n1861 9.3
R4416 GND.n1857 GND.n1856 9.3
R4417 GND.n1855 GND.n1854 9.3
R4418 GND.n1850 GND.n1849 9.3
R4419 GND.n1847 GND.n1846 9.3
R4420 GND.n1843 GND.n1842 9.3
R4421 GND.n1836 GND.n1835 9.3
R4422 GND.n1825 GND.n1824 9.3
R4423 GND.n1819 GND.n1818 9.3
R4424 GND.n1631 GND.n1630 9.3
R4425 GND.n1627 GND.n1626 9.3
R4426 GND.n1620 GND.n1619 9.3
R4427 GND.n1616 GND.n1615 9.3
R4428 GND.n1610 GND.n1609 9.3
R4429 GND.n1594 GND.n1593 9.3
R4430 GND.n1589 GND.n1588 9.3
R4431 GND.n1584 GND.n1583 9.3
R4432 GND.n1896 GND.n1895 9.3
R4433 GND.n1894 GND.n1893 9.3
R4434 GND.n8694 GND.n8693 9.3
R4435 GND.n8687 GND.n8686 9.3
R4436 GND.n8680 GND.n8679 9.3
R4437 GND.n8673 GND.n8672 9.3
R4438 GND.n8666 GND.n8665 9.3
R4439 GND.n8659 GND.n8658 9.3
R4440 GND.n8652 GND.n8651 9.3
R4441 GND.n8645 GND.n8644 9.3
R4442 GND.n8630 GND.n8629 9.3
R4443 GND.n8622 GND.n8621 9.3
R4444 GND.n8612 GND.n8611 9.3
R4445 GND.n8594 GND.n8593 9.3
R4446 GND.n8598 GND.n8597 9.3
R4447 GND.n8602 GND.n8601 9.3
R4448 GND.n8606 GND.n8605 9.3
R4449 GND.n8610 GND.n8609 9.3
R4450 GND.n8616 GND.n8615 9.3
R4451 GND.n8620 GND.n8619 9.3
R4452 GND.n8626 GND.n8625 9.3
R4453 GND.n8632 GND.n8631 9.3
R4454 GND.n8638 GND.n8637 9.3
R4455 GND.n8643 GND.n8642 9.3
R4456 GND.n8648 GND.n8647 9.3
R4457 GND.n8650 GND.n8649 9.3
R4458 GND.n8655 GND.n8654 9.3
R4459 GND.n8657 GND.n8656 9.3
R4460 GND.n8662 GND.n8661 9.3
R4461 GND.n8664 GND.n8663 9.3
R4462 GND.n8669 GND.n8668 9.3
R4463 GND.n8671 GND.n8670 9.3
R4464 GND.n8676 GND.n8675 9.3
R4465 GND.n8678 GND.n8677 9.3
R4466 GND.n8683 GND.n8682 9.3
R4467 GND.n8685 GND.n8684 9.3
R4468 GND.n8690 GND.n8689 9.3
R4469 GND.n8692 GND.n8691 9.3
R4470 GND.n8696 GND.n8695 9.3
R4471 GND.n8590 GND.n8589 9.3
R4472 GND.n1570 GND.n1569 9.3
R4473 GND.n1578 GND.n1577 9.3
R4474 GND.n1577 GND.n1576 9.3
R4475 GND.n1580 GND.n1579 9.3
R4476 GND.n1694 GND.n1693 9.3
R4477 GND.n1693 GND.n1692 9.3
R4478 GND.n1683 GND.n1682 9.3
R4479 GND.n1686 GND.n1685 9.3
R4480 GND.n10129 GND.n10128 9.3
R4481 GND.n10128 GND.n10127 9.3
R4482 GND.n10119 GND.n10118 9.3
R4483 GND.n10107 GND.n10106 9.3
R4484 GND.n10095 GND.n10094 9.3
R4485 GND.n10083 GND.n10082 9.3
R4486 GND.n10071 GND.n10070 9.3
R4487 GND.n10059 GND.n10058 9.3
R4488 GND.n10041 GND.n10040 9.3
R4489 GND.n10029 GND.n10028 9.3
R4490 GND.n10017 GND.n10016 9.3
R4491 GND.n10005 GND.n10004 9.3
R4492 GND.n9993 GND.n9992 9.3
R4493 GND.n9980 GND.n9979 9.3
R4494 GND.n9978 GND.n9977 9.3
R4495 GND.n9989 GND.n9988 9.3
R4496 GND.n9988 GND.n9987 9.3
R4497 GND.n9991 GND.n9990 9.3
R4498 GND.n10001 GND.n10000 9.3
R4499 GND.n10000 GND.n9999 9.3
R4500 GND.n10003 GND.n10002 9.3
R4501 GND.n10013 GND.n10012 9.3
R4502 GND.n10012 GND.n10011 9.3
R4503 GND.n10015 GND.n10014 9.3
R4504 GND.n10025 GND.n10024 9.3
R4505 GND.n10024 GND.n10023 9.3
R4506 GND.n10027 GND.n10026 9.3
R4507 GND.n10037 GND.n10036 9.3
R4508 GND.n10036 GND.n10035 9.3
R4509 GND.n10039 GND.n10038 9.3
R4510 GND.n10049 GND.n10048 9.3
R4511 GND.n10048 GND.n10047 9.3
R4512 GND.n10057 GND.n10056 9.3
R4513 GND.n10056 GND.n10055 9.3
R4514 GND.n10061 GND.n10060 9.3
R4515 GND.n10069 GND.n10068 9.3
R4516 GND.n10068 GND.n10067 9.3
R4517 GND.n10073 GND.n10072 9.3
R4518 GND.n10081 GND.n10080 9.3
R4519 GND.n10080 GND.n10079 9.3
R4520 GND.n10085 GND.n10084 9.3
R4521 GND.n10093 GND.n10092 9.3
R4522 GND.n10092 GND.n10091 9.3
R4523 GND.n10097 GND.n10096 9.3
R4524 GND.n10105 GND.n10104 9.3
R4525 GND.n10104 GND.n10103 9.3
R4526 GND.n10109 GND.n10108 9.3
R4527 GND.n10117 GND.n10116 9.3
R4528 GND.n10116 GND.n10115 9.3
R4529 GND.n10121 GND.n10120 9.3
R4530 GND.n9976 GND.n9975 9.3
R4531 GND.n9975 GND.n9974 9.3
R4532 GND.n9965 GND.n9964 9.3
R4533 GND.n9967 GND.n9966 9.3
R4534 GND.n10131 GND.n10130 9.3
R4535 GND.n10133 GND.n10132 9.3
R4536 GND.n9291 GND.n9290 9.3
R4537 GND.n9264 GND.n9263 9.3
R4538 GND.n9259 GND.n9258 9.3
R4539 GND.n9272 GND.n9271 9.3
R4540 GND.n9271 GND.n9270 9.3
R4541 GND.n9289 GND.n9288 9.3
R4542 GND.n9288 GND.n9287 9.3
R4543 GND.n9419 GND.n9418 9.3
R4544 GND.n9257 GND.n9256 9.3
R4545 GND.n9251 GND.n9250 9.3
R4546 GND.n8938 GND.n8937 9.3
R4547 GND.n8937 GND.n8936 9.3
R4548 GND.n8936 GND.n8935 9.3
R4549 GND.n8942 GND.n8941 9.3
R4550 GND.n8954 GND.n8953 9.3
R4551 GND.n8967 GND.n8966 9.3
R4552 GND.n8979 GND.n8978 9.3
R4553 GND.n8992 GND.n8991 9.3
R4554 GND.n9014 GND.n9013 9.3
R4555 GND.n9022 GND.n9021 9.3
R4556 GND.n9030 GND.n9029 9.3
R4557 GND.n9038 GND.n9037 9.3
R4558 GND.n9046 GND.n9045 9.3
R4559 GND.n9054 GND.n9053 9.3
R4560 GND.n9062 GND.n9061 9.3
R4561 GND.n9068 GND.n9067 9.3
R4562 GND.n9073 GND.n9072 9.3
R4563 GND.n9078 GND.n9077 9.3
R4564 GND.n9097 GND.n9096 9.3
R4565 GND.n9115 GND.n9114 9.3
R4566 GND.n9127 GND.n9126 9.3
R4567 GND.n9139 GND.n9138 9.3
R4568 GND.n9151 GND.n9150 9.3
R4569 GND.n9163 GND.n9162 9.3
R4570 GND.n9176 GND.n9175 9.3
R4571 GND.n9178 GND.n9177 9.3
R4572 GND.n9165 GND.n9164 9.3
R4573 GND.n9153 GND.n9152 9.3
R4574 GND.n9141 GND.n9140 9.3
R4575 GND.n9129 GND.n9128 9.3
R4576 GND.n9117 GND.n9116 9.3
R4577 GND.n9095 GND.n9094 9.3
R4578 GND.n9085 GND.n9084 9.3
R4579 GND.n9081 GND.n9080 9.3
R4580 GND.n9076 GND.n9075 9.3
R4581 GND.n9071 GND.n9070 9.3
R4582 GND.n9066 GND.n9065 9.3
R4583 GND.n9064 GND.n9063 9.3
R4584 GND.n9060 GND.n9059 9.3
R4585 GND.n8935 GND.n8934 9.3
R4586 GND.n9056 GND.n9055 9.3
R4587 GND.n9052 GND.n9051 9.3
R4588 GND.n9048 GND.n9047 9.3
R4589 GND.n9044 GND.n9043 9.3
R4590 GND.n9040 GND.n9039 9.3
R4591 GND.n9036 GND.n9035 9.3
R4592 GND.n9032 GND.n9031 9.3
R4593 GND.n9028 GND.n9027 9.3
R4594 GND.n9024 GND.n9023 9.3
R4595 GND.n9020 GND.n9019 9.3
R4596 GND.n9016 GND.n9015 9.3
R4597 GND.n9012 GND.n9011 9.3
R4598 GND.n9005 GND.n9004 9.3
R4599 GND.n9004 GND.n9003 9.3
R4600 GND.n8990 GND.n8989 9.3
R4601 GND.n8988 GND.n8987 9.3
R4602 GND.n8987 GND.n8986 9.3
R4603 GND.n8977 GND.n8976 9.3
R4604 GND.n8975 GND.n8974 9.3
R4605 GND.n8974 GND.n8973 9.3
R4606 GND.n8965 GND.n8964 9.3
R4607 GND.n8963 GND.n8962 9.3
R4608 GND.n8962 GND.n8961 9.3
R4609 GND.n8952 GND.n8951 9.3
R4610 GND.n8950 GND.n8949 9.3
R4611 GND.n8949 GND.n8948 9.3
R4612 GND.n8940 GND.n8939 9.3
R4613 GND.n9231 GND.n9230 9.3
R4614 GND.n9229 GND.n9228 9.3
R4615 GND.n8893 GND.n8892 9.3
R4616 GND.n8891 GND.n8890 9.3
R4617 GND.n9174 GND.n9173 9.3
R4618 GND.n9173 GND.n9172 9.3
R4619 GND.n9161 GND.n9160 9.3
R4620 GND.n9160 GND.n9159 9.3
R4621 GND.n9149 GND.n9148 9.3
R4622 GND.n9148 GND.n9147 9.3
R4623 GND.n9137 GND.n9136 9.3
R4624 GND.n9136 GND.n9135 9.3
R4625 GND.n9125 GND.n9124 9.3
R4626 GND.n9124 GND.n9123 9.3
R4627 GND.n9113 GND.n9112 9.3
R4628 GND.n9112 GND.n9111 9.3
R4629 GND.n9105 GND.n9104 9.3
R4630 GND.n9104 GND.n9103 9.3
R4631 GND.n9091 GND.n9090 9.3
R4632 GND.n9200 GND.n9199 9.3
R4633 GND.n9212 GND.n9211 9.3
R4634 GND.n9193 GND.n9192 9.3
R4635 GND.n9219 GND.n9218 9.3
R4636 GND.n9186 GND.n9185 9.3
R4637 GND.n9227 GND.n9226 9.3
R4638 GND.n9226 GND.n9225 9.3
R4639 GND.n4487 GND.n4486 9.3
R4640 GND.n4475 GND.n4474 9.3
R4641 GND.n4462 GND.n4461 9.3
R4642 GND.n4450 GND.n4449 9.3
R4643 GND.n4437 GND.n4436 9.3
R4644 GND.n4415 GND.n4414 9.3
R4645 GND.n4407 GND.n4406 9.3
R4646 GND.n4399 GND.n4398 9.3
R4647 GND.n4391 GND.n4390 9.3
R4648 GND.n4383 GND.n4382 9.3
R4649 GND.n4375 GND.n4374 9.3
R4650 GND.n4367 GND.n4366 9.3
R4651 GND.n4361 GND.n4360 9.3
R4652 GND.n4356 GND.n4355 9.3
R4653 GND.n4351 GND.n4350 9.3
R4654 GND.n4332 GND.n4331 9.3
R4655 GND.n4313 GND.n4312 9.3
R4656 GND.n4300 GND.n4299 9.3
R4657 GND.n4288 GND.n4287 9.3
R4658 GND.n4275 GND.n4274 9.3
R4659 GND.n4263 GND.n4262 9.3
R4660 GND.n4250 GND.n4249 9.3
R4661 GND.n4248 GND.n4247 9.3
R4662 GND.n4261 GND.n4260 9.3
R4663 GND.n4273 GND.n4272 9.3
R4664 GND.n4286 GND.n4285 9.3
R4665 GND.n4298 GND.n4297 9.3
R4666 GND.n4311 GND.n4310 9.3
R4667 GND.n4334 GND.n4333 9.3
R4668 GND.n4344 GND.n4343 9.3
R4669 GND.n4348 GND.n4347 9.3
R4670 GND.n4353 GND.n4352 9.3
R4671 GND.n4358 GND.n4357 9.3
R4672 GND.n4363 GND.n4362 9.3
R4673 GND.n4365 GND.n4364 9.3
R4674 GND.n4373 GND.n4372 9.3
R4675 GND.n4381 GND.n4380 9.3
R4676 GND.n4389 GND.n4388 9.3
R4677 GND.n4397 GND.n4396 9.3
R4678 GND.n4405 GND.n4404 9.3
R4679 GND.n4413 GND.n4412 9.3
R4680 GND.n4439 GND.n4438 9.3
R4681 GND.n4452 GND.n4451 9.3
R4682 GND.n4464 GND.n4463 9.3
R4683 GND.n4477 GND.n4476 9.3
R4684 GND.n4489 GND.n4488 9.3
R4685 GND.n1915 GND.n1914 9.3
R4686 GND.n4194 GND.n4193 9.3
R4687 GND.n4536 GND.n4535 9.3
R4688 GND.n4538 GND.n4537 9.3
R4689 GND.n4534 GND.n4533 9.3
R4690 GND.n4533 GND.n4532 9.3
R4691 GND.n4532 GND.n4531 9.3
R4692 GND.n4259 GND.n4258 9.3
R4693 GND.n4258 GND.n4257 9.3
R4694 GND.n4271 GND.n4270 9.3
R4695 GND.n4270 GND.n4269 9.3
R4696 GND.n4284 GND.n4283 9.3
R4697 GND.n4283 GND.n4282 9.3
R4698 GND.n4296 GND.n4295 9.3
R4699 GND.n4295 GND.n4294 9.3
R4700 GND.n4309 GND.n4308 9.3
R4701 GND.n4308 GND.n4307 9.3
R4702 GND.n4322 GND.n4321 9.3
R4703 GND.n4321 GND.n4320 9.3
R4704 GND.n4330 GND.n4329 9.3
R4705 GND.n4329 GND.n4328 9.3
R4706 GND.n4338 GND.n4337 9.3
R4707 GND.n4233 GND.n4232 9.3
R4708 GND.n4228 GND.n4227 9.3
R4709 GND.n4217 GND.n4216 9.3
R4710 GND.n4212 GND.n4211 9.3
R4711 GND.n4202 GND.n4201 9.3
R4712 GND.n4371 GND.n4370 9.3
R4713 GND.n4531 GND.n4530 9.3
R4714 GND.n4379 GND.n4378 9.3
R4715 GND.n4387 GND.n4386 9.3
R4716 GND.n4395 GND.n4394 9.3
R4717 GND.n4403 GND.n4402 9.3
R4718 GND.n4411 GND.n4410 9.3
R4719 GND.n4419 GND.n4418 9.3
R4720 GND.n4435 GND.n4434 9.3
R4721 GND.n4434 GND.n4433 9.3
R4722 GND.n4448 GND.n4447 9.3
R4723 GND.n4447 GND.n4446 9.3
R4724 GND.n4460 GND.n4459 9.3
R4725 GND.n4459 GND.n4458 9.3
R4726 GND.n4473 GND.n4472 9.3
R4727 GND.n4472 GND.n4471 9.3
R4728 GND.n4485 GND.n4484 9.3
R4729 GND.n4484 GND.n4483 9.3
R4730 GND.n4246 GND.n4245 9.3
R4731 GND.n4245 GND.n4244 9.3
R4732 GND.n2496 GND.n2495 9.3
R4733 GND.n2501 GND.n2500 9.3
R4734 GND.n2508 GND.n2507 9.3
R4735 GND.n2515 GND.n2514 9.3
R4736 GND.n2522 GND.n2521 9.3
R4737 GND.n2529 GND.n2528 9.3
R4738 GND.n2536 GND.n2535 9.3
R4739 GND.n2543 GND.n2542 9.3
R4740 GND.n2565 GND.n2564 9.3
R4741 GND.n2573 GND.n2572 9.3
R4742 GND.n2499 GND.n2498 9.3
R4743 GND.n2503 GND.n2502 9.3
R4744 GND.n2506 GND.n2505 9.3
R4745 GND.n2510 GND.n2509 9.3
R4746 GND.n2513 GND.n2512 9.3
R4747 GND.n2517 GND.n2516 9.3
R4748 GND.n2520 GND.n2519 9.3
R4749 GND.n2524 GND.n2523 9.3
R4750 GND.n2527 GND.n2526 9.3
R4751 GND.n2531 GND.n2530 9.3
R4752 GND.n2534 GND.n2533 9.3
R4753 GND.n2538 GND.n2537 9.3
R4754 GND.n2541 GND.n2540 9.3
R4755 GND.n2546 GND.n2545 9.3
R4756 GND.n2551 GND.n2550 9.3
R4757 GND.n2563 GND.n2562 9.3
R4758 GND.n2570 GND.n2569 9.3
R4759 GND.n2575 GND.n2574 9.3
R4760 GND.n2580 GND.n2579 9.3
R4761 GND.n2494 GND.n2493 9.3
R4762 GND.n2492 GND.n2491 9.3
R4763 GND.n2593 GND.n2592 9.3
R4764 GND.n2599 GND.n2598 9.3
R4765 GND.n2602 GND.n2601 9.3
R4766 GND.n2607 GND.n2606 9.3
R4767 GND.n2590 GND.n2589 9.3
R4768 GND.n2585 GND.n2584 9.3
R4769 GND.n2583 GND.n2582 9.3
R4770 GND.n2255 GND.n2254 9.3
R4771 GND.n2266 GND.n2265 9.3
R4772 GND.n3471 GND.n3470 9.3
R4773 GND.n3453 GND.n3452 9.3
R4774 GND.n3446 GND.n3445 9.3
R4775 GND.n3439 GND.n3438 9.3
R4776 GND.n3432 GND.n3431 9.3
R4777 GND.n3425 GND.n3424 9.3
R4778 GND.n3418 GND.n3417 9.3
R4779 GND.n3411 GND.n3410 9.3
R4780 GND.n3406 GND.n3405 9.3
R4781 GND.n3409 GND.n3408 9.3
R4782 GND.n3413 GND.n3412 9.3
R4783 GND.n3416 GND.n3415 9.3
R4784 GND.n3420 GND.n3419 9.3
R4785 GND.n3423 GND.n3422 9.3
R4786 GND.n3427 GND.n3426 9.3
R4787 GND.n3430 GND.n3429 9.3
R4788 GND.n3434 GND.n3433 9.3
R4789 GND.n3437 GND.n3436 9.3
R4790 GND.n3441 GND.n3440 9.3
R4791 GND.n3444 GND.n3443 9.3
R4792 GND.n3449 GND.n3448 9.3
R4793 GND.n3451 GND.n3450 9.3
R4794 GND.n3456 GND.n3455 9.3
R4795 GND.n3462 GND.n3461 9.3
R4796 GND.n3469 GND.n3468 9.3
R4797 GND.n3475 GND.n3474 9.3
R4798 GND.n2264 GND.n2263 9.3
R4799 GND.n2260 GND.n2259 9.3
R4800 GND.n2253 GND.n2252 9.3
R4801 GND.n2249 GND.n2248 9.3
R4802 GND.n2243 GND.n2242 9.3
R4803 GND.n2465 GND.n2464 9.3
R4804 GND.n2469 GND.n2468 9.3
R4805 GND.n2473 GND.n2472 9.3
R4806 GND.n3402 GND.n3401 9.3
R4807 GND.n3404 GND.n3403 9.3
R4808 GND.n2226 GND.n2225 9.3
R4809 GND.n2237 GND.n2236 9.3
R4810 GND.n2402 GND.n2401 9.3
R4811 GND.n2449 GND.n2448 9.3
R4812 GND.n2442 GND.n2441 9.3
R4813 GND.n2435 GND.n2434 9.3
R4814 GND.n2428 GND.n2427 9.3
R4815 GND.n2421 GND.n2420 9.3
R4816 GND.n2615 GND.n2614 9.3
R4817 GND.n2622 GND.n2621 9.3
R4818 GND.n2627 GND.n2626 9.3
R4819 GND.n2625 GND.n2624 9.3
R4820 GND.n2620 GND.n2619 9.3
R4821 GND.n2618 GND.n2617 9.3
R4822 GND.n2613 GND.n2612 9.3
R4823 GND.n2611 GND.n2610 9.3
R4824 GND.n2423 GND.n2422 9.3
R4825 GND.n2426 GND.n2425 9.3
R4826 GND.n2430 GND.n2429 9.3
R4827 GND.n2433 GND.n2432 9.3
R4828 GND.n2437 GND.n2436 9.3
R4829 GND.n2440 GND.n2439 9.3
R4830 GND.n2444 GND.n2443 9.3
R4831 GND.n2447 GND.n2446 9.3
R4832 GND.n2452 GND.n2451 9.3
R4833 GND.n2419 GND.n2418 9.3
R4834 GND.n2404 GND.n2403 9.3
R4835 GND.n2397 GND.n2396 9.3
R4836 GND.n2235 GND.n2234 9.3
R4837 GND.n2231 GND.n2230 9.3
R4838 GND.n2224 GND.n2223 9.3
R4839 GND.n2220 GND.n2219 9.3
R4840 GND.n2214 GND.n2213 9.3
R4841 GND.n2209 GND.n2208 9.3
R4842 GND.n2203 GND.n2202 9.3
R4843 GND.n3163 GND.n3162 9.3
R4844 GND.n2631 GND.n2630 9.3
R4845 GND.n2629 GND.n2628 9.3
R4846 GND.n2305 GND.n2304 9.3
R4847 GND.n3151 GND.n3150 9.3
R4848 GND.n2339 GND.n2338 9.3
R4849 GND.n2346 GND.n2345 9.3
R4850 GND.n2353 GND.n2352 9.3
R4851 GND.n2360 GND.n2359 9.3
R4852 GND.n2367 GND.n2366 9.3
R4853 GND.n2374 GND.n2373 9.3
R4854 GND.n2381 GND.n2380 9.3
R4855 GND.n2278 GND.n2277 9.3
R4856 GND.n2280 GND.n2279 9.3
R4857 GND.n2337 GND.n2336 9.3
R4858 GND.n2341 GND.n2340 9.3
R4859 GND.n2344 GND.n2343 9.3
R4860 GND.n2348 GND.n2347 9.3
R4861 GND.n2351 GND.n2350 9.3
R4862 GND.n2355 GND.n2354 9.3
R4863 GND.n2358 GND.n2357 9.3
R4864 GND.n2362 GND.n2361 9.3
R4865 GND.n2365 GND.n2364 9.3
R4866 GND.n2369 GND.n2368 9.3
R4867 GND.n2372 GND.n2371 9.3
R4868 GND.n2376 GND.n2375 9.3
R4869 GND.n2379 GND.n2378 9.3
R4870 GND.n2384 GND.n2383 9.3
R4871 GND.n2333 GND.n2332 9.3
R4872 GND.n2284 GND.n2283 9.3
R4873 GND.n2289 GND.n2288 9.3
R4874 GND.n2287 GND.n2286 9.3
R4875 GND.n2318 GND.n2317 9.3
R4876 GND.n2309 GND.n2308 9.3
R4877 GND.n2313 GND.n2312 9.3
R4878 GND.n2328 GND.n2327 9.3
R4879 GND.n2323 GND.n2322 9.3
R4880 GND.n2321 GND.n2320 9.3
R4881 GND.n3153 GND.n3152 9.3
R4882 GND.n3155 GND.n3154 9.3
R4883 GND.n2301 GND.n2300 9.3
R4884 GND.n2479 GND.n2478 9.3
R4885 GND.n3174 GND.n3173 9.3
R4886 GND.n3177 GND.n3176 9.3
R4887 GND.n3172 GND.n3171 9.3
R4888 GND.n3171 GND.n3170 9.3
R4889 GND.n2487 GND.n2486 9.3
R4890 GND.n2486 GND.n2485 9.3
R4891 GND.n2476 GND.n2475 9.3
R4892 GND.n1919 GND.n1918 9.3
R4893 GND.n4938 GND.n4937 9.3
R4894 GND.n4951 GND.n4950 9.3
R4895 GND.n4963 GND.n4962 9.3
R4896 GND.n4976 GND.n4975 9.3
R4897 GND.n4988 GND.n4987 9.3
R4898 GND.n5001 GND.n5000 9.3
R4899 GND.n5020 GND.n5019 9.3
R4900 GND.n5033 GND.n5032 9.3
R4901 GND.n5045 GND.n5044 9.3
R4902 GND.n5058 GND.n5057 9.3
R4903 GND.n5070 GND.n5069 9.3
R4904 GND.n5083 GND.n5082 9.3
R4905 GND.n5097 GND.n5096 9.3
R4906 GND.n4936 GND.n4935 9.3
R4907 GND.n4947 GND.n4946 9.3
R4908 GND.n4946 GND.n4945 9.3
R4909 GND.n4949 GND.n4948 9.3
R4910 GND.n4959 GND.n4958 9.3
R4911 GND.n4958 GND.n4957 9.3
R4912 GND.n4961 GND.n4960 9.3
R4913 GND.n4972 GND.n4971 9.3
R4914 GND.n4971 GND.n4970 9.3
R4915 GND.n4974 GND.n4973 9.3
R4916 GND.n4984 GND.n4983 9.3
R4917 GND.n4983 GND.n4982 9.3
R4918 GND.n4986 GND.n4985 9.3
R4919 GND.n4997 GND.n4996 9.3
R4920 GND.n4996 GND.n4995 9.3
R4921 GND.n4999 GND.n4998 9.3
R4922 GND.n5010 GND.n5009 9.3
R4923 GND.n5009 GND.n5008 9.3
R4924 GND.n5018 GND.n5017 9.3
R4925 GND.n5017 GND.n5016 9.3
R4926 GND.n5022 GND.n5021 9.3
R4927 GND.n5031 GND.n5030 9.3
R4928 GND.n5030 GND.n5029 9.3
R4929 GND.n5035 GND.n5034 9.3
R4930 GND.n5043 GND.n5042 9.3
R4931 GND.n5042 GND.n5041 9.3
R4932 GND.n5047 GND.n5046 9.3
R4933 GND.n5056 GND.n5055 9.3
R4934 GND.n5055 GND.n5054 9.3
R4935 GND.n5060 GND.n5059 9.3
R4936 GND.n5068 GND.n5067 9.3
R4937 GND.n5067 GND.n5066 9.3
R4938 GND.n5072 GND.n5071 9.3
R4939 GND.n5081 GND.n5080 9.3
R4940 GND.n5080 GND.n5079 9.3
R4941 GND.n5085 GND.n5084 9.3
R4942 GND.n5093 GND.n5092 9.3
R4943 GND.n5092 GND.n5091 9.3
R4944 GND.n5095 GND.n5094 9.3
R4945 GND.n4925 GND.n4924 9.3
R4946 GND.n4934 GND.n4933 9.3
R4947 GND.n4933 GND.n4932 9.3
R4948 GND.n3395 GND.n3394 9.3
R4949 GND.n3368 GND.n3367 9.3
R4950 GND.n3366 GND.n3365 9.3
R4951 GND.n3376 GND.n3375 9.3
R4952 GND.n3375 GND.n3374 9.3
R4953 GND.n3393 GND.n3392 9.3
R4954 GND.n3392 GND.n3391 9.3
R4955 GND.n3400 GND.n3399 9.3
R4956 GND.n5201 GND.n5200 9.3
R4957 GND.n5105 GND.n5104 9.3
R4958 GND.n5110 GND.n5109 9.3
R4959 GND.n5117 GND.n5116 9.3
R4960 GND.n5124 GND.n5123 9.3
R4961 GND.n5131 GND.n5130 9.3
R4962 GND.n5138 GND.n5137 9.3
R4963 GND.n5145 GND.n5144 9.3
R4964 GND.n5152 GND.n5151 9.3
R4965 GND.n5173 GND.n5172 9.3
R4966 GND.n5181 GND.n5180 9.3
R4967 GND.n5108 GND.n5107 9.3
R4968 GND.n5112 GND.n5111 9.3
R4969 GND.n5115 GND.n5114 9.3
R4970 GND.n5119 GND.n5118 9.3
R4971 GND.n5122 GND.n5121 9.3
R4972 GND.n5126 GND.n5125 9.3
R4973 GND.n5129 GND.n5128 9.3
R4974 GND.n5133 GND.n5132 9.3
R4975 GND.n5136 GND.n5135 9.3
R4976 GND.n5140 GND.n5139 9.3
R4977 GND.n5143 GND.n5142 9.3
R4978 GND.n5147 GND.n5146 9.3
R4979 GND.n5150 GND.n5149 9.3
R4980 GND.n5155 GND.n5154 9.3
R4981 GND.n5160 GND.n5159 9.3
R4982 GND.n5171 GND.n5170 9.3
R4983 GND.n5178 GND.n5177 9.3
R4984 GND.n5183 GND.n5182 9.3
R4985 GND.n5188 GND.n5187 9.3
R4986 GND.n5198 GND.n5197 9.3
R4987 GND.n5193 GND.n5192 9.3
R4988 GND.n5191 GND.n5190 9.3
R4989 GND.n5103 GND.n5102 9.3
R4990 GND.n5101 GND.n5100 9.3
R4991 GND.n5210 GND.n5209 9.3
R4992 GND.n5215 GND.n5214 9.3
R4993 GND.n5207 GND.n5206 9.3
R4994 GND.n2042 GND.n2041 9.3
R4995 GND.n2053 GND.n2052 9.3
R4996 GND.n2128 GND.n2127 9.3
R4997 GND.n2110 GND.n2109 9.3
R4998 GND.n2103 GND.n2102 9.3
R4999 GND.n2096 GND.n2095 9.3
R5000 GND.n2089 GND.n2088 9.3
R5001 GND.n2082 GND.n2081 9.3
R5002 GND.n2075 GND.n2074 9.3
R5003 GND.n2068 GND.n2067 9.3
R5004 GND.n2063 GND.n2062 9.3
R5005 GND.n2066 GND.n2065 9.3
R5006 GND.n2070 GND.n2069 9.3
R5007 GND.n2073 GND.n2072 9.3
R5008 GND.n2077 GND.n2076 9.3
R5009 GND.n2080 GND.n2079 9.3
R5010 GND.n2084 GND.n2083 9.3
R5011 GND.n2087 GND.n2086 9.3
R5012 GND.n2091 GND.n2090 9.3
R5013 GND.n2094 GND.n2093 9.3
R5014 GND.n2098 GND.n2097 9.3
R5015 GND.n2101 GND.n2100 9.3
R5016 GND.n2106 GND.n2105 9.3
R5017 GND.n2108 GND.n2107 9.3
R5018 GND.n2113 GND.n2112 9.3
R5019 GND.n2119 GND.n2118 9.3
R5020 GND.n2126 GND.n2125 9.3
R5021 GND.n2132 GND.n2131 9.3
R5022 GND.n2051 GND.n2050 9.3
R5023 GND.n2047 GND.n2046 9.3
R5024 GND.n2040 GND.n2039 9.3
R5025 GND.n2036 GND.n2035 9.3
R5026 GND.n2030 GND.n2029 9.3
R5027 GND.n2015 GND.n2014 9.3
R5028 GND.n2010 GND.n2009 9.3
R5029 GND.n2005 GND.n2004 9.3
R5030 GND.n1941 GND.n1940 9.3
R5031 GND.n2061 GND.n2060 9.3
R5032 GND.n1989 GND.n1988 9.3
R5033 GND.n2000 GND.n1999 9.3
R5034 GND.n2144 GND.n2143 9.3
R5035 GND.n2190 GND.n2189 9.3
R5036 GND.n2183 GND.n2182 9.3
R5037 GND.n2176 GND.n2175 9.3
R5038 GND.n2169 GND.n2168 9.3
R5039 GND.n2162 GND.n2161 9.3
R5040 GND.n2642 GND.n2641 9.3
R5041 GND.n2649 GND.n2648 9.3
R5042 GND.n2654 GND.n2653 9.3
R5043 GND.n2652 GND.n2651 9.3
R5044 GND.n2647 GND.n2646 9.3
R5045 GND.n2645 GND.n2644 9.3
R5046 GND.n2640 GND.n2639 9.3
R5047 GND.n2638 GND.n2637 9.3
R5048 GND.n2164 GND.n2163 9.3
R5049 GND.n2167 GND.n2166 9.3
R5050 GND.n2171 GND.n2170 9.3
R5051 GND.n2174 GND.n2173 9.3
R5052 GND.n2178 GND.n2177 9.3
R5053 GND.n2181 GND.n2180 9.3
R5054 GND.n2185 GND.n2184 9.3
R5055 GND.n2188 GND.n2187 9.3
R5056 GND.n2193 GND.n2192 9.3
R5057 GND.n2160 GND.n2159 9.3
R5058 GND.n2146 GND.n2145 9.3
R5059 GND.n2139 GND.n2138 9.3
R5060 GND.n1998 GND.n1997 9.3
R5061 GND.n1994 GND.n1993 9.3
R5062 GND.n1987 GND.n1986 9.3
R5063 GND.n1983 GND.n1982 9.3
R5064 GND.n1977 GND.n1976 9.3
R5065 GND.n1972 GND.n1971 9.3
R5066 GND.n1967 GND.n1966 9.3
R5067 GND.n1962 GND.n1961 9.3
R5068 GND.n2658 GND.n2657 9.3
R5069 GND.n2656 GND.n2655 9.3
R5070 GND.n2892 GND.n2891 9.3
R5071 GND.n2884 GND.n2883 9.3
R5072 GND.n2874 GND.n2873 9.3
R5073 GND.n2856 GND.n2855 9.3
R5074 GND.n2894 GND.n2893 9.3
R5075 GND.n2888 GND.n2887 9.3
R5076 GND.n2860 GND.n2859 9.3
R5077 GND.n2864 GND.n2863 9.3
R5078 GND.n2868 GND.n2867 9.3
R5079 GND.n2872 GND.n2871 9.3
R5080 GND.n2878 GND.n2877 9.3
R5081 GND.n2882 GND.n2881 9.3
R5082 GND.n2959 GND.n2958 9.3
R5083 GND.n2954 GND.n2953 9.3
R5084 GND.n2947 GND.n2946 9.3
R5085 GND.n2940 GND.n2939 9.3
R5086 GND.n2933 GND.n2932 9.3
R5087 GND.n2926 GND.n2925 9.3
R5088 GND.n2919 GND.n2918 9.3
R5089 GND.n2957 GND.n2956 9.3
R5090 GND.n2952 GND.n2951 9.3
R5091 GND.n2950 GND.n2949 9.3
R5092 GND.n2945 GND.n2944 9.3
R5093 GND.n2943 GND.n2942 9.3
R5094 GND.n2938 GND.n2937 9.3
R5095 GND.n2936 GND.n2935 9.3
R5096 GND.n2931 GND.n2930 9.3
R5097 GND.n2929 GND.n2928 9.3
R5098 GND.n2924 GND.n2923 9.3
R5099 GND.n2922 GND.n2921 9.3
R5100 GND.n2917 GND.n2916 9.3
R5101 GND.n2915 GND.n2914 9.3
R5102 GND.n2910 GND.n2909 9.3
R5103 GND.n2912 GND.n2911 9.3
R5104 GND.n2961 GND.n2960 9.3
R5105 GND.n2963 GND.n2962 9.3
R5106 GND.n2852 GND.n2851 9.3
R5107 GND.n2905 GND.n2904 9.3
R5108 GND.n4773 GND.n4772 9.3
R5109 GND.n1954 GND.n1953 9.3
R5110 GND.n1959 GND.n1958 9.3
R5111 GND.n1952 GND.n1951 9.3
R5112 GND.n1951 GND.n1950 9.3
R5113 GND.n4781 GND.n4780 9.3
R5114 GND.n4780 GND.n4779 9.3
R5115 GND.n4771 GND.n4770 9.3
R5116 GND.n4588 GND.n4587 9.3
R5117 GND.n4587 GND.n4586 9.3
R5118 GND.n4592 GND.n4591 9.3
R5119 GND.n4605 GND.n4604 9.3
R5120 GND.n4617 GND.n4616 9.3
R5121 GND.n4630 GND.n4629 9.3
R5122 GND.n4642 GND.n4641 9.3
R5123 GND.n4655 GND.n4654 9.3
R5124 GND.n4674 GND.n4673 9.3
R5125 GND.n4687 GND.n4686 9.3
R5126 GND.n4699 GND.n4698 9.3
R5127 GND.n4712 GND.n4711 9.3
R5128 GND.n4724 GND.n4723 9.3
R5129 GND.n4737 GND.n4736 9.3
R5130 GND.n4751 GND.n4750 9.3
R5131 GND.n4590 GND.n4589 9.3
R5132 GND.n4601 GND.n4600 9.3
R5133 GND.n4600 GND.n4599 9.3
R5134 GND.n4603 GND.n4602 9.3
R5135 GND.n4613 GND.n4612 9.3
R5136 GND.n4612 GND.n4611 9.3
R5137 GND.n4615 GND.n4614 9.3
R5138 GND.n4626 GND.n4625 9.3
R5139 GND.n4625 GND.n4624 9.3
R5140 GND.n4628 GND.n4627 9.3
R5141 GND.n4638 GND.n4637 9.3
R5142 GND.n4637 GND.n4636 9.3
R5143 GND.n4640 GND.n4639 9.3
R5144 GND.n4651 GND.n4650 9.3
R5145 GND.n4650 GND.n4649 9.3
R5146 GND.n4653 GND.n4652 9.3
R5147 GND.n4664 GND.n4663 9.3
R5148 GND.n4663 GND.n4662 9.3
R5149 GND.n4672 GND.n4671 9.3
R5150 GND.n4671 GND.n4670 9.3
R5151 GND.n4676 GND.n4675 9.3
R5152 GND.n4685 GND.n4684 9.3
R5153 GND.n4684 GND.n4683 9.3
R5154 GND.n4689 GND.n4688 9.3
R5155 GND.n4697 GND.n4696 9.3
R5156 GND.n4696 GND.n4695 9.3
R5157 GND.n4701 GND.n4700 9.3
R5158 GND.n4710 GND.n4709 9.3
R5159 GND.n4709 GND.n4708 9.3
R5160 GND.n4714 GND.n4713 9.3
R5161 GND.n4722 GND.n4721 9.3
R5162 GND.n4721 GND.n4720 9.3
R5163 GND.n4726 GND.n4725 9.3
R5164 GND.n4735 GND.n4734 9.3
R5165 GND.n4734 GND.n4733 9.3
R5166 GND.n4739 GND.n4738 9.3
R5167 GND.n4747 GND.n4746 9.3
R5168 GND.n4746 GND.n4745 9.3
R5169 GND.n4749 GND.n4748 9.3
R5170 GND.n4579 GND.n4578 9.3
R5171 GND.n1934 GND.n1933 9.3
R5172 GND.n4917 GND.n4916 9.3
R5173 GND.n2668 GND.n2667 9.3
R5174 GND.n4920 GND.n4919 9.3
R5175 GND.n4915 GND.n4914 9.3
R5176 GND.n4914 GND.n4913 9.3
R5177 GND.n2666 GND.n2665 9.3
R5178 GND.n2665 GND.n2664 9.3
R5179 GND.n2671 GND.n2670 9.3
R5180 GND.n2983 GND.n2982 9.3
R5181 GND.n2995 GND.n2994 9.3
R5182 GND.n3007 GND.n3006 9.3
R5183 GND.n3019 GND.n3018 9.3
R5184 GND.n3031 GND.n3030 9.3
R5185 GND.n3043 GND.n3042 9.3
R5186 GND.n3055 GND.n3054 9.3
R5187 GND.n3073 GND.n3072 9.3
R5188 GND.n3085 GND.n3084 9.3
R5189 GND.n3097 GND.n3096 9.3
R5190 GND.n3109 GND.n3108 9.3
R5191 GND.n3121 GND.n3120 9.3
R5192 GND.n3134 GND.n3133 9.3
R5193 GND.n3146 GND.n3145 9.3
R5194 GND.n3184 GND.n3183 9.3
R5195 GND.n3195 GND.n3194 9.3
R5196 GND.n3207 GND.n3206 9.3
R5197 GND.n3219 GND.n3218 9.3
R5198 GND.n3231 GND.n3230 9.3
R5199 GND.n3243 GND.n3242 9.3
R5200 GND.n3255 GND.n3254 9.3
R5201 GND.n3273 GND.n3272 9.3
R5202 GND.n3285 GND.n3284 9.3
R5203 GND.n3297 GND.n3296 9.3
R5204 GND.n3309 GND.n3308 9.3
R5205 GND.n3321 GND.n3320 9.3
R5206 GND.n3334 GND.n3333 9.3
R5207 GND.n3347 GND.n3346 9.3
R5208 GND.n3136 GND.n3135 9.3
R5209 GND.n3132 GND.n3131 9.3
R5210 GND.n3131 GND.n3130 9.3
R5211 GND.n3123 GND.n3122 9.3
R5212 GND.n3119 GND.n3118 9.3
R5213 GND.n3118 GND.n3117 9.3
R5214 GND.n3111 GND.n3110 9.3
R5215 GND.n3107 GND.n3106 9.3
R5216 GND.n3106 GND.n3105 9.3
R5217 GND.n3099 GND.n3098 9.3
R5218 GND.n3095 GND.n3094 9.3
R5219 GND.n3094 GND.n3093 9.3
R5220 GND.n3087 GND.n3086 9.3
R5221 GND.n3083 GND.n3082 9.3
R5222 GND.n3082 GND.n3081 9.3
R5223 GND.n3075 GND.n3074 9.3
R5224 GND.n3071 GND.n3070 9.3
R5225 GND.n3070 GND.n3069 9.3
R5226 GND.n3063 GND.n3062 9.3
R5227 GND.n3062 GND.n3061 9.3
R5228 GND.n3053 GND.n3052 9.3
R5229 GND.n3051 GND.n3050 9.3
R5230 GND.n3050 GND.n3049 9.3
R5231 GND.n3041 GND.n3040 9.3
R5232 GND.n3039 GND.n3038 9.3
R5233 GND.n3038 GND.n3037 9.3
R5234 GND.n3029 GND.n3028 9.3
R5235 GND.n3027 GND.n3026 9.3
R5236 GND.n3026 GND.n3025 9.3
R5237 GND.n3017 GND.n3016 9.3
R5238 GND.n3015 GND.n3014 9.3
R5239 GND.n3014 GND.n3013 9.3
R5240 GND.n3005 GND.n3004 9.3
R5241 GND.n3003 GND.n3002 9.3
R5242 GND.n3002 GND.n3001 9.3
R5243 GND.n2993 GND.n2992 9.3
R5244 GND.n2991 GND.n2990 9.3
R5245 GND.n2990 GND.n2989 9.3
R5246 GND.n2981 GND.n2980 9.3
R5247 GND.n3144 GND.n3143 9.3
R5248 GND.n3148 GND.n3147 9.3
R5249 GND.n3182 GND.n3181 9.3
R5250 GND.n3191 GND.n3190 9.3
R5251 GND.n3336 GND.n3335 9.3
R5252 GND.n3332 GND.n3331 9.3
R5253 GND.n3331 GND.n3330 9.3
R5254 GND.n3323 GND.n3322 9.3
R5255 GND.n3319 GND.n3318 9.3
R5256 GND.n3318 GND.n3317 9.3
R5257 GND.n3311 GND.n3310 9.3
R5258 GND.n3307 GND.n3306 9.3
R5259 GND.n3306 GND.n3305 9.3
R5260 GND.n3299 GND.n3298 9.3
R5261 GND.n3295 GND.n3294 9.3
R5262 GND.n3294 GND.n3293 9.3
R5263 GND.n3287 GND.n3286 9.3
R5264 GND.n3283 GND.n3282 9.3
R5265 GND.n3282 GND.n3281 9.3
R5266 GND.n3275 GND.n3274 9.3
R5267 GND.n3271 GND.n3270 9.3
R5268 GND.n3270 GND.n3269 9.3
R5269 GND.n3263 GND.n3262 9.3
R5270 GND.n3262 GND.n3261 9.3
R5271 GND.n3253 GND.n3252 9.3
R5272 GND.n3251 GND.n3250 9.3
R5273 GND.n3250 GND.n3249 9.3
R5274 GND.n3241 GND.n3240 9.3
R5275 GND.n3239 GND.n3238 9.3
R5276 GND.n3238 GND.n3237 9.3
R5277 GND.n3229 GND.n3228 9.3
R5278 GND.n3227 GND.n3226 9.3
R5279 GND.n3226 GND.n3225 9.3
R5280 GND.n3217 GND.n3216 9.3
R5281 GND.n3215 GND.n3214 9.3
R5282 GND.n3214 GND.n3213 9.3
R5283 GND.n3205 GND.n3204 9.3
R5284 GND.n3203 GND.n3202 9.3
R5285 GND.n3202 GND.n3201 9.3
R5286 GND.n3193 GND.n3192 9.3
R5287 GND.n3345 GND.n3344 9.3
R5288 GND.n3344 GND.n3343 9.3
R5289 GND.n3349 GND.n3348 9.3
R5290 GND.n14911 GND.n14910 9.3
R5291 GND.n14899 GND.n14898 9.3
R5292 GND.n14886 GND.n14885 9.3
R5293 GND.n14874 GND.n14873 9.3
R5294 GND.n14861 GND.n14860 9.3
R5295 GND.n14849 GND.n14848 9.3
R5296 GND.n14836 GND.n14835 9.3
R5297 GND.n14817 GND.n14816 9.3
R5298 GND.n14804 GND.n14803 9.3
R5299 GND.n14792 GND.n14791 9.3
R5300 GND.n14779 GND.n14778 9.3
R5301 GND.n14767 GND.n14766 9.3
R5302 GND.n14754 GND.n14753 9.3
R5303 GND.n14752 GND.n14751 9.3
R5304 GND.n14763 GND.n14762 9.3
R5305 GND.n14762 GND.n14761 9.3
R5306 GND.n14765 GND.n14764 9.3
R5307 GND.n14775 GND.n14774 9.3
R5308 GND.n14774 GND.n14773 9.3
R5309 GND.n14777 GND.n14776 9.3
R5310 GND.n14788 GND.n14787 9.3
R5311 GND.n14787 GND.n14786 9.3
R5312 GND.n14790 GND.n14789 9.3
R5313 GND.n14800 GND.n14799 9.3
R5314 GND.n14799 GND.n14798 9.3
R5315 GND.n14802 GND.n14801 9.3
R5316 GND.n14813 GND.n14812 9.3
R5317 GND.n14812 GND.n14811 9.3
R5318 GND.n14815 GND.n14814 9.3
R5319 GND.n14826 GND.n14825 9.3
R5320 GND.n14825 GND.n14824 9.3
R5321 GND.n14834 GND.n14833 9.3
R5322 GND.n14833 GND.n14832 9.3
R5323 GND.n14838 GND.n14837 9.3
R5324 GND.n14847 GND.n14846 9.3
R5325 GND.n14846 GND.n14845 9.3
R5326 GND.n14851 GND.n14850 9.3
R5327 GND.n14859 GND.n14858 9.3
R5328 GND.n14858 GND.n14857 9.3
R5329 GND.n14863 GND.n14862 9.3
R5330 GND.n14872 GND.n14871 9.3
R5331 GND.n14871 GND.n14870 9.3
R5332 GND.n14876 GND.n14875 9.3
R5333 GND.n14884 GND.n14883 9.3
R5334 GND.n14883 GND.n14882 9.3
R5335 GND.n14888 GND.n14887 9.3
R5336 GND.n14897 GND.n14896 9.3
R5337 GND.n14896 GND.n14895 9.3
R5338 GND.n14901 GND.n14900 9.3
R5339 GND.n14909 GND.n14908 9.3
R5340 GND.n14908 GND.n14907 9.3
R5341 GND.n14913 GND.n14912 9.3
R5342 GND.n14750 GND.n14749 9.3
R5343 GND.n14749 GND.n14748 9.3
R5344 GND.n14739 GND.n14738 9.3
R5345 GND.n14741 GND.n14740 9.3
R5346 GND.n10415 GND.n10414 9.3
R5347 GND.n10414 GND.n10413 9.3
R5348 GND.n10427 GND.n10426 9.3
R5349 GND.n10426 GND.n10425 9.3
R5350 GND.n10431 GND.n10430 9.3
R5351 GND.n10443 GND.n10442 9.3
R5352 GND.n10455 GND.n10454 9.3
R5353 GND.n10467 GND.n10466 9.3
R5354 GND.n10479 GND.n10478 9.3
R5355 GND.n10497 GND.n10496 9.3
R5356 GND.n10509 GND.n10508 9.3
R5357 GND.n10521 GND.n10520 9.3
R5358 GND.n10533 GND.n10532 9.3
R5359 GND.n10545 GND.n10544 9.3
R5360 GND.n10557 GND.n10556 9.3
R5361 GND.n10429 GND.n10428 9.3
R5362 GND.n10439 GND.n10438 9.3
R5363 GND.n10438 GND.n10437 9.3
R5364 GND.n10441 GND.n10440 9.3
R5365 GND.n10451 GND.n10450 9.3
R5366 GND.n10450 GND.n10449 9.3
R5367 GND.n10453 GND.n10452 9.3
R5368 GND.n10463 GND.n10462 9.3
R5369 GND.n10462 GND.n10461 9.3
R5370 GND.n10465 GND.n10464 9.3
R5371 GND.n10475 GND.n10474 9.3
R5372 GND.n10474 GND.n10473 9.3
R5373 GND.n10477 GND.n10476 9.3
R5374 GND.n10487 GND.n10486 9.3
R5375 GND.n10486 GND.n10485 9.3
R5376 GND.n10495 GND.n10494 9.3
R5377 GND.n10494 GND.n10493 9.3
R5378 GND.n10499 GND.n10498 9.3
R5379 GND.n10507 GND.n10506 9.3
R5380 GND.n10506 GND.n10505 9.3
R5381 GND.n10511 GND.n10510 9.3
R5382 GND.n10519 GND.n10518 9.3
R5383 GND.n10518 GND.n10517 9.3
R5384 GND.n10523 GND.n10522 9.3
R5385 GND.n10531 GND.n10530 9.3
R5386 GND.n10530 GND.n10529 9.3
R5387 GND.n10535 GND.n10534 9.3
R5388 GND.n10543 GND.n10542 9.3
R5389 GND.n10542 GND.n10541 9.3
R5390 GND.n10547 GND.n10546 9.3
R5391 GND.n10555 GND.n10554 9.3
R5392 GND.n10554 GND.n10553 9.3
R5393 GND.n10559 GND.n10558 9.3
R5394 GND.n10568 GND.n10567 9.3
R5395 GND.n10567 GND.n10566 9.3
R5396 GND.n10566 GND.n10565 9.3
R5397 GND.n10572 GND.n10571 9.3
R5398 GND.n10570 GND.n10569 9.3
R5399 GND.n10395 GND.n10394 9.3
R5400 GND.n10407 GND.n10406 9.3
R5401 GND.n10419 GND.n10418 9.3
R5402 GND.n10417 GND.n10416 9.3
R5403 GND.n14084 GND.n14083 9.3
R5404 GND.n14094 GND.n14093 9.3
R5405 GND.n14093 GND.n14092 9.3
R5406 GND.n14086 GND.n14085 9.3
R5407 GND.n14111 GND.n14110 9.3
R5408 GND.n14110 GND.n14109 9.3
R5409 GND.n14118 GND.n14117 9.3
R5410 GND.n14113 GND.n14112 9.3
R5411 GND.n15549 GND.n15548 9.3
R5412 GND.n15561 GND.n15560 9.3
R5413 GND.n15574 GND.n15573 9.3
R5414 GND.n15586 GND.n15585 9.3
R5415 GND.n15599 GND.n15598 9.3
R5416 GND.n15611 GND.n15610 9.3
R5417 GND.n15624 GND.n15623 9.3
R5418 GND.n15643 GND.n15642 9.3
R5419 GND.n15656 GND.n15655 9.3
R5420 GND.n15668 GND.n15667 9.3
R5421 GND.n15681 GND.n15680 9.3
R5422 GND.n15693 GND.n15692 9.3
R5423 GND.n15706 GND.n15705 9.3
R5424 GND.n15547 GND.n15546 9.3
R5425 GND.n15557 GND.n15556 9.3
R5426 GND.n15556 GND.n15555 9.3
R5427 GND.n15708 GND.n15707 9.3
R5428 GND.n15704 GND.n15703 9.3
R5429 GND.n15703 GND.n15702 9.3
R5430 GND.n15695 GND.n15694 9.3
R5431 GND.n15691 GND.n15690 9.3
R5432 GND.n15690 GND.n15689 9.3
R5433 GND.n15683 GND.n15682 9.3
R5434 GND.n15679 GND.n15678 9.3
R5435 GND.n15678 GND.n15677 9.3
R5436 GND.n15670 GND.n15669 9.3
R5437 GND.n15666 GND.n15665 9.3
R5438 GND.n15665 GND.n15664 9.3
R5439 GND.n15658 GND.n15657 9.3
R5440 GND.n15654 GND.n15653 9.3
R5441 GND.n15653 GND.n15652 9.3
R5442 GND.n15645 GND.n15644 9.3
R5443 GND.n15641 GND.n15640 9.3
R5444 GND.n15640 GND.n15639 9.3
R5445 GND.n15632 GND.n15631 9.3
R5446 GND.n15631 GND.n15630 9.3
R5447 GND.n15622 GND.n15621 9.3
R5448 GND.n15620 GND.n15619 9.3
R5449 GND.n15619 GND.n15618 9.3
R5450 GND.n15609 GND.n15608 9.3
R5451 GND.n15607 GND.n15606 9.3
R5452 GND.n15606 GND.n15605 9.3
R5453 GND.n15597 GND.n15596 9.3
R5454 GND.n15595 GND.n15594 9.3
R5455 GND.n15594 GND.n15593 9.3
R5456 GND.n15584 GND.n15583 9.3
R5457 GND.n15582 GND.n15581 9.3
R5458 GND.n15581 GND.n15580 9.3
R5459 GND.n15572 GND.n15571 9.3
R5460 GND.n15570 GND.n15569 9.3
R5461 GND.n15569 GND.n15568 9.3
R5462 GND.n15559 GND.n15558 9.3
R5463 GND.n15716 GND.n15715 9.3
R5464 GND.n15728 GND.n15727 9.3
R5465 GND.n15749 GND.n15748 9.3
R5466 GND.n15752 GND.n15751 9.3
R5467 GND.n15747 GND.n15746 9.3
R5468 GND.n15746 GND.n15745 9.3
R5469 GND.n15736 GND.n15735 9.3
R5470 GND.n15735 GND.n15734 9.3
R5471 GND.n15725 GND.n15724 9.3
R5472 GND.n15869 GND.n15868 9.3
R5473 GND.n15862 GND.n15861 9.3
R5474 GND.n15855 GND.n15854 9.3
R5475 GND.n15848 GND.n15847 9.3
R5476 GND.n15841 GND.n15840 9.3
R5477 GND.n15834 GND.n15833 9.3
R5478 GND.n15827 GND.n15826 9.3
R5479 GND.n15820 GND.n15819 9.3
R5480 GND.n15800 GND.n15799 9.3
R5481 GND.n15792 GND.n15791 9.3
R5482 GND.n15802 GND.n15801 9.3
R5483 GND.n15796 GND.n15795 9.3
R5484 GND.n15790 GND.n15789 9.3
R5485 GND.n15786 GND.n15785 9.3
R5486 GND.n15813 GND.n15812 9.3
R5487 GND.n15818 GND.n15817 9.3
R5488 GND.n15823 GND.n15822 9.3
R5489 GND.n15825 GND.n15824 9.3
R5490 GND.n15830 GND.n15829 9.3
R5491 GND.n15832 GND.n15831 9.3
R5492 GND.n15837 GND.n15836 9.3
R5493 GND.n15839 GND.n15838 9.3
R5494 GND.n15844 GND.n15843 9.3
R5495 GND.n15846 GND.n15845 9.3
R5496 GND.n15851 GND.n15850 9.3
R5497 GND.n15853 GND.n15852 9.3
R5498 GND.n15858 GND.n15857 9.3
R5499 GND.n15860 GND.n15859 9.3
R5500 GND.n15865 GND.n15864 9.3
R5501 GND.n15867 GND.n15866 9.3
R5502 GND.n15871 GND.n15870 9.3
R5503 GND.n15773 GND.n15772 9.3
R5504 GND.n15769 GND.n15768 9.3
R5505 GND.n15765 GND.n15764 9.3
R5506 GND.n15761 GND.n15760 9.3
R5507 GND.n15777 GND.n15776 9.3
R5508 GND.n15780 GND.n15779 9.3
R5509 GND.n15782 GND.n15781 9.3
R5510 GND.n15422 GND.n15421 9.3
R5511 GND.n15417 GND.n15416 9.3
R5512 GND.n15410 GND.n15409 9.3
R5513 GND.n15403 GND.n15402 9.3
R5514 GND.n15396 GND.n15395 9.3
R5515 GND.n15389 GND.n15388 9.3
R5516 GND.n15382 GND.n15381 9.3
R5517 GND.n15375 GND.n15374 9.3
R5518 GND.n15354 GND.n15353 9.3
R5519 GND.n15346 GND.n15345 9.3
R5520 GND.n15420 GND.n15419 9.3
R5521 GND.n15415 GND.n15414 9.3
R5522 GND.n15413 GND.n15412 9.3
R5523 GND.n15408 GND.n15407 9.3
R5524 GND.n15406 GND.n15405 9.3
R5525 GND.n15401 GND.n15400 9.3
R5526 GND.n15399 GND.n15398 9.3
R5527 GND.n15394 GND.n15393 9.3
R5528 GND.n15392 GND.n15391 9.3
R5529 GND.n15387 GND.n15386 9.3
R5530 GND.n15385 GND.n15384 9.3
R5531 GND.n15380 GND.n15379 9.3
R5532 GND.n15378 GND.n15377 9.3
R5533 GND.n15373 GND.n15372 9.3
R5534 GND.n15368 GND.n15367 9.3
R5535 GND.n15356 GND.n15355 9.3
R5536 GND.n15350 GND.n15349 9.3
R5537 GND.n15344 GND.n15343 9.3
R5538 GND.n15340 GND.n15339 9.3
R5539 GND.n15424 GND.n15423 9.3
R5540 GND.n15426 GND.n15425 9.3
R5541 GND.n15327 GND.n15326 9.3
R5542 GND.n15323 GND.n15322 9.3
R5543 GND.n15319 GND.n15318 9.3
R5544 GND.n15315 GND.n15314 9.3
R5545 GND.n15331 GND.n15330 9.3
R5546 GND.n15334 GND.n15333 9.3
R5547 GND.n15336 GND.n15335 9.3
R5548 GND.n14926 GND.n14925 9.3
R5549 GND.n14931 GND.n14930 9.3
R5550 GND.n14938 GND.n14937 9.3
R5551 GND.n14945 GND.n14944 9.3
R5552 GND.n14952 GND.n14951 9.3
R5553 GND.n14959 GND.n14958 9.3
R5554 GND.n14966 GND.n14965 9.3
R5555 GND.n14973 GND.n14972 9.3
R5556 GND.n14422 GND.n14421 9.3
R5557 GND.n14430 GND.n14429 9.3
R5558 GND.n14929 GND.n14928 9.3
R5559 GND.n14933 GND.n14932 9.3
R5560 GND.n14936 GND.n14935 9.3
R5561 GND.n14940 GND.n14939 9.3
R5562 GND.n14943 GND.n14942 9.3
R5563 GND.n14947 GND.n14946 9.3
R5564 GND.n14950 GND.n14949 9.3
R5565 GND.n14954 GND.n14953 9.3
R5566 GND.n14957 GND.n14956 9.3
R5567 GND.n14961 GND.n14960 9.3
R5568 GND.n14964 GND.n14963 9.3
R5569 GND.n14968 GND.n14967 9.3
R5570 GND.n14971 GND.n14970 9.3
R5571 GND.n14976 GND.n14975 9.3
R5572 GND.n14980 GND.n14979 9.3
R5573 GND.n14420 GND.n14419 9.3
R5574 GND.n14427 GND.n14426 9.3
R5575 GND.n14432 GND.n14431 9.3
R5576 GND.n14437 GND.n14436 9.3
R5577 GND.n14924 GND.n14923 9.3
R5578 GND.n14922 GND.n14921 9.3
R5579 GND.n14450 GND.n14449 9.3
R5580 GND.n14456 GND.n14455 9.3
R5581 GND.n14459 GND.n14458 9.3
R5582 GND.n14463 GND.n14462 9.3
R5583 GND.n14447 GND.n14446 9.3
R5584 GND.n14442 GND.n14441 9.3
R5585 GND.n14440 GND.n14439 9.3
R5586 GND.n14478 GND.n14477 9.3
R5587 GND.n14486 GND.n14485 9.3
R5588 GND.n14485 GND.n14484 9.3
R5589 GND.n14488 GND.n14487 9.3
R5590 GND.n15437 GND.n15436 9.3
R5591 GND.n15436 GND.n15435 9.3
R5592 GND.n15446 GND.n15445 9.3
R5593 GND.n15439 GND.n15438 9.3
R5594 GND.n15108 GND.n15107 9.3
R5595 GND.n15103 GND.n15102 9.3
R5596 GND.n15096 GND.n15095 9.3
R5597 GND.n15089 GND.n15088 9.3
R5598 GND.n15082 GND.n15081 9.3
R5599 GND.n15075 GND.n15074 9.3
R5600 GND.n15068 GND.n15067 9.3
R5601 GND.n15061 GND.n15060 9.3
R5602 GND.n15046 GND.n15045 9.3
R5603 GND.n15038 GND.n15037 9.3
R5604 GND.n15106 GND.n15105 9.3
R5605 GND.n15101 GND.n15100 9.3
R5606 GND.n15099 GND.n15098 9.3
R5607 GND.n15094 GND.n15093 9.3
R5608 GND.n15092 GND.n15091 9.3
R5609 GND.n15087 GND.n15086 9.3
R5610 GND.n15085 GND.n15084 9.3
R5611 GND.n15080 GND.n15079 9.3
R5612 GND.n15078 GND.n15077 9.3
R5613 GND.n15073 GND.n15072 9.3
R5614 GND.n15071 GND.n15070 9.3
R5615 GND.n15066 GND.n15065 9.3
R5616 GND.n15064 GND.n15063 9.3
R5617 GND.n15059 GND.n15058 9.3
R5618 GND.n15054 GND.n15053 9.3
R5619 GND.n15048 GND.n15047 9.3
R5620 GND.n15042 GND.n15041 9.3
R5621 GND.n15036 GND.n15035 9.3
R5622 GND.n15032 GND.n15031 9.3
R5623 GND.n15110 GND.n15109 9.3
R5624 GND.n15112 GND.n15111 9.3
R5625 GND.n15019 GND.n15018 9.3
R5626 GND.n15015 GND.n15014 9.3
R5627 GND.n15011 GND.n15010 9.3
R5628 GND.n15007 GND.n15006 9.3
R5629 GND.n15023 GND.n15022 9.3
R5630 GND.n15026 GND.n15025 9.3
R5631 GND.n15028 GND.n15027 9.3
R5632 GND.n15298 GND.n15297 9.3
R5633 GND.n14474 GND.n14473 9.3
R5634 GND.n14719 GND.n14718 9.3
R5635 GND.n14472 GND.n14471 9.3
R5636 GND.n14471 GND.n14470 9.3
R5637 GND.n15305 GND.n15304 9.3
R5638 GND.n15304 GND.n15303 9.3
R5639 GND.n15296 GND.n15295 9.3
R5640 GND.n15275 GND.n15274 9.3
R5641 GND.n15274 GND.n15273 9.3
R5642 GND.n15267 GND.n15266 9.3
R5643 GND.n15253 GND.n15252 9.3
R5644 GND.n15240 GND.n15239 9.3
R5645 GND.n15228 GND.n15227 9.3
R5646 GND.n15216 GND.n15215 9.3
R5647 GND.n15204 GND.n15203 9.3
R5648 GND.n15186 GND.n15185 9.3
R5649 GND.n15174 GND.n15173 9.3
R5650 GND.n15162 GND.n15161 9.3
R5651 GND.n15150 GND.n15149 9.3
R5652 GND.n15138 GND.n15137 9.3
R5653 GND.n15126 GND.n15125 9.3
R5654 GND.n15255 GND.n15254 9.3
R5655 GND.n15251 GND.n15250 9.3
R5656 GND.n15250 GND.n15249 9.3
R5657 GND.n15242 GND.n15241 9.3
R5658 GND.n15238 GND.n15237 9.3
R5659 GND.n15237 GND.n15236 9.3
R5660 GND.n15230 GND.n15229 9.3
R5661 GND.n15226 GND.n15225 9.3
R5662 GND.n15225 GND.n15224 9.3
R5663 GND.n15218 GND.n15217 9.3
R5664 GND.n15214 GND.n15213 9.3
R5665 GND.n15213 GND.n15212 9.3
R5666 GND.n15206 GND.n15205 9.3
R5667 GND.n15202 GND.n15201 9.3
R5668 GND.n15201 GND.n15200 9.3
R5669 GND.n15194 GND.n15193 9.3
R5670 GND.n15193 GND.n15192 9.3
R5671 GND.n15184 GND.n15183 9.3
R5672 GND.n15182 GND.n15181 9.3
R5673 GND.n15181 GND.n15180 9.3
R5674 GND.n15172 GND.n15171 9.3
R5675 GND.n15170 GND.n15169 9.3
R5676 GND.n15169 GND.n15168 9.3
R5677 GND.n15160 GND.n15159 9.3
R5678 GND.n15158 GND.n15157 9.3
R5679 GND.n15157 GND.n15156 9.3
R5680 GND.n15148 GND.n15147 9.3
R5681 GND.n15146 GND.n15145 9.3
R5682 GND.n15145 GND.n15144 9.3
R5683 GND.n15136 GND.n15135 9.3
R5684 GND.n15134 GND.n15133 9.3
R5685 GND.n15133 GND.n15132 9.3
R5686 GND.n15124 GND.n15123 9.3
R5687 GND.n15121 GND.n15120 9.3
R5688 GND.n15265 GND.n15264 9.3
R5689 GND.n15263 GND.n15262 9.3
R5690 GND.n15262 GND.n15261 9.3
R5691 GND.n15277 GND.n15276 9.3
R5692 GND.n15279 GND.n15278 9.3
R5693 GND.n3949 GND.n3948 9.3
R5694 GND.n3948 GND.n3947 9.3
R5695 GND.n3947 GND.n3946 9.3
R5696 GND.n3906 GND.n3905 9.3
R5697 GND.n3894 GND.n3893 9.3
R5698 GND.n3882 GND.n3881 9.3
R5699 GND.n3870 GND.n3869 9.3
R5700 GND.n3858 GND.n3857 9.3
R5701 GND.n3836 GND.n3835 9.3
R5702 GND.n3828 GND.n3827 9.3
R5703 GND.n3820 GND.n3819 9.3
R5704 GND.n3812 GND.n3811 9.3
R5705 GND.n3804 GND.n3803 9.3
R5706 GND.n3796 GND.n3795 9.3
R5707 GND.n3788 GND.n3787 9.3
R5708 GND.n3782 GND.n3781 9.3
R5709 GND.n3777 GND.n3776 9.3
R5710 GND.n3772 GND.n3771 9.3
R5711 GND.n3753 GND.n3752 9.3
R5712 GND.n3735 GND.n3734 9.3
R5713 GND.n3723 GND.n3722 9.3
R5714 GND.n3711 GND.n3710 9.3
R5715 GND.n3699 GND.n3698 9.3
R5716 GND.n3687 GND.n3686 9.3
R5717 GND.n3674 GND.n3673 9.3
R5718 GND.n3672 GND.n3671 9.3
R5719 GND.n3683 GND.n3682 9.3
R5720 GND.n3682 GND.n3681 9.3
R5721 GND.n3685 GND.n3684 9.3
R5722 GND.n3695 GND.n3694 9.3
R5723 GND.n3694 GND.n3693 9.3
R5724 GND.n3697 GND.n3696 9.3
R5725 GND.n3707 GND.n3706 9.3
R5726 GND.n3706 GND.n3705 9.3
R5727 GND.n3709 GND.n3708 9.3
R5728 GND.n3719 GND.n3718 9.3
R5729 GND.n3718 GND.n3717 9.3
R5730 GND.n3721 GND.n3720 9.3
R5731 GND.n3731 GND.n3730 9.3
R5732 GND.n3730 GND.n3729 9.3
R5733 GND.n3733 GND.n3732 9.3
R5734 GND.n3743 GND.n3742 9.3
R5735 GND.n3742 GND.n3741 9.3
R5736 GND.n3751 GND.n3750 9.3
R5737 GND.n3750 GND.n3749 9.3
R5738 GND.n3755 GND.n3754 9.3
R5739 GND.n3759 GND.n3758 9.3
R5740 GND.n3641 GND.n3640 9.3
R5741 GND.n3765 GND.n3764 9.3
R5742 GND.n3653 GND.n3652 9.3
R5743 GND.n3769 GND.n3768 9.3
R5744 GND.n3634 GND.n3633 9.3
R5745 GND.n3774 GND.n3773 9.3
R5746 GND.n3660 GND.n3659 9.3
R5747 GND.n3779 GND.n3778 9.3
R5748 GND.n3627 GND.n3626 9.3
R5749 GND.n3784 GND.n3783 9.3
R5750 GND.n3786 GND.n3785 9.3
R5751 GND.n3792 GND.n3791 9.3
R5752 GND.n3946 GND.n3933 9.3
R5753 GND.n3794 GND.n3793 9.3
R5754 GND.n3800 GND.n3799 9.3
R5755 GND.n3946 GND.n3937 9.3
R5756 GND.n3802 GND.n3801 9.3
R5757 GND.n3808 GND.n3807 9.3
R5758 GND.n3946 GND.n3929 9.3
R5759 GND.n3810 GND.n3809 9.3
R5760 GND.n3816 GND.n3815 9.3
R5761 GND.n3946 GND.n3941 9.3
R5762 GND.n3818 GND.n3817 9.3
R5763 GND.n3824 GND.n3823 9.3
R5764 GND.n3946 GND.n3925 9.3
R5765 GND.n3826 GND.n3825 9.3
R5766 GND.n3832 GND.n3831 9.3
R5767 GND.n3946 GND.n3945 9.3
R5768 GND.n3834 GND.n3833 9.3
R5769 GND.n3840 GND.n3839 9.3
R5770 GND.n3946 GND.n3921 9.3
R5771 GND.n3856 GND.n3855 9.3
R5772 GND.n3855 GND.n3854 9.3
R5773 GND.n3860 GND.n3859 9.3
R5774 GND.n3868 GND.n3867 9.3
R5775 GND.n3867 GND.n3866 9.3
R5776 GND.n3872 GND.n3871 9.3
R5777 GND.n3880 GND.n3879 9.3
R5778 GND.n3879 GND.n3878 9.3
R5779 GND.n3884 GND.n3883 9.3
R5780 GND.n3892 GND.n3891 9.3
R5781 GND.n3891 GND.n3890 9.3
R5782 GND.n3896 GND.n3895 9.3
R5783 GND.n3904 GND.n3903 9.3
R5784 GND.n3903 GND.n3902 9.3
R5785 GND.n3908 GND.n3907 9.3
R5786 GND.n3670 GND.n3669 9.3
R5787 GND.n3669 GND.n3668 9.3
R5788 GND.n1917 GND.n1916 9.3
R5789 GND.n3621 GND.n3620 9.3
R5790 GND.n3951 GND.n3950 9.3
R5791 GND.n3953 GND.n3952 9.3
R5792 GND.n5787 GND.n5786 9.3
R5793 GND.n5786 GND.n5785 9.3
R5794 GND.n5785 GND.n5784 9.3
R5795 GND.n5744 GND.n5743 9.3
R5796 GND.n5732 GND.n5731 9.3
R5797 GND.n5720 GND.n5719 9.3
R5798 GND.n5708 GND.n5707 9.3
R5799 GND.n5696 GND.n5695 9.3
R5800 GND.n5674 GND.n5673 9.3
R5801 GND.n5666 GND.n5665 9.3
R5802 GND.n5658 GND.n5657 9.3
R5803 GND.n5650 GND.n5649 9.3
R5804 GND.n5642 GND.n5641 9.3
R5805 GND.n5634 GND.n5633 9.3
R5806 GND.n5626 GND.n5625 9.3
R5807 GND.n5620 GND.n5619 9.3
R5808 GND.n5615 GND.n5614 9.3
R5809 GND.n5610 GND.n5609 9.3
R5810 GND.n5591 GND.n5590 9.3
R5811 GND.n5572 GND.n5571 9.3
R5812 GND.n5559 GND.n5558 9.3
R5813 GND.n5547 GND.n5546 9.3
R5814 GND.n5534 GND.n5533 9.3
R5815 GND.n5522 GND.n5521 9.3
R5816 GND.n5509 GND.n5508 9.3
R5817 GND.n5507 GND.n5506 9.3
R5818 GND.n5518 GND.n5517 9.3
R5819 GND.n5517 GND.n5516 9.3
R5820 GND.n5520 GND.n5519 9.3
R5821 GND.n5530 GND.n5529 9.3
R5822 GND.n5529 GND.n5528 9.3
R5823 GND.n5532 GND.n5531 9.3
R5824 GND.n5543 GND.n5542 9.3
R5825 GND.n5542 GND.n5541 9.3
R5826 GND.n5545 GND.n5544 9.3
R5827 GND.n5555 GND.n5554 9.3
R5828 GND.n5554 GND.n5553 9.3
R5829 GND.n5557 GND.n5556 9.3
R5830 GND.n5568 GND.n5567 9.3
R5831 GND.n5567 GND.n5566 9.3
R5832 GND.n5570 GND.n5569 9.3
R5833 GND.n5581 GND.n5580 9.3
R5834 GND.n5580 GND.n5579 9.3
R5835 GND.n5589 GND.n5588 9.3
R5836 GND.n5588 GND.n5587 9.3
R5837 GND.n5593 GND.n5592 9.3
R5838 GND.n5597 GND.n5596 9.3
R5839 GND.n5492 GND.n5491 9.3
R5840 GND.n5603 GND.n5602 9.3
R5841 GND.n5487 GND.n5486 9.3
R5842 GND.n5607 GND.n5606 9.3
R5843 GND.n5476 GND.n5475 9.3
R5844 GND.n5612 GND.n5611 9.3
R5845 GND.n5471 GND.n5470 9.3
R5846 GND.n5617 GND.n5616 9.3
R5847 GND.n5461 GND.n5460 9.3
R5848 GND.n5622 GND.n5621 9.3
R5849 GND.n5624 GND.n5623 9.3
R5850 GND.n5630 GND.n5629 9.3
R5851 GND.n5784 GND.n5771 9.3
R5852 GND.n5632 GND.n5631 9.3
R5853 GND.n5638 GND.n5637 9.3
R5854 GND.n5784 GND.n5775 9.3
R5855 GND.n5640 GND.n5639 9.3
R5856 GND.n5646 GND.n5645 9.3
R5857 GND.n5784 GND.n5767 9.3
R5858 GND.n5648 GND.n5647 9.3
R5859 GND.n5654 GND.n5653 9.3
R5860 GND.n5784 GND.n5779 9.3
R5861 GND.n5656 GND.n5655 9.3
R5862 GND.n5662 GND.n5661 9.3
R5863 GND.n5784 GND.n5763 9.3
R5864 GND.n5664 GND.n5663 9.3
R5865 GND.n5670 GND.n5669 9.3
R5866 GND.n5784 GND.n5783 9.3
R5867 GND.n5672 GND.n5671 9.3
R5868 GND.n5678 GND.n5677 9.3
R5869 GND.n5784 GND.n5759 9.3
R5870 GND.n5694 GND.n5693 9.3
R5871 GND.n5693 GND.n5692 9.3
R5872 GND.n5698 GND.n5697 9.3
R5873 GND.n5706 GND.n5705 9.3
R5874 GND.n5705 GND.n5704 9.3
R5875 GND.n5710 GND.n5709 9.3
R5876 GND.n5718 GND.n5717 9.3
R5877 GND.n5717 GND.n5716 9.3
R5878 GND.n5722 GND.n5721 9.3
R5879 GND.n5730 GND.n5729 9.3
R5880 GND.n5729 GND.n5728 9.3
R5881 GND.n5734 GND.n5733 9.3
R5882 GND.n5742 GND.n5741 9.3
R5883 GND.n5741 GND.n5740 9.3
R5884 GND.n5746 GND.n5745 9.3
R5885 GND.n5505 GND.n5504 9.3
R5886 GND.n5504 GND.n5503 9.3
R5887 GND.n5451 GND.n5450 9.3
R5888 GND.n5453 GND.n5452 9.3
R5889 GND.n5789 GND.n5788 9.3
R5890 GND.n5791 GND.n5790 9.3
R5891 GND.n16434 GND.n16433 9.3
R5892 GND.n16423 GND.n16422 9.3
R5893 GND.n16458 GND.n16457 9.3
R5894 GND.n16446 GND.n16445 9.3
R5895 GND.n16463 GND.n16462 9.3
R5896 GND.n16467 GND.n16466 9.3
R5897 GND.n16469 GND.n16468 9.3
R5898 GND.n16475 GND.n16474 9.3
R5899 GND.n16456 GND.n16455 9.3
R5900 GND.n16440 GND.n16439 9.3
R5901 GND.n16481 GND.n16480 9.3
R5902 GND.n16479 GND.n16478 9.3
R5903 GND.n16417 GND.n16416 9.3
R5904 GND.n16429 GND.n16428 9.3
R5905 GND.n16550 GND.n16549 9.3
R5906 GND.n16546 GND.n16545 9.3
R5907 GND.n16514 GND.n16513 9.3
R5908 GND.n16516 GND.n16515 9.3
R5909 GND.n16505 GND.n16504 9.3
R5910 GND.n16520 GND.n16519 9.3
R5911 GND.n16500 GND.n16499 9.3
R5912 GND.n16535 GND.n16534 9.3
R5913 GND.n16539 GND.n16538 9.3
R5914 GND.n16541 GND.n16540 9.3
R5915 GND.n16526 GND.n16525 9.3
R5916 GND.n16552 GND.n16551 9.3
R5917 GND.n16560 GND.n16559 9.3
R5918 GND.n16332 GND.n16331 9.3
R5919 GND.n16377 GND.n16376 9.3
R5920 GND.n16375 GND.n16374 9.3
R5921 GND.n16366 GND.n16365 9.3
R5922 GND.n16386 GND.n16385 9.3
R5923 GND.n16371 GND.n16370 9.3
R5924 GND.n16364 GND.n16363 9.3
R5925 GND.n16360 GND.n16359 9.3
R5926 GND.n16338 GND.n16337 9.3
R5927 GND.n16343 GND.n16342 9.3
R5928 GND.n16349 GND.n16348 9.3
R5929 GND.n16353 GND.n16352 9.3
R5930 GND.n16355 GND.n16354 9.3
R5931 GND.n16327 GND.n16326 9.3
R5932 GND.n16695 GND.n16694 9.3
R5933 GND.n16684 GND.n16683 9.3
R5934 GND.n16719 GND.n16718 9.3
R5935 GND.n16707 GND.n16706 9.3
R5936 GND.n16724 GND.n16723 9.3
R5937 GND.n16728 GND.n16727 9.3
R5938 GND.n16730 GND.n16729 9.3
R5939 GND.n16736 GND.n16735 9.3
R5940 GND.n16717 GND.n16716 9.3
R5941 GND.n16701 GND.n16700 9.3
R5942 GND.n16742 GND.n16741 9.3
R5943 GND.n16740 GND.n16739 9.3
R5944 GND.n16678 GND.n16677 9.3
R5945 GND.n16690 GND.n16689 9.3
R5946 GND.n16811 GND.n16810 9.3
R5947 GND.n16807 GND.n16806 9.3
R5948 GND.n16775 GND.n16774 9.3
R5949 GND.n16777 GND.n16776 9.3
R5950 GND.n16766 GND.n16765 9.3
R5951 GND.n16781 GND.n16780 9.3
R5952 GND.n16761 GND.n16760 9.3
R5953 GND.n16796 GND.n16795 9.3
R5954 GND.n16800 GND.n16799 9.3
R5955 GND.n16802 GND.n16801 9.3
R5956 GND.n16787 GND.n16786 9.3
R5957 GND.n16813 GND.n16812 9.3
R5958 GND.n16821 GND.n16820 9.3
R5959 GND.n16593 GND.n16592 9.3
R5960 GND.n16638 GND.n16637 9.3
R5961 GND.n16636 GND.n16635 9.3
R5962 GND.n16627 GND.n16626 9.3
R5963 GND.n16647 GND.n16646 9.3
R5964 GND.n16632 GND.n16631 9.3
R5965 GND.n16625 GND.n16624 9.3
R5966 GND.n16621 GND.n16620 9.3
R5967 GND.n16599 GND.n16598 9.3
R5968 GND.n16604 GND.n16603 9.3
R5969 GND.n16610 GND.n16609 9.3
R5970 GND.n16614 GND.n16613 9.3
R5971 GND.n16616 GND.n16615 9.3
R5972 GND.n16588 GND.n16587 9.3
R5973 GND.n16956 GND.n16955 9.3
R5974 GND.n16945 GND.n16944 9.3
R5975 GND.n16980 GND.n16979 9.3
R5976 GND.n16968 GND.n16967 9.3
R5977 GND.n16985 GND.n16984 9.3
R5978 GND.n16989 GND.n16988 9.3
R5979 GND.n16991 GND.n16990 9.3
R5980 GND.n16997 GND.n16996 9.3
R5981 GND.n16978 GND.n16977 9.3
R5982 GND.n16962 GND.n16961 9.3
R5983 GND.n17003 GND.n17002 9.3
R5984 GND.n17001 GND.n17000 9.3
R5985 GND.n16939 GND.n16938 9.3
R5986 GND.n16951 GND.n16950 9.3
R5987 GND.n17072 GND.n17071 9.3
R5988 GND.n17068 GND.n17067 9.3
R5989 GND.n17036 GND.n17035 9.3
R5990 GND.n17038 GND.n17037 9.3
R5991 GND.n17027 GND.n17026 9.3
R5992 GND.n17042 GND.n17041 9.3
R5993 GND.n17022 GND.n17021 9.3
R5994 GND.n17057 GND.n17056 9.3
R5995 GND.n17061 GND.n17060 9.3
R5996 GND.n17063 GND.n17062 9.3
R5997 GND.n17048 GND.n17047 9.3
R5998 GND.n17074 GND.n17073 9.3
R5999 GND.n17082 GND.n17081 9.3
R6000 GND.n16854 GND.n16853 9.3
R6001 GND.n16899 GND.n16898 9.3
R6002 GND.n16897 GND.n16896 9.3
R6003 GND.n16888 GND.n16887 9.3
R6004 GND.n16908 GND.n16907 9.3
R6005 GND.n16893 GND.n16892 9.3
R6006 GND.n16886 GND.n16885 9.3
R6007 GND.n16882 GND.n16881 9.3
R6008 GND.n16860 GND.n16859 9.3
R6009 GND.n16865 GND.n16864 9.3
R6010 GND.n16871 GND.n16870 9.3
R6011 GND.n16875 GND.n16874 9.3
R6012 GND.n16877 GND.n16876 9.3
R6013 GND.n16849 GND.n16848 9.3
R6014 GND.n17217 GND.n17216 9.3
R6015 GND.n17206 GND.n17205 9.3
R6016 GND.n17241 GND.n17240 9.3
R6017 GND.n17229 GND.n17228 9.3
R6018 GND.n17246 GND.n17245 9.3
R6019 GND.n17250 GND.n17249 9.3
R6020 GND.n17252 GND.n17251 9.3
R6021 GND.n17258 GND.n17257 9.3
R6022 GND.n17239 GND.n17238 9.3
R6023 GND.n17223 GND.n17222 9.3
R6024 GND.n17264 GND.n17263 9.3
R6025 GND.n17262 GND.n17261 9.3
R6026 GND.n17200 GND.n17199 9.3
R6027 GND.n17212 GND.n17211 9.3
R6028 GND.n17333 GND.n17332 9.3
R6029 GND.n17329 GND.n17328 9.3
R6030 GND.n17297 GND.n17296 9.3
R6031 GND.n17299 GND.n17298 9.3
R6032 GND.n17288 GND.n17287 9.3
R6033 GND.n17303 GND.n17302 9.3
R6034 GND.n17283 GND.n17282 9.3
R6035 GND.n17318 GND.n17317 9.3
R6036 GND.n17322 GND.n17321 9.3
R6037 GND.n17324 GND.n17323 9.3
R6038 GND.n17309 GND.n17308 9.3
R6039 GND.n17335 GND.n17334 9.3
R6040 GND.n17343 GND.n17342 9.3
R6041 GND.n17115 GND.n17114 9.3
R6042 GND.n17160 GND.n17159 9.3
R6043 GND.n17158 GND.n17157 9.3
R6044 GND.n17149 GND.n17148 9.3
R6045 GND.n17169 GND.n17168 9.3
R6046 GND.n17154 GND.n17153 9.3
R6047 GND.n17147 GND.n17146 9.3
R6048 GND.n17143 GND.n17142 9.3
R6049 GND.n17121 GND.n17120 9.3
R6050 GND.n17126 GND.n17125 9.3
R6051 GND.n17132 GND.n17131 9.3
R6052 GND.n17136 GND.n17135 9.3
R6053 GND.n17138 GND.n17137 9.3
R6054 GND.n17110 GND.n17109 9.3
R6055 GND.n17478 GND.n17477 9.3
R6056 GND.n17467 GND.n17466 9.3
R6057 GND.n17502 GND.n17501 9.3
R6058 GND.n17490 GND.n17489 9.3
R6059 GND.n17507 GND.n17506 9.3
R6060 GND.n17511 GND.n17510 9.3
R6061 GND.n17513 GND.n17512 9.3
R6062 GND.n17519 GND.n17518 9.3
R6063 GND.n17500 GND.n17499 9.3
R6064 GND.n17484 GND.n17483 9.3
R6065 GND.n17525 GND.n17524 9.3
R6066 GND.n17523 GND.n17522 9.3
R6067 GND.n17461 GND.n17460 9.3
R6068 GND.n17473 GND.n17472 9.3
R6069 GND.n17594 GND.n17593 9.3
R6070 GND.n17590 GND.n17589 9.3
R6071 GND.n17558 GND.n17557 9.3
R6072 GND.n17560 GND.n17559 9.3
R6073 GND.n17549 GND.n17548 9.3
R6074 GND.n17564 GND.n17563 9.3
R6075 GND.n17544 GND.n17543 9.3
R6076 GND.n17579 GND.n17578 9.3
R6077 GND.n17583 GND.n17582 9.3
R6078 GND.n17585 GND.n17584 9.3
R6079 GND.n17570 GND.n17569 9.3
R6080 GND.n17596 GND.n17595 9.3
R6081 GND.n17604 GND.n17603 9.3
R6082 GND.n17376 GND.n17375 9.3
R6083 GND.n17421 GND.n17420 9.3
R6084 GND.n17419 GND.n17418 9.3
R6085 GND.n17410 GND.n17409 9.3
R6086 GND.n17430 GND.n17429 9.3
R6087 GND.n17415 GND.n17414 9.3
R6088 GND.n17408 GND.n17407 9.3
R6089 GND.n17404 GND.n17403 9.3
R6090 GND.n17382 GND.n17381 9.3
R6091 GND.n17387 GND.n17386 9.3
R6092 GND.n17393 GND.n17392 9.3
R6093 GND.n17397 GND.n17396 9.3
R6094 GND.n17399 GND.n17398 9.3
R6095 GND.n17371 GND.n17370 9.3
R6096 GND.n643 GND.n642 9.3
R6097 GND.n640 GND.n639 9.3
R6098 GND.n699 GND.n698 9.3
R6099 GND.n688 GND.n687 9.3
R6100 GND.n694 GND.n693 9.3
R6101 GND.n654 GND.n653 9.3
R6102 GND.n652 GND.n651 9.3
R6103 GND.n663 GND.n662 9.3
R6104 GND.n673 GND.n672 9.3
R6105 GND.n659 GND.n658 9.3
R6106 GND.n665 GND.n664 9.3
R6107 GND.n648 GND.n647 9.3
R6108 GND.n636 GND.n635 9.3
R6109 GND.n766 GND.n765 9.3
R6110 GND.n762 GND.n761 9.3
R6111 GND.n726 GND.n725 9.3
R6112 GND.n750 GND.n749 9.3
R6113 GND.n757 GND.n756 9.3
R6114 GND.n721 GND.n720 9.3
R6115 GND.n714 GND.n713 9.3
R6116 GND.n738 GND.n737 9.3
R6117 GND.n742 GND.n741 9.3
R6118 GND.n745 GND.n744 9.3
R6119 GND.n755 GND.n754 9.3
R6120 GND.n768 GND.n767 9.3
R6121 GND.n776 GND.n775 9.3
R6122 GND.n555 GND.n554 9.3
R6123 GND.n589 GND.n588 9.3
R6124 GND.n607 GND.n606 9.3
R6125 GND.n597 GND.n596 9.3
R6126 GND.n599 GND.n598 9.3
R6127 GND.n594 GND.n593 9.3
R6128 GND.n587 GND.n586 9.3
R6129 GND.n582 GND.n581 9.3
R6130 GND.n561 GND.n560 9.3
R6131 GND.n565 GND.n564 9.3
R6132 GND.n570 GND.n569 9.3
R6133 GND.n574 GND.n573 9.3
R6134 GND.n577 GND.n576 9.3
R6135 GND.n549 GND.n548 9.3
R6136 GND.n385 GND.n384 9.3
R6137 GND.n382 GND.n381 9.3
R6138 GND.n441 GND.n440 9.3
R6139 GND.n430 GND.n429 9.3
R6140 GND.n436 GND.n435 9.3
R6141 GND.n396 GND.n395 9.3
R6142 GND.n394 GND.n393 9.3
R6143 GND.n405 GND.n404 9.3
R6144 GND.n415 GND.n414 9.3
R6145 GND.n401 GND.n400 9.3
R6146 GND.n407 GND.n406 9.3
R6147 GND.n390 GND.n389 9.3
R6148 GND.n378 GND.n377 9.3
R6149 GND.n508 GND.n507 9.3
R6150 GND.n504 GND.n503 9.3
R6151 GND.n468 GND.n467 9.3
R6152 GND.n492 GND.n491 9.3
R6153 GND.n499 GND.n498 9.3
R6154 GND.n463 GND.n462 9.3
R6155 GND.n456 GND.n455 9.3
R6156 GND.n480 GND.n479 9.3
R6157 GND.n484 GND.n483 9.3
R6158 GND.n487 GND.n486 9.3
R6159 GND.n497 GND.n496 9.3
R6160 GND.n510 GND.n509 9.3
R6161 GND.n518 GND.n517 9.3
R6162 GND.n297 GND.n296 9.3
R6163 GND.n331 GND.n330 9.3
R6164 GND.n349 GND.n348 9.3
R6165 GND.n339 GND.n338 9.3
R6166 GND.n341 GND.n340 9.3
R6167 GND.n336 GND.n335 9.3
R6168 GND.n329 GND.n328 9.3
R6169 GND.n324 GND.n323 9.3
R6170 GND.n303 GND.n302 9.3
R6171 GND.n307 GND.n306 9.3
R6172 GND.n312 GND.n311 9.3
R6173 GND.n316 GND.n315 9.3
R6174 GND.n319 GND.n318 9.3
R6175 GND.n291 GND.n290 9.3
R6176 GND.n127 GND.n126 9.3
R6177 GND.n124 GND.n123 9.3
R6178 GND.n183 GND.n182 9.3
R6179 GND.n172 GND.n171 9.3
R6180 GND.n178 GND.n177 9.3
R6181 GND.n138 GND.n137 9.3
R6182 GND.n136 GND.n135 9.3
R6183 GND.n147 GND.n146 9.3
R6184 GND.n157 GND.n156 9.3
R6185 GND.n143 GND.n142 9.3
R6186 GND.n149 GND.n148 9.3
R6187 GND.n132 GND.n131 9.3
R6188 GND.n120 GND.n119 9.3
R6189 GND.n250 GND.n249 9.3
R6190 GND.n246 GND.n245 9.3
R6191 GND.n210 GND.n209 9.3
R6192 GND.n234 GND.n233 9.3
R6193 GND.n241 GND.n240 9.3
R6194 GND.n205 GND.n204 9.3
R6195 GND.n198 GND.n197 9.3
R6196 GND.n222 GND.n221 9.3
R6197 GND.n226 GND.n225 9.3
R6198 GND.n229 GND.n228 9.3
R6199 GND.n239 GND.n238 9.3
R6200 GND.n252 GND.n251 9.3
R6201 GND.n260 GND.n259 9.3
R6202 GND.n39 GND.n38 9.3
R6203 GND.n73 GND.n72 9.3
R6204 GND.n91 GND.n90 9.3
R6205 GND.n81 GND.n80 9.3
R6206 GND.n83 GND.n82 9.3
R6207 GND.n78 GND.n77 9.3
R6208 GND.n71 GND.n70 9.3
R6209 GND.n66 GND.n65 9.3
R6210 GND.n45 GND.n44 9.3
R6211 GND.n49 GND.n48 9.3
R6212 GND.n54 GND.n53 9.3
R6213 GND.n58 GND.n57 9.3
R6214 GND.n61 GND.n60 9.3
R6215 GND.n33 GND.n32 9.3
R6216 GND.n17742 GND.n17741 9.3
R6217 GND.n17739 GND.n17738 9.3
R6218 GND.n17798 GND.n17797 9.3
R6219 GND.n17787 GND.n17786 9.3
R6220 GND.n17793 GND.n17792 9.3
R6221 GND.n17753 GND.n17752 9.3
R6222 GND.n17751 GND.n17750 9.3
R6223 GND.n17762 GND.n17761 9.3
R6224 GND.n17772 GND.n17771 9.3
R6225 GND.n17758 GND.n17757 9.3
R6226 GND.n17764 GND.n17763 9.3
R6227 GND.n17747 GND.n17746 9.3
R6228 GND.n17735 GND.n17734 9.3
R6229 GND.n17839 GND.n17838 9.3
R6230 GND.n17835 GND.n17834 9.3
R6231 GND.n17720 GND.n17719 9.3
R6232 GND.n17823 GND.n17822 9.3
R6233 GND.n17830 GND.n17829 9.3
R6234 GND.n17715 GND.n17714 9.3
R6235 GND.n17708 GND.n17707 9.3
R6236 GND.n17811 GND.n17810 9.3
R6237 GND.n17815 GND.n17814 9.3
R6238 GND.n17818 GND.n17817 9.3
R6239 GND.n17828 GND.n17827 9.3
R6240 GND.n17841 GND.n17840 9.3
R6241 GND.n17849 GND.n17848 9.3
R6242 GND.n17875 GND.n17874 9.3
R6243 GND.n17909 GND.n17908 9.3
R6244 GND.n17927 GND.n17926 9.3
R6245 GND.n17917 GND.n17916 9.3
R6246 GND.n17919 GND.n17918 9.3
R6247 GND.n17914 GND.n17913 9.3
R6248 GND.n17907 GND.n17906 9.3
R6249 GND.n17902 GND.n17901 9.3
R6250 GND.n17881 GND.n17880 9.3
R6251 GND.n17885 GND.n17884 9.3
R6252 GND.n17890 GND.n17889 9.3
R6253 GND.n17894 GND.n17893 9.3
R6254 GND.n17897 GND.n17896 9.3
R6255 GND.n17869 GND.n17868 9.3
R6256 GND.n2813 GND.n2812 9.154
R6257 GND.n2835 GND.n2834 9.154
R6258 GND.n2832 GND.n2831 9.154
R6259 GND.n2829 GND.n2828 9.154
R6260 GND.n2826 GND.n2825 9.154
R6261 GND.n2822 GND.n2821 9.154
R6262 GND.n2819 GND.n2818 9.154
R6263 GND.n2816 GND.n2815 9.154
R6264 GND.n2838 GND.n2837 9.154
R6265 GND.n2679 GND.n2678 9.154
R6266 GND.n2684 GND.n2683 9.154
R6267 GND.n2689 GND.n2688 9.154
R6268 GND.n2694 GND.n2693 9.154
R6269 GND.n2699 GND.n2698 9.154
R6270 GND.n2704 GND.n2703 9.154
R6271 GND.n2707 GND.n2706 9.154
R6272 GND.n2712 GND.n2711 9.154
R6273 GND.n2717 GND.n2716 9.154
R6274 GND.n2722 GND.n2721 9.154
R6275 GND.n2729 GND.n2728 9.154
R6276 GND.n2750 GND.n2749 9.154
R6277 GND.n2753 GND.n2752 9.154
R6278 GND.n2758 GND.n2757 9.154
R6279 GND.n2763 GND.n2762 9.154
R6280 GND.n2768 GND.n2767 9.154
R6281 GND.n2773 GND.n2772 9.154
R6282 GND.n2776 GND.n2775 9.154
R6283 GND.n2781 GND.n2780 9.154
R6284 GND.n2786 GND.n2785 9.154
R6285 GND.n2791 GND.n2790 9.154
R6286 GND.n2796 GND.n2795 9.154
R6287 GND.n2803 GND.n2802 9.154
R6288 GND.n2735 GND.n2734 9.154
R6289 GND.n3963 GND.n3962 9.154
R6290 GND.n3962 GND.n3961 9.154
R6291 GND.n3970 GND.n3969 9.154
R6292 GND.n3969 GND.n3968 9.154
R6293 GND.n3977 GND.n3976 9.154
R6294 GND.n3976 GND.n3975 9.154
R6295 GND.n3984 GND.n3983 9.154
R6296 GND.n3983 GND.n3982 9.154
R6297 GND.n3991 GND.n3990 9.154
R6298 GND.n3990 GND.n3989 9.154
R6299 GND.n4005 GND.n4004 9.154
R6300 GND.n4004 GND.n4003 9.154
R6301 GND.n4012 GND.n4011 9.154
R6302 GND.n4011 GND.n4010 9.154
R6303 GND.n4019 GND.n4018 9.154
R6304 GND.n4018 GND.n4017 9.154
R6305 GND.n4026 GND.n4025 9.154
R6306 GND.n4025 GND.n4024 9.154
R6307 GND.n4033 GND.n4032 9.154
R6308 GND.n4032 GND.n4031 9.154
R6309 GND.n4043 GND.n4042 9.154
R6310 GND.n4042 GND.n4041 9.154
R6311 GND.n4153 GND.n4152 9.154
R6312 GND.n4152 GND.n4151 9.154
R6313 GND.n4143 GND.n4142 9.154
R6314 GND.n4142 GND.n4141 9.154
R6315 GND.n4136 GND.n4135 9.154
R6316 GND.n4135 GND.n4134 9.154
R6317 GND.n4129 GND.n4128 9.154
R6318 GND.n4128 GND.n4127 9.154
R6319 GND.n4122 GND.n4121 9.154
R6320 GND.n4121 GND.n4120 9.154
R6321 GND.n4115 GND.n4114 9.154
R6322 GND.n4114 GND.n4113 9.154
R6323 GND.n4101 GND.n4100 9.154
R6324 GND.n4100 GND.n4099 9.154
R6325 GND.n4094 GND.n4093 9.154
R6326 GND.n4093 GND.n4092 9.154
R6327 GND.n4087 GND.n4086 9.154
R6328 GND.n4086 GND.n4085 9.154
R6329 GND.n4080 GND.n4079 9.154
R6330 GND.n4079 GND.n4078 9.154
R6331 GND.n4073 GND.n4072 9.154
R6332 GND.n4072 GND.n4071 9.154
R6333 GND.n4069 GND.n4068 9.154
R6334 GND.n4068 GND.n4067 9.154
R6335 GND.n4049 GND.n4048 9.154
R6336 GND.n4048 GND.n4047 9.154
R6337 GND.n4167 GND.n4166 9.154
R6338 GND.n4170 GND.n4169 9.154
R6339 GND.n4173 GND.n4172 9.154
R6340 GND.n4176 GND.n4175 9.154
R6341 GND.n4179 GND.n4178 9.154
R6342 GND.n4182 GND.n4181 9.154
R6343 GND.n4185 GND.n4184 9.154
R6344 GND.n4188 GND.n4187 9.154
R6345 GND.n4164 GND.n4163 9.154
R6346 GND.n11726 GND.n11725 9.154
R6347 GND.n12703 GND.n12702 9.154
R6348 GND.n11723 GND.n11722 9.154
R6349 GND.n13025 GND.n13024 9.154
R6350 GND.n11920 GND.n11919 9.154
R6351 GND.n11917 GND.n11916 9.154
R6352 GND.n11914 GND.n11913 9.154
R6353 GND.n12301 GND.n12300 9.154
R6354 GND.n12304 GND.n12303 9.154
R6355 GND.n12307 GND.n12306 9.154
R6356 GND.n13022 GND.n13021 9.154
R6357 GND.n13019 GND.n13018 9.154
R6358 GND.n7790 GND.n7789 9.154
R6359 GND.n7793 GND.n7792 9.154
R6360 GND.n7796 GND.n7795 9.154
R6361 GND.n5850 GND.n5849 9.154
R6362 GND.n5853 GND.n5852 9.154
R6363 GND.n7161 GND.n7160 9.154
R6364 GND.n6333 GND.n6332 9.154
R6365 GND.n6526 GND.n6525 9.154
R6366 GND.n6529 GND.n6528 9.154
R6367 GND.n7377 GND.n7376 9.154
R6368 GND.n7428 GND.n7427 9.154
R6369 GND.n7415 GND.n7414 9.154
R6370 GND.n7402 GND.n7401 9.154
R6371 GND.n7396 GND.n7395 9.154
R6372 GND.n7381 GND.n7380 9.154
R6373 GND.n7585 GND.n7584 9.154
R6374 GND.n7591 GND.n7590 9.154
R6375 GND.n7594 GND.n7593 9.154
R6376 GND.n7617 GND.n7616 9.154
R6377 GND.n7612 GND.n7611 9.154
R6378 GND.n7609 GND.n7608 9.154
R6379 GND.n7606 GND.n7605 9.154
R6380 GND.n7603 GND.n7602 9.154
R6381 GND.n7600 GND.n7599 9.154
R6382 GND.n7597 GND.n7596 9.154
R6383 GND.n11743 GND.n11742 9.154
R6384 GND.n12122 GND.n12121 9.154
R6385 GND.n12119 GND.n12118 9.154
R6386 GND.n12113 GND.n12112 9.154
R6387 GND.n12110 GND.n12109 9.154
R6388 GND.n12107 GND.n12106 9.154
R6389 GND.n12104 GND.n12103 9.154
R6390 GND.n12101 GND.n12100 9.154
R6391 GND.n12098 GND.n12097 9.154
R6392 GND.n11728 GND.n11727 9.154
R6393 GND.n13200 GND.n13199 9.154
R6394 GND.n13203 GND.n13202 9.154
R6395 GND.n13335 GND.n13334 9.154
R6396 GND.n13332 GND.n13331 9.154
R6397 GND.n13327 GND.n13326 9.154
R6398 GND.n11122 GND.n11121 9.154
R6399 GND.n11128 GND.n11127 9.154
R6400 GND.n11143 GND.n11142 9.154
R6401 GND.n11317 GND.n11316 9.154
R6402 GND.n11314 GND.n11313 9.154
R6403 GND.n13548 GND.n13547 9.154
R6404 GND.n13551 GND.n13550 9.154
R6405 GND.n13721 GND.n13720 9.154
R6406 GND.n14015 GND.n14014 9.154
R6407 GND.n14018 GND.n14017 9.154
R6408 GND.n14021 GND.n14020 9.154
R6409 GND.n14024 GND.n14023 9.154
R6410 GND.n14012 GND.n14011 9.154
R6411 GND.n14027 GND.n14026 9.154
R6412 GND.n8386 GND.n8385 9.154
R6413 GND.n8379 GND.n8378 9.154
R6414 GND.n5826 GND.n5825 9.154
R6415 GND.n6042 GND.n6041 9.154
R6416 GND.n6049 GND.n6048 9.154
R6417 GND.n6110 GND.n6109 9.154
R6418 GND.n6119 GND.n6118 9.154
R6419 GND.n7971 GND.n7970 9.154
R6420 GND.n7966 GND.n7965 9.154
R6421 GND.n6142 GND.n6141 9.154
R6422 GND.n6137 GND.n6136 9.154
R6423 GND.n6134 GND.n6133 9.154
R6424 GND.n6131 GND.n6130 9.154
R6425 GND.n6128 GND.n6127 9.154
R6426 GND.n6125 GND.n6124 9.154
R6427 GND.n6122 GND.n6121 9.154
R6428 GND.n12484 GND.n12483 9.154
R6429 GND.n12488 GND.n12487 9.154
R6430 GND.n12493 GND.n12492 9.154
R6431 GND.n12497 GND.n12496 9.154
R6432 GND.n12500 GND.n12499 9.154
R6433 GND.n12503 GND.n12502 9.154
R6434 GND.n12506 GND.n12505 9.154
R6435 GND.n12509 GND.n12508 9.154
R6436 GND.n12512 GND.n12511 9.154
R6437 GND.n12515 GND.n12514 9.154
R6438 GND.n12843 GND.n12842 9.154
R6439 GND.n12838 GND.n12837 9.154
R6440 GND.n12834 GND.n12833 9.154
R6441 GND.n12831 GND.n12830 9.154
R6442 GND.n12526 GND.n12525 9.154
R6443 GND.n10889 GND.n10888 9.154
R6444 GND.n10900 GND.n10899 9.154
R6445 GND.n13998 GND.n13997 9.154
R6446 GND.n14003 GND.n14002 9.154
R6447 GND.n14008 GND.n14007 9.154
R6448 GND.n8405 GND.n8404 9.154
R6449 GND.n8402 GND.n8401 9.154
R6450 GND.n8399 GND.n8398 9.154
R6451 GND.n8396 GND.n8395 9.154
R6452 GND.n8393 GND.n8392 9.154
R6453 GND.n8390 GND.n8389 9.154
R6454 GND.n4756 GND.n4755 9.154
R6455 GND.n4759 GND.n4758 9.154
R6456 GND.n4768 GND.n4767 9.154
R6457 GND.n4783 GND.n4782 9.154
R6458 GND.n3499 GND.n3498 9.154
R6459 GND.n1956 GND.n1955 9.154
R6460 GND.n2971 GND.n2970 9.154
R6461 GND.n2977 GND.n2976 9.154
R6462 GND.n15879 GND.n15878 9.154
R6463 GND.n15874 GND.n15873 9.154
R6464 GND.n14081 GND.n14080 9.154
R6465 GND.n14096 GND.n14095 9.154
R6466 GND.n14102 GND.n14101 9.154
R6467 GND.n14115 GND.n14114 9.154
R6468 GND.n15538 GND.n15537 9.154
R6469 GND.n15543 GND.n15542 9.154
R6470 GND.n15281 GND.n15280 9.154
R6471 GND.n15284 GND.n15283 9.154
R6472 GND.n15293 GND.n15292 9.154
R6473 GND.n15307 GND.n15306 9.154
R6474 GND.n14378 GND.n14377 9.154
R6475 GND.n14721 GND.n14720 9.154
R6476 GND.n14730 GND.n14729 9.154
R6477 GND.n14735 GND.n14734 9.154
R6478 GND.n14416 GND.n14415 9.154
R6479 GND.n811 GND.n810 9.154
R6480 GND.n16235 GND.n16234 9.154
R6481 GND.n16244 GND.n16243 9.154
R6482 GND.n16242 GND.n16241 9.154
R6483 GND.n16239 GND.n16238 9.154
R6484 GND.n806 GND.n805 9.154
R6485 GND.n825 GND.n824 9.154
R6486 GND.n828 GND.n827 9.154
R6487 GND.n822 GND.n821 9.154
R6488 GND.n9588 GND.n9587 9.154
R6489 GND.n9937 GND.n9936 9.154
R6490 GND.n9940 GND.n9939 9.154
R6491 GND.n9943 GND.n9942 9.154
R6492 GND.n9584 GND.n9583 9.154
R6493 GND.n9582 GND.n9581 9.154
R6494 GND.n9579 GND.n9578 9.154
R6495 GND.n9947 GND.n9946 9.154
R6496 GND.n9952 GND.n9951 9.154
R6497 GND.n9956 GND.n9955 9.154
R6498 GND.n9961 GND.n9960 9.154
R6499 GND.n9243 GND.n9242 9.154
R6500 GND.n9248 GND.n9247 9.154
R6501 GND.n9261 GND.n9260 9.154
R6502 GND.n9274 GND.n9273 9.154
R6503 GND.n9280 GND.n9279 9.154
R6504 GND.n9416 GND.n9415 9.154
R6505 GND.n1184 GND.n1183 9.154
R6506 GND.n3351 GND.n3350 9.154
R6507 GND.n3354 GND.n3353 9.154
R6508 GND.n3363 GND.n3362 9.154
R6509 GND.n3378 GND.n3377 9.154
R6510 GND.n3384 GND.n3383 9.154
R6511 GND.n3397 GND.n3396 9.154
R6512 GND.n5219 GND.n5218 9.154
R6513 GND.n5224 GND.n5223 9.154
R6514 GND.n5302 GND.n5301 9.154
R6515 GND.n5305 GND.n5304 9.154
R6516 GND.n1903 GND.n1902 9.154
R6517 GND.n9234 GND.n9233 9.154
R6518 GND.n9239 GND.n9238 9.154
R6519 GND.n10329 GND.n10328 9.154
R6520 GND.n10332 GND.n10331 9.154
R6521 GND.n10338 GND.n10337 9.154
R6522 GND.n10341 GND.n10340 9.154
R6523 GND.n10344 GND.n10343 9.154
R6524 GND.n10347 GND.n10346 9.154
R6525 GND.n10350 GND.n10349 9.154
R6526 GND.n10353 GND.n10352 9.154
R6527 GND.n10356 GND.n10355 9.154
R6528 GND.n10361 GND.n10360 9.154
R6529 GND.n10365 GND.n10364 9.154
R6530 GND.n10370 GND.n10369 9.154
R6531 GND.n10374 GND.n10373 9.154
R6532 GND.n10377 GND.n10376 9.154
R6533 GND.n10380 GND.n10379 9.154
R6534 GND.n10383 GND.n10382 9.154
R6535 GND.n10386 GND.n10385 9.154
R6536 GND.n10389 GND.n10388 9.154
R6537 GND.n10392 GND.n10391 9.154
R6538 GND.n15888 GND.n15887 9.154
R6539 GND.n15883 GND.n15882 9.154
R6540 GND.n10323 GND.n10322 9.154
R6541 GND.n10320 GND.n10319 9.154
R6542 GND.n10317 GND.n10316 9.154
R6543 GND.n10314 GND.n10313 9.154
R6544 GND.n10311 GND.n10310 9.154
R6545 GND.n8874 GND.n8873 9.154
R6546 GND.n8877 GND.n8876 9.154
R6547 GND.n8884 GND.n8883 9.154
R6548 GND.n8887 GND.n8886 9.154
R6549 GND.n5819 GND.n5818 9.154
R6550 GND.n5814 GND.n5813 9.154
R6551 GND.n5811 GND.n5810 9.154
R6552 GND.n5808 GND.n5807 9.154
R6553 GND.n5805 GND.n5804 9.154
R6554 GND.n5802 GND.n5801 9.154
R6555 GND.n5799 GND.n5798 9.154
R6556 GND.n5796 GND.n5795 9.154
R6557 GND.n1909 GND.n1908 9.154
R6558 GND.n4542 GND.n4541 9.154
R6559 GND.n4546 GND.n4545 9.154
R6560 GND.n4549 GND.n4548 9.154
R6561 GND.n4552 GND.n4551 9.154
R6562 GND.n4557 GND.n4556 9.154
R6563 GND.n4561 GND.n4560 9.154
R6564 GND.n4564 GND.n4563 9.154
R6565 GND.n4567 GND.n4566 9.154
R6566 GND.n4573 GND.n4572 9.154
R6567 GND.n4576 GND.n4575 9.154
R6568 GND.n5430 GND.n5429 9.154
R6569 GND.n5436 GND.n5435 9.154
R6570 GND.n5439 GND.n5438 9.154
R6571 GND.n5447 GND.n5446 9.154
R6572 GND.n5442 GND.n5441 9.154
R6573 GND.n5293 GND.n5292 9.154
R6574 GND.n5296 GND.n5295 9.154
R6575 GND.n5299 GND.n5298 9.154
R6576 GND.n5228 GND.n5227 9.154
R6577 GND.n5233 GND.n5232 9.154
R6578 GND.n5237 GND.n5236 9.154
R6579 GND.n5240 GND.n5239 9.154
R6580 GND.n5243 GND.n5242 9.154
R6581 GND.n5246 GND.n5245 9.154
R6582 GND.n5248 GND.n5247 9.154
R6583 GND.n5426 GND.n5425 9.154
R6584 GND.n12915 GND.n12914 9.103
R6585 GND.n13188 GND.n13137 9.103
R6586 GND.n11810 GND.n11782 9.103
R6587 GND.n12472 GND.n12471 9.103
R6588 GND.n12472 GND.n12467 9.103
R6589 GND.n12915 GND.n12910 9.103
R6590 GND.n7683 GND.n7632 9.103
R6591 GND.n7955 GND.n7927 9.103
R6592 GND.n1165 GND.n1136 9.103
R6593 GND.n1228 GND.n1199 9.103
R6594 GND.n5784 GND.n5755 9.103
R6595 GND.n3946 GND.n3917 9.103
R6596 GND.n12088 GND.n12050 9.001
R6597 GND.n11810 GND.n11794 9.001
R6598 GND.n12192 GND.n12154 9.001
R6599 GND.n7955 GND.n7939 9.001
R6600 GND.n15936 GND.n15913 9.001
R6601 GND.n16224 GND.n16208 9.001
R6602 GND.n9636 GND.n9613 9.001
R6603 GND.n9924 GND.n9908 9.001
R6604 GND.n8935 GND.n8912 9.001
R6605 GND.n9223 GND.n9207 9.001
R6606 GND.n4531 GND.n4508 9.001
R6607 GND.n3664 GND.n3648 9.001
R6608 GND.n14123 GND.n14122 9
R6609 GND.n14133 GND.n14079 9
R6610 GND.n14143 GND.n14142 9
R6611 GND.n14154 GND.n14153 9
R6612 GND.n14298 GND.n14297 9
R6613 GND.n14305 GND.n14304 9
R6614 GND.n14357 GND.n14356 9
R6615 GND.n14292 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/DRAIN 9
R6616 GND.n14165 GND.n14164 9
R6617 GND.n14186 GND.n14160 9
R6618 GND.n14196 GND.n14195 9
R6619 GND.n14207 GND.n14206 9
R6620 GND.n14286 GND.n14212 9
R6621 GND.n14281 GND.n14280 9
R6622 GND.n14274 GND.n14273 9
R6623 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/DRAIN GND.n14291 9
R6624 GND.n10787 GND.n10786 9
R6625 GND.n10797 GND.n10796 9
R6626 GND.n10805 GND.n10804 9
R6627 GND.n10765 GND.n10734 9
R6628 GND.n10815 GND.n10814 9
R6629 GND.n10825 GND.n10824 9
R6630 GND.n10831 GND.n10830 9
R6631 GND.n13937 GND.n13936 9
R6632 GND.n13896 GND.n10843 9
R6633 GND.n13904 GND.n13903 9
R6634 GND.n13914 GND.n13913 9
R6635 GND.n13924 GND.n13923 9
R6636 GND.n13930 GND.n13929 9
R6637 GND.n13887 GND.n13886 9
R6638 GND.n10908 GND.n10848 9
R6639 GND.n10917 GND.n10847 9
R6640 GND.n10924 GND.n10846 9
R6641 GND.n13809 GND.n10844 9
R6642 GND.n10949 GND.n10845 9
R6643 GND.n10944 GND.n10943 9
R6644 GND.n10934 GND.n10933 9
R6645 GND.n10957 GND.n10954 9
R6646 GND.n10966 GND.n10953 9
R6647 GND.n10973 GND.n10952 9
R6648 GND.n13781 GND.n10999 9
R6649 GND.n10998 GND.n10951 9
R6650 GND.n10993 GND.n10992 9
R6651 GND.n10983 GND.n10982 9
R6652 GND.n12769 GND.n12768 9
R6653 GND.n12825 GND.n12824 9
R6654 GND.n12815 GND.n12814 9
R6655 GND.n12807 GND.n12806 9
R6656 GND.n12781 GND.n12780 9
R6657 GND.n12787 GND.n12786 9
R6658 GND.n12797 GND.n12796 9
R6659 GND.n11448 GND.n11447 9
R6660 GND.n11458 GND.n11457 9
R6661 GND.n11466 GND.n11465 9
R6662 GND.n11663 GND.n11662 9
R6663 GND.n11476 GND.n11475 9
R6664 GND.n11486 GND.n11485 9
R6665 GND.n11492 GND.n11491 9
R6666 GND.n11559 GND.n11558 9
R6667 GND.n11518 GND.n11504 9
R6668 GND.n11526 GND.n11525 9
R6669 GND.n11536 GND.n11535 9
R6670 GND.n11546 GND.n11545 9
R6671 GND.n11552 GND.n11551 9
R6672 GND.n11509 GND.n11508 9
R6673 GND.n13264 GND.n13205 9
R6674 GND.n11650 GND.n11649 9
R6675 GND.n11640 GND.n11639 9
R6676 GND.n11632 GND.n11631 9
R6677 GND.n11051 GND.n11016 9
R6678 GND.n11028 GND.n11017 9
R6679 GND.n11023 GND.n11022 9
R6680 GND.n11622 GND.n11621 9
R6681 GND.n13212 GND.n13209 9
R6682 GND.n13221 GND.n13208 9
R6683 GND.n13228 GND.n13207 9
R6684 GND.n13253 GND.n13206 9
R6685 GND.n13248 GND.n13247 9
R6686 GND.n13238 GND.n13237 9
R6687 GND.n11431 GND.n11007 9
R6688 GND.n11422 GND.n11421 9
R6689 GND.n11414 GND.n11413 9
R6690 GND.n11377 GND.n11011 9
R6691 GND.n11388 GND.n11387 9
R6692 GND.n11394 GND.n11393 9
R6693 GND.n11404 GND.n11403 9
R6694 GND.n6103 GND.n6102 9
R6695 GND.n6093 GND.n6092 9
R6696 GND.n6085 GND.n6084 9
R6697 GND.n8218 GND.n8217 9
R6698 GND.n5831 GND.n5830 9
R6699 GND.n6065 GND.n6064 9
R6700 GND.n6075 GND.n6074 9
R6701 GND.n8307 GND.n8306 9
R6702 GND.n8364 GND.n8363 9
R6703 GND.n8354 GND.n8353 9
R6704 GND.n8346 GND.n8345 9
R6705 GND.n8320 GND.n8319 9
R6706 GND.n8326 GND.n8325 9
R6707 GND.n8336 GND.n8335 9
R6708 GND.n5973 GND.n5972 9
R6709 GND.n5845 GND.n5834 9
R6710 GND.n5836 GND.n5835 9
R6711 GND.n5927 GND.n5926 9
R6712 GND.n5935 GND.n5934 9
R6713 GND.n5945 GND.n5944 9
R6714 GND.n5955 GND.n5954 9
R6715 GND.n5961 GND.n5960 9
R6716 GND.n6395 GND.n6384 9
R6717 GND.n6386 GND.n6385 9
R6718 GND.n6376 GND.n6375 9
R6719 GND.n6382 GND.n6381 9
R6720 GND.n6358 GND.n6357 9
R6721 GND.n5917 GND.n5916 9
R6722 GND.n6514 GND.n6334 9
R6723 GND.n6505 GND.n6335 9
R6724 GND.n6498 GND.n6336 9
R6725 GND.n6468 GND.n6343 9
R6726 GND.n6489 GND.n6337 9
R6727 GND.n6480 GND.n6338 9
R6728 GND.n6475 GND.n6474 9
R6729 GND.n6885 GND.n6884 9
R6730 GND.n6840 GND.n6839 9
R6731 GND.n6848 GND.n6847 9
R6732 GND.n6858 GND.n6857 9
R6733 GND.n6868 GND.n6867 9
R6734 GND.n6874 GND.n6873 9
R6735 GND.n6830 GND.n6829 9
R6736 GND.n6595 GND.n6594 9
R6737 GND.n6605 GND.n6604 9
R6738 GND.n6613 GND.n6612 9
R6739 GND.n6650 GND.n6649 9
R6740 GND.n6623 GND.n6622 9
R6741 GND.n6633 GND.n6632 9
R6742 GND.n6639 GND.n6638 9
R6743 GND.n6823 GND.n6822 9
R6744 GND.n6813 GND.n6812 9
R6745 GND.n6805 GND.n6804 9
R6746 GND.n6766 GND.n6765 9
R6747 GND.n6779 GND.n6778 9
R6748 GND.n6785 GND.n6784 9
R6749 GND.n6795 GND.n6794 9
R6750 GND.n7490 GND.n7489 9
R6751 GND.n6573 GND.n6572 9
R6752 GND.n6563 GND.n6562 9
R6753 GND.n6555 GND.n6554 9
R6754 GND.n6163 GND.n6162 9
R6755 GND.n6535 GND.n6534 9
R6756 GND.n6545 GND.n6544 9
R6757 GND.n6982 GND.n6981 9
R6758 GND.n6972 GND.n6971 9
R6759 GND.n6964 GND.n6963 9
R6760 GND.n7525 GND.n6155 9
R6761 GND.n7519 GND.n7514 9
R6762 GND.n6944 GND.n6943 9
R6763 GND.n6954 GND.n6953 9
R6764 GND.n1678 GND.n1643 9
R6765 GND.n1668 GND.n1644 9
R6766 GND.n1659 GND.n1645 9
R6767 GND.n1649 GND.n1646 9
R6768 GND.n9491 GND.n1637 9
R6769 GND.n9486 GND.n9485 9
R6770 GND.n9479 GND.n9478 9
R6771 GND.n1586 GND.n1585 9
R6772 GND.n1608 GND.n1607 9
R6773 GND.n1618 GND.n1617 9
R6774 GND.n1629 GND.n1628 9
R6775 GND.n1821 GND.n1820 9
R6776 GND.n1827 GND.n1826 9
R6777 GND.n1838 GND.n1837 9
R6778 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN GND.n1634 9
R6779 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN GND.n9496 9
R6780 GND.n9351 GND.n9350 9
R6781 GND.n9362 GND.n9361 9
R6782 GND.n9368 GND.n9367 9
R6783 GND.n9378 GND.n9377 9
R6784 GND.n9388 GND.n9387 9
R6785 GND.n9396 GND.n9395 9
R6786 GND.n9405 GND.n9292 9
R6787 GND.n1756 GND.n1755 9
R6788 GND.n1769 GND.n1768 9
R6789 GND.n1775 GND.n1774 9
R6790 GND.n1785 GND.n1784 9
R6791 GND.n1795 GND.n1794 9
R6792 GND.n1803 GND.n1802 9
R6793 GND.n1812 GND.n1642 9
R6794 GND.n8639 GND.n8580 9
R6795 GND.n8633 GND.n8586 9
R6796 GND.n8628 GND.n8627 9
R6797 GND.n8618 GND.n8617 9
R6798 GND.n8608 GND.n8607 9
R6799 GND.n8600 GND.n8587 9
R6800 GND.n8591 GND.n8588 9
R6801 GND.n5213 GND.n5212 9
R6802 GND.n2605 GND.n2604 9
R6803 GND.n2595 GND.n2594 9
R6804 GND.n2311 GND.n2297 9
R6805 GND.n2334 GND.n2330 9
R6806 GND.n5195 GND.n5194 9
R6807 GND.n5158 GND.n5157 9
R6808 GND.n5169 GND.n5168 9
R6809 GND.n5175 GND.n5174 9
R6810 GND.n5185 GND.n5184 9
R6811 GND.n5203 GND.n5202 9
R6812 GND.n2587 GND.n2586 9
R6813 GND.n2549 GND.n2548 9
R6814 GND.n2561 GND.n2560 9
R6815 GND.n2567 GND.n2566 9
R6816 GND.n2577 GND.n2576 9
R6817 GND.n2325 GND.n2324 9
R6818 GND.n2285 GND.n2276 9
R6819 GND.n2290 GND.n2275 9
R6820 GND.n2315 GND.n2314 9
R6821 GND.n2302 GND.n2298 9
R6822 GND.n3161 GND.n3160 9
R6823 GND.n2212 GND.n2211 9
R6824 GND.n2222 GND.n2221 9
R6825 GND.n2233 GND.n2232 9
R6826 GND.n2399 GND.n2398 9
R6827 GND.n2406 GND.n2405 9
R6828 GND.n2456 GND.n2455 9
R6829 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/DRAIN GND.n2238 9
R6830 GND.n2471 GND.n2462 9
R6831 GND.n2241 GND.n2240 9
R6832 GND.n2251 GND.n2250 9
R6833 GND.n2262 GND.n2261 9
R6834 GND.n3472 GND.n2267 9
R6835 GND.n3467 GND.n3466 9
R6836 GND.n3460 GND.n3459 9
R6837 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/DRAIN GND.n3477 9
R6838 GND.n1964 GND.n1963 9
R6839 GND.n1975 GND.n1974 9
R6840 GND.n1985 GND.n1984 9
R6841 GND.n1996 GND.n1995 9
R6842 GND.n2141 GND.n2140 9
R6843 GND.n2148 GND.n2147 9
R6844 GND.n2197 GND.n2196 9
R6845 GND.n2135 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/DRAIN 9
R6846 GND.n2007 GND.n2006 9
R6847 GND.n2028 GND.n2002 9
R6848 GND.n2038 GND.n2037 9
R6849 GND.n2049 GND.n2048 9
R6850 GND.n2129 GND.n2054 9
R6851 GND.n2124 GND.n2123 9
R6852 GND.n2117 GND.n2116 9
R6853 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/DRAIN GND.n2134 9
R6854 GND.n4858 GND.n4857 9
R6855 GND.n4864 GND.n4863 9
R6856 GND.n4874 GND.n4873 9
R6857 GND.n4884 GND.n4883 9
R6858 GND.n4892 GND.n4891 9
R6859 GND.n4901 GND.n1942 9
R6860 GND.n4846 GND.n4845 9
R6861 GND.n3549 GND.n3502 9
R6862 GND.n3544 GND.n3543 9
R6863 GND.n3534 GND.n3533 9
R6864 GND.n3524 GND.n3523 9
R6865 GND.n3516 GND.n3503 9
R6866 GND.n3507 GND.n3504 9
R6867 GND.n3559 GND.n3501 9
R6868 GND.n2895 GND.n2847 9
R6869 GND.n2890 GND.n2889 9
R6870 GND.n2880 GND.n2879 9
R6871 GND.n2870 GND.n2869 9
R6872 GND.n2862 GND.n2848 9
R6873 GND.n2853 GND.n2849 9
R6874 GND.n2906 GND.n2840 9
R6875 GND.n15814 GND.n10401 9
R6876 GND.n14036 GND.n14033 9
R6877 GND.n14045 GND.n14032 9
R6878 GND.n14052 GND.n14031 9
R6879 GND.n15473 GND.n14029 9
R6880 GND.n14077 GND.n14030 9
R6881 GND.n14072 GND.n14071 9
R6882 GND.n14062 GND.n14061 9
R6883 GND.n10691 GND.n10690 9
R6884 GND.n10681 GND.n10680 9
R6885 GND.n10673 GND.n10672 9
R6886 GND.n10634 GND.n10633 9
R6887 GND.n10647 GND.n10646 9
R6888 GND.n10653 GND.n10652 9
R6889 GND.n10663 GND.n10662 9
R6890 GND.n15762 GND.n10405 9
R6891 GND.n15771 GND.n10404 9
R6892 GND.n15778 GND.n10403 9
R6893 GND.n15803 GND.n10402 9
R6894 GND.n15798 GND.n15797 9
R6895 GND.n15788 GND.n15787 9
R6896 GND.n14628 GND.n14592 9
R6897 GND.n14544 GND.n14543 9
R6898 GND.n14554 GND.n14553 9
R6899 GND.n14565 GND.n14564 9
R6900 GND.n14576 GND.n14575 9
R6901 GND.n14582 GND.n14581 9
R6902 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/DRAIN GND.n14570 9
R6903 GND.n15452 GND.n15451 9
R6904 GND.n14659 GND.n14658 9
R6905 GND.n14527 GND.n14503 9
R6906 GND.n14518 GND.n14504 9
R6907 GND.n14508 GND.n14505 9
R6908 GND.n14642 GND.n14641 9
R6909 GND.n14648 GND.n14647 9
R6910 GND.n14636 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/DRAIN 9
R6911 GND.n14494 GND.n14493 9
R6912 GND.n15316 GND.n14376 9
R6913 GND.n15325 GND.n14375 9
R6914 GND.n15332 GND.n14374 9
R6915 GND.n15369 GND.n14372 9
R6916 GND.n15357 GND.n14373 9
R6917 GND.n15352 GND.n15351 9
R6918 GND.n15342 GND.n15341 9
R6919 GND.n14461 GND.n14418 9
R6920 GND.n14452 GND.n14451 9
R6921 GND.n14444 GND.n14443 9
R6922 GND.n14978 GND.n14414 9
R6923 GND.n14413 GND.n14412 9
R6924 GND.n14424 GND.n14423 9
R6925 GND.n14434 GND.n14433 9
R6926 GND.n15008 GND.n15005 9
R6927 GND.n15017 GND.n15004 9
R6928 GND.n15024 GND.n15003 9
R6929 GND.n15055 GND.n14404 9
R6930 GND.n15049 GND.n15002 9
R6931 GND.n15044 GND.n15043 9
R6932 GND.n15034 GND.n15033 9
R6933 GND.n16384 GND.n16383 9
R6934 GND.n16339 GND.n16325 9
R6935 GND.n16351 GND.n16324 9
R6936 GND.n16361 GND.n16323 9
R6937 GND.n16379 GND.n16378 9
R6938 GND.n16373 GND.n16372 9
R6939 GND.n16497 GND.n16496 9
R6940 GND.n16536 GND.n16531 9
R6941 GND.n16442 GND.n16414 9
R6942 GND.n16444 GND.n16443 9
R6943 GND.n16472 GND.n16471 9
R6944 GND.n16460 GND.n16459 9
R6945 GND.n16454 GND.n16453 9
R6946 GND.n16510 GND.n16509 9
R6947 GND.n16528 GND.n16517 9
R6948 GND.n16419 GND.n16418 9
R6949 GND.n16430 GND.n16415 9
R6950 GND.n16548 GND.n16547 9
R6951 GND.n16553 GND.n16530 9
R6952 GND.n16558 GND.n16557 9
R6953 GND.n16329 GND.n16328 9
R6954 GND.n16645 GND.n16644 9
R6955 GND.n16600 GND.n16586 9
R6956 GND.n16612 GND.n16585 9
R6957 GND.n16622 GND.n16584 9
R6958 GND.n16640 GND.n16639 9
R6959 GND.n16634 GND.n16633 9
R6960 GND.n16758 GND.n16757 9
R6961 GND.n16797 GND.n16792 9
R6962 GND.n16703 GND.n16675 9
R6963 GND.n16705 GND.n16704 9
R6964 GND.n16733 GND.n16732 9
R6965 GND.n16721 GND.n16720 9
R6966 GND.n16715 GND.n16714 9
R6967 GND.n16771 GND.n16770 9
R6968 GND.n16789 GND.n16778 9
R6969 GND.n16680 GND.n16679 9
R6970 GND.n16691 GND.n16676 9
R6971 GND.n16809 GND.n16808 9
R6972 GND.n16814 GND.n16791 9
R6973 GND.n16819 GND.n16818 9
R6974 GND.n16590 GND.n16589 9
R6975 GND.n16906 GND.n16905 9
R6976 GND.n16861 GND.n16847 9
R6977 GND.n16873 GND.n16846 9
R6978 GND.n16883 GND.n16845 9
R6979 GND.n16901 GND.n16900 9
R6980 GND.n16895 GND.n16894 9
R6981 GND.n17019 GND.n17018 9
R6982 GND.n17058 GND.n17053 9
R6983 GND.n16964 GND.n16936 9
R6984 GND.n16966 GND.n16965 9
R6985 GND.n16994 GND.n16993 9
R6986 GND.n16982 GND.n16981 9
R6987 GND.n16976 GND.n16975 9
R6988 GND.n17032 GND.n17031 9
R6989 GND.n17050 GND.n17039 9
R6990 GND.n16941 GND.n16940 9
R6991 GND.n16952 GND.n16937 9
R6992 GND.n17070 GND.n17069 9
R6993 GND.n17075 GND.n17052 9
R6994 GND.n17080 GND.n17079 9
R6995 GND.n16851 GND.n16850 9
R6996 GND.n17167 GND.n17166 9
R6997 GND.n17122 GND.n17108 9
R6998 GND.n17134 GND.n17107 9
R6999 GND.n17144 GND.n17106 9
R7000 GND.n17162 GND.n17161 9
R7001 GND.n17156 GND.n17155 9
R7002 GND.n17280 GND.n17279 9
R7003 GND.n17319 GND.n17314 9
R7004 GND.n17225 GND.n17197 9
R7005 GND.n17227 GND.n17226 9
R7006 GND.n17255 GND.n17254 9
R7007 GND.n17243 GND.n17242 9
R7008 GND.n17237 GND.n17236 9
R7009 GND.n17293 GND.n17292 9
R7010 GND.n17311 GND.n17300 9
R7011 GND.n17202 GND.n17201 9
R7012 GND.n17213 GND.n17198 9
R7013 GND.n17331 GND.n17330 9
R7014 GND.n17336 GND.n17313 9
R7015 GND.n17341 GND.n17340 9
R7016 GND.n17112 GND.n17111 9
R7017 GND.n17428 GND.n17427 9
R7018 GND.n17383 GND.n17369 9
R7019 GND.n17395 GND.n17368 9
R7020 GND.n17405 GND.n17367 9
R7021 GND.n17423 GND.n17422 9
R7022 GND.n17417 GND.n17416 9
R7023 GND.n17541 GND.n17540 9
R7024 GND.n17580 GND.n17575 9
R7025 GND.n17486 GND.n17458 9
R7026 GND.n17488 GND.n17487 9
R7027 GND.n17516 GND.n17515 9
R7028 GND.n17504 GND.n17503 9
R7029 GND.n17498 GND.n17497 9
R7030 GND.n17554 GND.n17553 9
R7031 GND.n17572 GND.n17561 9
R7032 GND.n17463 GND.n17462 9
R7033 GND.n17474 GND.n17459 9
R7034 GND.n17592 GND.n17591 9
R7035 GND.n17597 GND.n17574 9
R7036 GND.n17602 GND.n17601 9
R7037 GND.n17373 GND.n17372 9
R7038 GND.n605 GND.n604 9
R7039 GND.n595 GND.n545 9
R7040 GND.n584 GND.n583 9
R7041 GND.n718 GND.n717 9
R7042 GND.n562 GND.n547 9
R7043 GND.n572 GND.n546 9
R7044 GND.n600 GND.n544 9
R7045 GND.n740 GND.n734 9
R7046 GND.n691 GND.n690 9
R7047 GND.n671 GND.n670 9
R7048 GND.n661 GND.n660 9
R7049 GND.n666 GND.n630 9
R7050 GND.n649 GND.n631 9
R7051 GND.n752 GND.n751 9
R7052 GND.n731 GND.n730 9
R7053 GND.n685 GND.n684 9
R7054 GND.n638 GND.n632 9
R7055 GND.n764 GND.n763 9
R7056 GND.n769 GND.n733 9
R7057 GND.n774 GND.n773 9
R7058 GND.n551 GND.n550 9
R7059 GND.n347 GND.n346 9
R7060 GND.n337 GND.n287 9
R7061 GND.n326 GND.n325 9
R7062 GND.n460 GND.n459 9
R7063 GND.n304 GND.n289 9
R7064 GND.n314 GND.n288 9
R7065 GND.n342 GND.n286 9
R7066 GND.n482 GND.n476 9
R7067 GND.n433 GND.n432 9
R7068 GND.n413 GND.n412 9
R7069 GND.n403 GND.n402 9
R7070 GND.n408 GND.n372 9
R7071 GND.n391 GND.n373 9
R7072 GND.n494 GND.n493 9
R7073 GND.n473 GND.n472 9
R7074 GND.n427 GND.n426 9
R7075 GND.n380 GND.n374 9
R7076 GND.n506 GND.n505 9
R7077 GND.n511 GND.n475 9
R7078 GND.n516 GND.n515 9
R7079 GND.n293 GND.n292 9
R7080 GND.n89 GND.n88 9
R7081 GND.n79 GND.n29 9
R7082 GND.n68 GND.n67 9
R7083 GND.n202 GND.n201 9
R7084 GND.n46 GND.n31 9
R7085 GND.n56 GND.n30 9
R7086 GND.n84 GND.n28 9
R7087 GND.n224 GND.n218 9
R7088 GND.n175 GND.n174 9
R7089 GND.n155 GND.n154 9
R7090 GND.n145 GND.n144 9
R7091 GND.n150 GND.n114 9
R7092 GND.n133 GND.n115 9
R7093 GND.n236 GND.n235 9
R7094 GND.n215 GND.n214 9
R7095 GND.n169 GND.n168 9
R7096 GND.n122 GND.n116 9
R7097 GND.n248 GND.n247 9
R7098 GND.n253 GND.n217 9
R7099 GND.n258 GND.n257 9
R7100 GND.n35 GND.n34 9
R7101 GND.n17925 GND.n17924 9
R7102 GND.n17915 GND.n17865 9
R7103 GND.n17904 GND.n17903 9
R7104 GND.n17712 GND.n17711 9
R7105 GND.n17882 GND.n17867 9
R7106 GND.n17892 GND.n17866 9
R7107 GND.n17920 GND.n17864 9
R7108 GND.n17813 GND.n17807 9
R7109 GND.n17790 GND.n17789 9
R7110 GND.n17770 GND.n17769 9
R7111 GND.n17760 GND.n17759 9
R7112 GND.n17765 GND.n17729 9
R7113 GND.n17748 GND.n17730 9
R7114 GND.n17825 GND.n17824 9
R7115 GND.n17725 GND.n17724 9
R7116 GND.n17784 GND.n17783 9
R7117 GND.n17737 GND.n17731 9
R7118 GND.n17837 GND.n17836 9
R7119 GND.n17842 GND.n17806 9
R7120 GND.n17847 GND.n17846 9
R7121 GND.n17871 GND.n17870 9
R7122 GND.n11810 GND.n11774 8.901
R7123 GND.n12472 GND.n12449 8.901
R7124 GND.n12915 GND.n12892 8.901
R7125 GND.n7955 GND.n7919 8.901
R7126 GND.n16224 GND.n16204 8.901
R7127 GND.n882 GND.n876 8.901
R7128 GND.n9924 GND.n9904 8.901
R7129 GND.n1520 GND.n1514 8.901
R7130 GND.n9223 GND.n9203 8.901
R7131 GND.n4242 GND.n4236 8.901
R7132 GND.n3664 GND.n3644 8.901
R7133 GND.n5501 GND.n5495 8.901
R7134 GND.n12088 GND.n12065 8.803
R7135 GND.n11810 GND.n11802 8.803
R7136 GND.n12192 GND.n12169 8.803
R7137 GND.n7955 GND.n7947 8.803
R7138 GND.n15936 GND.n15922 8.803
R7139 GND.n16224 GND.n16216 8.803
R7140 GND.n9636 GND.n9622 8.803
R7141 GND.n9924 GND.n9916 8.803
R7142 GND.n8935 GND.n8921 8.803
R7143 GND.n9223 GND.n9215 8.803
R7144 GND.n4531 GND.n4517 8.803
R7145 GND.n3664 GND.n3656 8.803
R7146 GND.n10903 GND.n10902 8.764
R7147 GND.n13868 GND.n13867 8.764
R7148 GND.n13530 GND.n13529 8.764
R7149 GND.n11125 GND.n11124 8.764
R7150 GND.n5911 GND.n5910 8.764
R7151 GND.n6046 GND.n6045 8.764
R7152 GND.n7399 GND.n7398 8.764
R7153 GND.n7183 GND.n7182 8.764
R7154 GND.n1696 GND.n1695 8.764
R7155 GND.n9277 GND.n9276 8.764
R7156 GND.n2489 GND.n2488 8.764
R7157 GND.n3381 GND.n3380 8.764
R7158 GND.n4786 GND.n4785 8.764
R7159 GND.n4906 GND.n4905 8.764
R7160 GND.n14099 GND.n14098 8.764
R7161 GND.n15738 GND.n15737 8.764
R7162 GND.n15428 GND.n15427 8.764
R7163 GND.n15311 GND.n15310 8.764
R7164 GND.n11810 GND.n11766 8.707
R7165 GND.n12472 GND.n12432 8.707
R7166 GND.n12915 GND.n12875 8.707
R7167 GND.n7955 GND.n7911 8.707
R7168 GND.n16224 GND.n16197 8.707
R7169 GND.n882 GND.n860 8.707
R7170 GND.n9924 GND.n9897 8.707
R7171 GND.n1520 GND.n1498 8.707
R7172 GND.n9223 GND.n9196 8.707
R7173 GND.n4242 GND.n4220 8.707
R7174 GND.n3664 GND.n3637 8.707
R7175 GND.n5501 GND.n5479 8.707
R7176 GND.n4005 GND.n4002 8.704
R7177 GND.n12088 GND.n12080 8.613
R7178 GND.n11810 GND.n11809 8.613
R7179 GND.n12192 GND.n12184 8.613
R7180 GND.n7955 GND.n7954 8.613
R7181 GND.n15936 GND.n15931 8.613
R7182 GND.n16224 GND.n16223 8.613
R7183 GND.n9636 GND.n9631 8.613
R7184 GND.n9924 GND.n9923 8.613
R7185 GND.n8935 GND.n8930 8.613
R7186 GND.n9223 GND.n9222 8.613
R7187 GND.n4531 GND.n4526 8.613
R7188 GND.n3664 GND.n3663 8.613
R7189 GND.n12522 GND.n12521 8.522
R7190 GND.n13343 GND.n13342 8.522
R7191 GND.n12916 GND.n12915 8.522
R7192 GND.n11810 GND.n11759 8.522
R7193 GND.n11813 GND.n11810 8.522
R7194 GND.n12089 GND.n12088 8.522
R7195 GND.n12473 GND.n12472 8.522
R7196 GND.n12472 GND.n12417 8.522
R7197 GND.n12193 GND.n12192 8.522
R7198 GND.n12915 GND.n12860 8.522
R7199 GND.n7956 GND.n7955 8.522
R7200 GND.n7955 GND.n7904 8.522
R7201 GND.n7983 GND.n7982 8.522
R7202 GND.n7152 GND.n7151 8.522
R7203 GND.n6171 GND.n6170 8.522
R7204 GND.n16224 GND.n16190 8.522
R7205 GND.n16225 GND.n16224 8.522
R7206 GND.n883 GND.n882 8.522
R7207 GND.n882 GND.n845 8.522
R7208 GND.n9924 GND.n9890 8.522
R7209 GND.n9925 GND.n9924 8.522
R7210 GND.n1521 GND.n1520 8.522
R7211 GND.n1520 GND.n1483 8.522
R7212 GND.n9973 GND.n9970 8.522
R7213 GND.n9223 GND.n9189 8.522
R7214 GND.n9224 GND.n9223 8.522
R7215 GND.n5502 GND.n5501 8.522
R7216 GND.n4242 GND.n4205 8.522
R7217 GND.n4243 GND.n4242 8.522
R7218 GND.n15714 GND.n15713 8.522
R7219 GND.n4585 GND.n4584 8.522
R7220 GND.n4931 GND.n4930 8.522
R7221 GND.n3142 GND.n3141 8.522
R7222 GND.n3342 GND.n3341 8.522
R7223 GND.n14747 GND.n14746 8.522
R7224 GND.n15119 GND.n15116 8.522
R7225 GND.n3664 GND.n3630 8.522
R7226 GND.n3667 GND.n3664 8.522
R7227 GND.n5501 GND.n5464 8.522
R7228 GND.n12119 GND.n12116 8.282
R7229 GND.n12493 GND.n12490 8.282
R7230 GND.n10370 GND.n10367 8.282
R7231 GND.n822 GND.n819 8.282
R7232 GND.n14651 GND.n14650 7.99
R7233 GND.n14585 GND.n14584 7.99
R7234 GND.n15808 GND.n15807 7.99
R7235 GND.n10642 GND.n10641 7.99
R7236 GND.n15467 GND.n15466 7.99
R7237 GND.n14310 GND.n14309 7.99
R7238 GND.n14214 GND.n14213 7.99
R7239 GND.n2900 GND.n2899 7.99
R7240 GND.n3553 GND.n3552 7.99
R7241 GND.n4853 GND.n4852 7.99
R7242 GND.n12776 GND.n12775 7.99
R7243 GND.n10731 GND.n10730 7.99
R7244 GND.n10727 GND.n10726 7.99
R7245 GND.n13803 GND.n13802 7.99
R7246 GND.n13787 GND.n13786 7.99
R7247 GND.n11655 GND.n11654 7.99
R7248 GND.n11441 GND.n11440 7.99
R7249 GND.n11045 GND.n11044 7.99
R7250 GND.n13258 GND.n13257 7.99
R7251 GND.n11383 GND.n11382 7.99
R7252 GND.n8224 GND.n8223 7.99
R7253 GND.n8315 GND.n8314 7.99
R7254 GND.n5965 GND.n5964 7.99
R7255 GND.n6877 GND.n6876 7.99
R7256 GND.n6642 GND.n6641 7.99
R7257 GND.n6774 GND.n6773 7.99
R7258 GND.n7497 GND.n7496 7.99
R7259 GND.n6158 GND.n6157 7.99
R7260 GND.n9357 GND.n9356 7.99
R7261 GND.n1764 GND.n1763 7.99
R7262 GND.n1639 GND.n1638 7.99
R7263 GND.n1830 GND.n1829 7.99
R7264 GND.n8584 GND.n8583 7.99
R7265 GND.n2556 GND.n2555 7.99
R7266 GND.n2270 GND.n2269 7.99
R7267 GND.n2412 GND.n2411 7.99
R7268 GND.n2293 GND.n2292 7.99
R7269 GND.n5164 GND.n5163 7.99
R7270 GND.n2057 GND.n2056 7.99
R7271 GND.n2153 GND.n2152 7.99
R7272 GND.n15363 GND.n15362 7.99
R7273 GND.n14985 GND.n14984 7.99
R7274 GND.n14407 GND.n14406 7.99
R7275 GND.n6341 GND.n6340 7.99
R7276 GND.n6363 GND.n6362 7.99
R7277 GND.n4557 GND.n4554 7.905
R7278 GND.n4153 GND.n4148 7.68
R7279 GND.n2803 GND.n2800 7.68
R7280 GND.n8884 GND.n8881 7.529
R7281 GND.n9239 GND.n9236 7.529
R7282 GND.n12915 GND.n12868 7.027
R7283 GND.n12915 GND.n12884 7.027
R7284 GND.n12915 GND.n12901 7.027
R7285 GND.n12088 GND.n12033 7.027
R7286 GND.n12088 GND.n12042 7.027
R7287 GND.n12088 GND.n12058 7.027
R7288 GND.n12088 GND.n12073 7.027
R7289 GND.n12192 GND.n12137 7.027
R7290 GND.n12472 GND.n12425 7.027
R7291 GND.n12472 GND.n12441 7.027
R7292 GND.n12472 GND.n12458 7.027
R7293 GND.n12192 GND.n12146 7.027
R7294 GND.n12192 GND.n12162 7.027
R7295 GND.n12192 GND.n12177 7.027
R7296 GND.n15936 GND.n15927 7.027
R7297 GND.n15936 GND.n15918 7.027
R7298 GND.n15936 GND.n15909 7.027
R7299 GND.n15936 GND.n15904 7.027
R7300 GND.n882 GND.n881 7.027
R7301 GND.n882 GND.n869 7.027
R7302 GND.n882 GND.n853 7.027
R7303 GND.n9636 GND.n9627 7.027
R7304 GND.n9636 GND.n9618 7.027
R7305 GND.n9636 GND.n9609 7.027
R7306 GND.n9636 GND.n9604 7.027
R7307 GND.n1520 GND.n1519 7.027
R7308 GND.n1520 GND.n1507 7.027
R7309 GND.n1520 GND.n1491 7.027
R7310 GND.n8935 GND.n8926 7.027
R7311 GND.n8935 GND.n8917 7.027
R7312 GND.n8935 GND.n8908 7.027
R7313 GND.n8935 GND.n8903 7.027
R7314 GND.n5501 GND.n5500 7.027
R7315 GND.n5501 GND.n5488 7.027
R7316 GND.n5501 GND.n5472 7.027
R7317 GND.n4242 GND.n4241 7.027
R7318 GND.n4242 GND.n4229 7.027
R7319 GND.n4242 GND.n4213 7.027
R7320 GND.n4531 GND.n4522 7.027
R7321 GND.n4531 GND.n4513 7.027
R7322 GND.n4531 GND.n4504 7.027
R7323 GND.n4531 GND.n4499 7.027
R7324 GND.n4069 GND.n4065 6.912
R7325 GND.n2750 GND.n2747 6.912
R7326 GND.n14468 GND.n14467 6.885
R7327 GND.n14482 GND.n14481 6.885
R7328 GND.n15433 GND.n15432 6.885
R7329 GND.n15743 GND.n15742 6.885
R7330 GND.n15732 GND.n15731 6.885
R7331 GND.n14090 GND.n14089 6.885
R7332 GND.n14107 GND.n14106 6.885
R7333 GND.n2662 GND.n2661 6.885
R7334 GND.n4911 GND.n4910 6.885
R7335 GND.n1948 GND.n1947 6.885
R7336 GND.n4777 GND.n4776 6.885
R7337 GND.n7188 GND.n7187 6.885
R7338 GND.n7177 GND.n7176 6.885
R7339 GND.n7407 GND.n7406 6.885
R7340 GND.n7390 GND.n7389 6.885
R7341 GND.n10775 GND.n10774 6.885
R7342 GND.n13873 GND.n13872 6.885
R7343 GND.n10883 GND.n10882 6.885
R7344 GND.n10894 GND.n10893 6.885
R7345 GND.n11116 GND.n11115 6.885
R7346 GND.n11133 GND.n11132 6.885
R7347 GND.n13524 GND.n13523 6.885
R7348 GND.n13535 GND.n13534 6.885
R7349 GND.n6036 GND.n6035 6.885
R7350 GND.n8241 GND.n8240 6.885
R7351 GND.n5905 GND.n5904 6.885
R7352 GND.n9268 GND.n9267 6.885
R7353 GND.n9285 GND.n9284 6.885
R7354 GND.n1574 GND.n1573 6.885
R7355 GND.n1690 GND.n1689 6.885
R7356 GND.n3372 GND.n3371 6.885
R7357 GND.n3389 GND.n3388 6.885
R7358 GND.n3168 GND.n3167 6.885
R7359 GND.n2483 GND.n2482 6.885
R7360 GND.n4573 GND.n4570 6.776
R7361 GND.n5796 GND.n5793 6.776
R7362 GND.n5233 GND.n5230 6.776
R7363 GND.n5447 GND.n5444 6.776
R7364 GND.n3912 GND.n3911 6.716
R7365 GND.n3932 GND.n3931 6.716
R7366 GND.n7627 GND.n7626 6.716
R7367 GND.n7657 GND.n7656 6.716
R7368 GND.n13132 GND.n13131 6.716
R7369 GND.n13162 GND.n13161 6.716
R7370 GND.n13161 GND.n13160 6.716
R7371 GND.n13133 GND.n13132 6.716
R7372 GND.n12082 GND.n12081 6.716
R7373 GND.n12083 GND.n12082 6.716
R7374 GND.n12186 GND.n12185 6.716
R7375 GND.n12187 GND.n12186 6.716
R7376 GND.n7656 GND.n7655 6.716
R7377 GND.n7628 GND.n7627 6.716
R7378 GND.n7208 GND.n7207 6.716
R7379 GND.n7209 GND.n7208 6.716
R7380 GND.n11152 GND.n11151 6.716
R7381 GND.n13559 GND.n13558 6.716
R7382 GND.n11151 GND.n11150 6.716
R7383 GND.n13558 GND.n13557 6.716
R7384 GND.n10411 GND.n10410 6.716
R7385 GND.n10564 GND.n10563 6.716
R7386 GND.n8898 GND.n8897 6.716
R7387 GND.n8932 GND.n8931 6.716
R7388 GND.n9599 GND.n9598 6.716
R7389 GND.n9633 GND.n9632 6.716
R7390 GND.n15899 GND.n15898 6.716
R7391 GND.n15933 GND.n15932 6.716
R7392 GND.n15934 GND.n15933 6.716
R7393 GND.n15898 GND.n15897 6.716
R7394 GND.n1131 GND.n1130 6.716
R7395 GND.n1151 GND.n1150 6.716
R7396 GND.n1150 GND.n1149 6.716
R7397 GND.n1132 GND.n1131 6.716
R7398 GND.n9634 GND.n9633 6.716
R7399 GND.n9598 GND.n9597 6.716
R7400 GND.n1194 GND.n1193 6.716
R7401 GND.n1214 GND.n1213 6.716
R7402 GND.n1213 GND.n1212 6.716
R7403 GND.n1195 GND.n1194 6.716
R7404 GND.n10302 GND.n10301 6.716
R7405 GND.n10142 GND.n10141 6.716
R7406 GND.n10125 GND.n10124 6.716
R7407 GND.n10143 GND.n10142 6.716
R7408 GND.n10301 GND.n10300 6.716
R7409 GND.n10126 GND.n10125 6.716
R7410 GND.n8864 GND.n8863 6.716
R7411 GND.n8712 GND.n8711 6.716
R7412 GND.n8412 GND.n8411 6.716
R7413 GND.n8711 GND.n8710 6.716
R7414 GND.n8865 GND.n8864 6.716
R7415 GND.n8413 GND.n8412 6.716
R7416 GND.n8933 GND.n8932 6.716
R7417 GND.n8897 GND.n8896 6.716
R7418 GND.n5750 GND.n5749 6.716
R7419 GND.n5770 GND.n5769 6.716
R7420 GND.n5769 GND.n5768 6.716
R7421 GND.n5751 GND.n5750 6.716
R7422 GND.n4494 GND.n4493 6.716
R7423 GND.n4528 GND.n4527 6.716
R7424 GND.n4529 GND.n4528 6.716
R7425 GND.n4493 GND.n4492 6.716
R7426 GND.n10563 GND.n10562 6.716
R7427 GND.n10412 GND.n10411 6.716
R7428 GND.n3931 GND.n3930 6.716
R7429 GND.n3913 GND.n3912 6.716
R7430 GND.n4112 GND.n4105 6.656
R7431 GND.n4108 GND.n4107 6.656
R7432 GND.n2977 GND.n2973 6.4
R7433 GND.n14726 GND.n14723 6.276
R7434 GND.n15290 GND.n15287 6.276
R7435 GND.n14918 GND.n14915 6.276
R7436 GND.n15443 GND.n15440 6.276
R7437 GND.n15756 GND.n15753 6.276
R7438 GND.n15722 GND.n15719 6.276
R7439 GND.n10399 GND.n10396 6.276
R7440 GND.n15534 GND.n15531 6.276
R7441 GND.n2635 GND.n2632 6.276
R7442 GND.n1939 GND.n1936 6.276
R7443 GND.n2967 GND.n2964 6.276
R7444 GND.n4765 GND.n4762 6.276
R7445 GND.n6580 GND.n6577 6.276
R7446 GND.n7167 GND.n7164 6.276
R7447 GND.n7422 GND.n7419 6.276
R7448 GND.n6153 GND.n6150 6.276
R7449 GND.n12708 GND.n12705 6.276
R7450 GND.n11003 GND.n11000 6.276
R7451 GND.n12531 GND.n12528 6.276
R7452 GND.n10722 GND.n10719 6.276
R7453 GND.n13325 GND.n13322 6.276
R7454 GND.n11015 GND.n11012 6.276
R7455 GND.n13514 GND.n13511 6.276
R7456 GND.n11438 GND.n11435 6.276
R7457 GND.n8373 GND.n8370 6.276
R7458 GND.n6115 GND.n6112 6.276
R7459 GND.n6521 GND.n6518 6.276
R7460 GND.n8155 GND.n8152 6.276
R7461 GND.n9255 GND.n9252 6.276
R7462 GND.n9413 GND.n9410 6.276
R7463 GND.n8700 GND.n8697 6.276
R7464 GND.n1180 GND.n1177 6.276
R7465 GND.n3360 GND.n3357 6.276
R7466 GND.n1923 GND.n1920 6.276
R7467 GND.n3159 GND.n3156 6.276
R7468 GND.n1931 GND.n1928 6.276
R7469 GND.n16245 GND.n16242 6.197
R7470 GND.n9585 GND.n9582 6.197
R7471 GND.n15626 GND.n15625 6.023
R7472 GND.n15634 GND.n15633 6.023
R7473 GND.n11230 GND.n11229 6.023
R7474 GND.n11222 GND.n11221 6.023
R7475 GND.n13637 GND.n13636 6.023
R7476 GND.n13629 GND.n13628 6.023
R7477 GND.n13414 GND.n13413 6.023
R7478 GND.n13422 GND.n13421 6.023
R7479 GND.n12616 GND.n12615 6.023
R7480 GND.n12607 GND.n12606 6.023
R7481 GND.n13068 GND.n13067 6.023
R7482 GND.n13065 GND.n13064 6.023
R7483 GND.n13142 GND.n13141 6.023
R7484 GND.n12904 GND.n12903 6.023
R7485 GND.n11731 GND.n11730 6.023
R7486 GND.n12983 GND.n11733 6.023
R7487 GND.n11962 GND.n11961 6.023
R7488 GND.n11959 GND.n11958 6.023
R7489 GND.n12038 GND.n12037 6.023
R7490 GND.n11777 GND.n11776 6.023
R7491 GND.n11746 GND.n11745 6.023
R7492 GND.n11878 GND.n11748 6.023
R7493 GND.n12255 GND.n12254 6.023
R7494 GND.n12252 GND.n12251 6.023
R7495 GND.n12142 GND.n12141 6.023
R7496 GND.n12461 GND.n12460 6.023
R7497 GND.n11737 GND.n11736 6.023
R7498 GND.n12343 GND.n11739 6.023
R7499 GND.n7743 GND.n7742 6.023
R7500 GND.n7740 GND.n7739 6.023
R7501 GND.n7637 GND.n7636 6.023
R7502 GND.n7922 GND.n7921 6.023
R7503 GND.n6145 GND.n6144 6.023
R7504 GND.n7832 GND.n6147 6.023
R7505 GND.n7617 GND.n7614 6.023
R7506 GND.n7290 GND.n7289 6.023
R7507 GND.n7281 GND.n7280 6.023
R7508 GND.n6249 GND.n6248 6.023
R7509 GND.n6241 GND.n6240 6.023
R7510 GND.n6142 GND.n6139 6.023
R7511 GND.n7064 GND.n7063 6.023
R7512 GND.n7072 GND.n7071 6.023
R7513 GND.n8063 GND.n8062 6.023
R7514 GND.n8055 GND.n8054 6.023
R7515 GND.n15998 GND.n15997 6.023
R7516 GND.n15995 GND.n15994 6.023
R7517 GND.n16011 GND.n16010 6.023
R7518 GND.n16100 GND.n16099 6.023
R7519 GND.n16108 GND.n16107 6.023
R7520 GND.n1067 GND.n1066 6.023
R7521 GND.n1064 GND.n1063 6.023
R7522 GND.n1057 GND.n1056 6.023
R7523 GND.n964 GND.n963 6.023
R7524 GND.n955 GND.n954 6.023
R7525 GND.n9698 GND.n9697 6.023
R7526 GND.n9695 GND.n9694 6.023
R7527 GND.n9711 GND.n9710 6.023
R7528 GND.n9800 GND.n9799 6.023
R7529 GND.n9808 GND.n9807 6.023
R7530 GND.n1288 GND.n1287 6.023
R7531 GND.n1285 GND.n1284 6.023
R7532 GND.n1301 GND.n1300 6.023
R7533 GND.n1390 GND.n1389 6.023
R7534 GND.n1398 GND.n1397 6.023
R7535 GND.n10224 GND.n10223 6.023
R7536 GND.n10215 GND.n10214 6.023
R7537 GND.n10051 GND.n10050 6.023
R7538 GND.n10043 GND.n10042 6.023
R7539 GND.n8790 GND.n8789 6.023
R7540 GND.n8782 GND.n8781 6.023
R7541 GND.n8494 GND.n8493 6.023
R7542 GND.n8485 GND.n8484 6.023
R7543 GND.n8997 GND.n8996 6.023
R7544 GND.n8994 GND.n8993 6.023
R7545 GND.n9010 GND.n9009 6.023
R7546 GND.n9099 GND.n9098 6.023
R7547 GND.n9107 GND.n9106 6.023
R7548 GND.n5686 GND.n5685 6.023
R7549 GND.n5683 GND.n5682 6.023
R7550 GND.n5676 GND.n5675 6.023
R7551 GND.n5583 GND.n5582 6.023
R7552 GND.n5574 GND.n5573 6.023
R7553 GND.n4427 GND.n4426 6.023
R7554 GND.n4424 GND.n4423 6.023
R7555 GND.n4417 GND.n4416 6.023
R7556 GND.n4324 GND.n4323 6.023
R7557 GND.n4315 GND.n4314 6.023
R7558 GND.n4666 GND.n4665 6.023
R7559 GND.n4657 GND.n4656 6.023
R7560 GND.n5012 GND.n5011 6.023
R7561 GND.n5003 GND.n5002 6.023
R7562 GND.n3057 GND.n3056 6.023
R7563 GND.n3065 GND.n3064 6.023
R7564 GND.n3257 GND.n3256 6.023
R7565 GND.n3265 GND.n3264 6.023
R7566 GND.n10338 GND.n10335 6.023
R7567 GND.n10481 GND.n10480 6.023
R7568 GND.n10489 GND.n10488 6.023
R7569 GND.n14828 GND.n14827 6.023
R7570 GND.n14819 GND.n14818 6.023
R7571 GND.n15188 GND.n15187 6.023
R7572 GND.n15196 GND.n15195 6.023
R7573 GND.n9952 GND.n9949 6.023
R7574 GND.n3848 GND.n3847 6.023
R7575 GND.n3845 GND.n3844 6.023
R7576 GND.n3838 GND.n3837 6.023
R7577 GND.n3745 GND.n3744 6.023
R7578 GND.n3737 GND.n3736 6.023
R7579 GND.n14466 GND.n14465 5.647
R7580 GND.n15300 GND.n15299 5.647
R7581 GND.n14480 GND.n14479 5.647
R7582 GND.n15431 GND.n15430 5.647
R7583 GND.n15741 GND.n15740 5.647
R7584 GND.n15730 GND.n15729 5.647
R7585 GND.n14088 GND.n14087 5.647
R7586 GND.n14105 GND.n14104 5.647
R7587 GND.n2660 GND.n2659 5.647
R7588 GND.n4909 GND.n4908 5.647
R7589 GND.n1946 GND.n1945 5.647
R7590 GND.n4775 GND.n4774 5.647
R7591 GND.n7186 GND.n7185 5.647
R7592 GND.n7175 GND.n7174 5.647
R7593 GND.n7405 GND.n7404 5.647
R7594 GND.n7388 GND.n7387 5.647
R7595 GND.n10773 GND.n10772 5.647
R7596 GND.n13871 GND.n13870 5.647
R7597 GND.n10881 GND.n10880 5.647
R7598 GND.n10892 GND.n10891 5.647
R7599 GND.n11114 GND.n11113 5.647
R7600 GND.n11131 GND.n11130 5.647
R7601 GND.n13522 GND.n13521 5.647
R7602 GND.n13533 GND.n13532 5.647
R7603 GND.n6034 GND.n6033 5.647
R7604 GND.n6052 GND.n6051 5.647
R7605 GND.n8239 GND.n8238 5.647
R7606 GND.n5903 GND.n5902 5.647
R7607 GND.n9266 GND.n9265 5.647
R7608 GND.n9283 GND.n9282 5.647
R7609 GND.n1572 GND.n1571 5.647
R7610 GND.n1688 GND.n1687 5.647
R7611 GND.n3370 GND.n3369 5.647
R7612 GND.n3387 GND.n3386 5.647
R7613 GND.n3166 GND.n3165 5.647
R7614 GND.n2481 GND.n2480 5.647
R7615 GND.n15613 GND.n15612 5.27
R7616 GND.n15647 GND.n15646 5.27
R7617 GND.n11242 GND.n11241 5.27
R7618 GND.n11210 GND.n11209 5.27
R7619 GND.n13649 GND.n13648 5.27
R7620 GND.n13617 GND.n13616 5.27
R7621 GND.n13401 GND.n13400 5.27
R7622 GND.n13435 GND.n13434 5.27
R7623 GND.n12628 GND.n12627 5.27
R7624 GND.n12594 GND.n12593 5.27
R7625 GND.n13070 GND.n13069 5.27
R7626 GND.n13185 GND.n13184 5.27
R7627 GND.n12898 GND.n12897 5.27
R7628 GND.n12982 GND.n12981 5.27
R7629 GND.n11964 GND.n11963 5.27
R7630 GND.n12046 GND.n12045 5.27
R7631 GND.n11789 GND.n11788 5.27
R7632 GND.n11877 GND.n11876 5.27
R7633 GND.n12257 GND.n12256 5.27
R7634 GND.n12150 GND.n12149 5.27
R7635 GND.n12455 GND.n12454 5.27
R7636 GND.n12345 GND.n12344 5.27
R7637 GND.n7745 GND.n7744 5.27
R7638 GND.n7680 GND.n7679 5.27
R7639 GND.n7934 GND.n7933 5.27
R7640 GND.n7834 GND.n7833 5.27
R7641 GND.n7303 GND.n7302 5.27
R7642 GND.n7269 GND.n7268 5.27
R7643 GND.n6261 GND.n6260 5.27
R7644 GND.n6229 GND.n6228 5.27
R7645 GND.n7051 GND.n7050 5.27
R7646 GND.n7085 GND.n7084 5.27
R7647 GND.n8076 GND.n8075 5.27
R7648 GND.n8042 GND.n8041 5.27
R7649 GND.n16000 GND.n15999 5.27
R7650 GND.n16019 GND.n16018 5.27
R7651 GND.n815 GND.n814 5.27
R7652 GND.n16094 GND.n16093 5.27
R7653 GND.n16120 GND.n16119 5.27
R7654 GND.n1069 GND.n1068 5.27
R7655 GND.n1049 GND.n1048 5.27
R7656 GND.n818 GND.n817 5.27
R7657 GND.n976 GND.n975 5.27
R7658 GND.n942 GND.n941 5.27
R7659 GND.n9700 GND.n9699 5.27
R7660 GND.n9719 GND.n9718 5.27
R7661 GND.n9592 GND.n9591 5.27
R7662 GND.n9794 GND.n9793 5.27
R7663 GND.n9820 GND.n9819 5.27
R7664 GND.n1290 GND.n1289 5.27
R7665 GND.n1309 GND.n1308 5.27
R7666 GND.n1188 GND.n1187 5.27
R7667 GND.n1384 GND.n1383 5.27
R7668 GND.n1411 GND.n1410 5.27
R7669 GND.n10237 GND.n10236 5.27
R7670 GND.n10203 GND.n10202 5.27
R7671 GND.n10063 GND.n10062 5.27
R7672 GND.n10031 GND.n10030 5.27
R7673 GND.n8802 GND.n8801 5.27
R7674 GND.n8770 GND.n8769 5.27
R7675 GND.n8507 GND.n8506 5.27
R7676 GND.n8473 GND.n8472 5.27
R7677 GND.n8999 GND.n8998 5.27
R7678 GND.n9018 GND.n9017 5.27
R7679 GND.n1907 GND.n1906 5.27
R7680 GND.n9093 GND.n9092 5.27
R7681 GND.n9119 GND.n9118 5.27
R7682 GND.n5688 GND.n5687 5.27
R7683 GND.n5668 GND.n5667 5.27
R7684 GND.n1913 GND.n1912 5.27
R7685 GND.n5595 GND.n5594 5.27
R7686 GND.n5561 GND.n5560 5.27
R7687 GND.n4429 GND.n4428 5.27
R7688 GND.n4409 GND.n4408 5.27
R7689 GND.n4192 GND.n4191 5.27
R7690 GND.n4336 GND.n4335 5.27
R7691 GND.n4302 GND.n4301 5.27
R7692 GND.n4678 GND.n4677 5.27
R7693 GND.n4644 GND.n4643 5.27
R7694 GND.n5024 GND.n5023 5.27
R7695 GND.n4990 GND.n4989 5.27
R7696 GND.n3045 GND.n3044 5.27
R7697 GND.n3077 GND.n3076 5.27
R7698 GND.n3245 GND.n3244 5.27
R7699 GND.n3277 GND.n3276 5.27
R7700 GND.n15879 GND.n15876 5.27
R7701 GND.n10469 GND.n10468 5.27
R7702 GND.n10501 GND.n10500 5.27
R7703 GND.n14840 GND.n14839 5.27
R7704 GND.n14806 GND.n14805 5.27
R7705 GND.n15176 GND.n15175 5.27
R7706 GND.n15208 GND.n15207 5.27
R7707 GND.n14735 GND.n14732 5.27
R7708 GND.n3850 GND.n3849 5.27
R7709 GND.n3830 GND.n3829 5.27
R7710 GND.n3619 GND.n3618 5.27
R7711 GND.n3757 GND.n3756 5.27
R7712 GND.n3725 GND.n3724 5.27
R7713 GND.n3963 GND.n3957 5.12
R7714 GND.n2679 GND.n2675 5.12
R7715 GND.n15556 GND.n15551 4.894
R7716 GND.n15716 GND.n15710 4.894
R7717 GND.n11307 GND.n11302 4.894
R7718 GND.n11155 GND.n11149 4.894
R7719 GND.n13714 GND.n13709 4.894
R7720 GND.n13562 GND.n13556 4.894
R7721 GND.n13344 GND.n13339 4.894
R7722 GND.n13503 GND.n13498 4.894
R7723 GND.n12696 GND.n12691 4.894
R7724 GND.n12523 GND.n12518 4.894
R7725 GND.n13190 GND.n13130 4.894
R7726 GND.n13165 GND.n13164 4.894
R7727 GND.n12856 GND.n12855 4.894
R7728 GND.n12918 GND.n12851 4.894
R7729 GND.n12091 GND.n12026 4.894
R7730 GND.n12086 GND.n12085 4.894
R7731 GND.n11755 GND.n11754 4.894
R7732 GND.n11815 GND.n11752 4.894
R7733 GND.n12195 GND.n12130 4.894
R7734 GND.n12190 GND.n12189 4.894
R7735 GND.n12413 GND.n12412 4.894
R7736 GND.n12475 GND.n12408 4.894
R7737 GND.n7685 GND.n7625 4.894
R7738 GND.n7660 GND.n7659 4.894
R7739 GND.n7900 GND.n7899 4.894
R7740 GND.n7958 GND.n7895 4.894
R7741 GND.n7370 GND.n7365 4.894
R7742 GND.n7212 GND.n7206 4.894
R7743 GND.n6326 GND.n6321 4.894
R7744 GND.n6173 GND.n6167 4.894
R7745 GND.n6994 GND.n6989 4.894
R7746 GND.n7154 GND.n7148 4.894
R7747 GND.n8144 GND.n8139 4.894
R7748 GND.n7985 GND.n7979 4.894
R7749 GND.n15938 GND.n15896 4.894
R7750 GND.n16060 GND.n16059 4.894
R7751 GND.n16186 GND.n16185 4.894
R7752 GND.n16227 GND.n16181 4.894
R7753 GND.n1167 GND.n1129 4.894
R7754 GND.n1010 GND.n1009 4.894
R7755 GND.n841 GND.n840 4.894
R7756 GND.n885 GND.n836 4.894
R7757 GND.n9638 GND.n9596 4.894
R7758 GND.n9760 GND.n9759 4.894
R7759 GND.n9886 GND.n9885 4.894
R7760 GND.n9927 GND.n9881 4.894
R7761 GND.n1230 GND.n1192 4.894
R7762 GND.n1350 GND.n1349 4.894
R7763 GND.n1479 GND.n1478 4.894
R7764 GND.n1523 GND.n1474 4.894
R7765 GND.n10304 GND.n10299 4.894
R7766 GND.n10146 GND.n10140 4.894
R7767 GND.n10128 GND.n10123 4.894
R7768 GND.n9975 GND.n9969 4.894
R7769 GND.n8867 GND.n8862 4.894
R7770 GND.n8715 GND.n8709 4.894
R7771 GND.n8574 GND.n8569 4.894
R7772 GND.n8416 GND.n8410 4.894
R7773 GND.n8937 GND.n8895 4.894
R7774 GND.n9059 GND.n9058 4.894
R7775 GND.n9185 GND.n9184 4.894
R7776 GND.n9226 GND.n9180 4.894
R7777 GND.n5786 GND.n5748 4.894
R7778 GND.n5629 GND.n5628 4.894
R7779 GND.n5460 GND.n5459 4.894
R7780 GND.n5504 GND.n5455 4.894
R7781 GND.n4533 GND.n4491 4.894
R7782 GND.n4370 GND.n4369 4.894
R7783 GND.n4201 GND.n4200 4.894
R7784 GND.n4245 GND.n4196 4.894
R7785 GND.n4746 GND.n4741 4.894
R7786 GND.n4587 GND.n4581 4.894
R7787 GND.n5092 GND.n5087 4.894
R7788 GND.n4933 GND.n4927 4.894
R7789 GND.n2990 GND.n2985 4.894
R7790 GND.n3143 GND.n3138 4.894
R7791 GND.n3190 GND.n3186 4.894
R7792 GND.n3344 GND.n3338 4.894
R7793 GND.n10414 GND.n10409 4.894
R7794 GND.n10567 GND.n10561 4.894
R7795 GND.n14908 GND.n14903 4.894
R7796 GND.n14749 GND.n14743 4.894
R7797 GND.n15121 GND.n15115 4.894
R7798 GND.n15274 GND.n15269 4.894
R7799 GND.n3948 GND.n3910 4.894
R7800 GND.n3791 GND.n3790 4.894
R7801 GND.n3626 GND.n3625 4.894
R7802 GND.n3669 GND.n3623 4.894
R7803 GND.n2680 GND.n2674 4.801
R7804 GND.n3964 GND.n3956 4.801
R7805 GND.n15717 GND.n15716 4.786
R7806 GND.n13345 GND.n13344 4.786
R7807 GND.n12524 GND.n12523 4.786
R7808 GND.n15122 GND.n15121 4.786
R7809 GND.n4168 GND.n4167 4.65
R7810 GND.n4161 GND.n4160 4.65
R7811 GND.n4058 GND.n4057 4.65
R7812 GND.n4156 GND.n4155 4.65
R7813 GND.n2809 GND.n2808 4.65
R7814 GND.n2806 GND.n2805 4.65
R7815 GND.n2741 GND.n2740 4.65
R7816 GND.n2814 GND.n2813 4.65
R7817 GND.n2836 GND.n2835 4.65
R7818 GND.n2833 GND.n2832 4.65
R7819 GND.n2830 GND.n2829 4.65
R7820 GND.n2827 GND.n2826 4.65
R7821 GND.n2823 GND.n2822 4.65
R7822 GND.n2820 GND.n2819 4.65
R7823 GND.n2817 GND.n2816 4.65
R7824 GND.n2839 GND.n2838 4.65
R7825 GND.n2736 GND.n2735 4.65
R7826 GND.n2751 GND.n2750 4.65
R7827 GND.n4070 GND.n4069 4.65
R7828 GND.n4050 GND.n4049 4.65
R7829 GND.n4171 GND.n4170 4.65
R7830 GND.n4174 GND.n4173 4.65
R7831 GND.n4177 GND.n4176 4.65
R7832 GND.n4180 GND.n4179 4.65
R7833 GND.n4183 GND.n4182 4.65
R7834 GND.n4186 GND.n4185 4.65
R7835 GND.n4189 GND.n4188 4.65
R7836 GND.n4165 GND.n4164 4.65
R7837 GND.n13552 GND.n13551 4.65
R7838 GND.n14025 GND.n14024 4.65
R7839 GND.n10904 GND.n10903 4.65
R7840 GND.n13869 GND.n13868 4.65
R7841 GND.n11724 GND.n11723 4.65
R7842 GND.n12704 GND.n12703 4.65
R7843 GND.n13509 GND.n11726 4.65
R7844 GND.n13531 GND.n13530 4.65
R7845 GND.n11126 GND.n11125 4.65
R7846 GND.n11921 GND.n11920 4.65
R7847 GND.n11918 GND.n11917 4.65
R7848 GND.n11915 GND.n11914 4.65
R7849 GND.n12302 GND.n12301 4.65
R7850 GND.n12305 GND.n12304 4.65
R7851 GND.n12308 GND.n12307 4.65
R7852 GND.n13026 GND.n13025 4.65
R7853 GND.n13023 GND.n13022 4.65
R7854 GND.n13020 GND.n13019 4.65
R7855 GND.n7791 GND.n7790 4.65
R7856 GND.n7794 GND.n7793 4.65
R7857 GND.n7797 GND.n7796 4.65
R7858 GND.n6527 GND.n6526 4.65
R7859 GND.n6524 GND.n6333 4.65
R7860 GND.n5912 GND.n5911 4.65
R7861 GND.n6047 GND.n6046 4.65
R7862 GND.n8391 GND.n8390 4.65
R7863 GND.n5851 GND.n5850 4.65
R7864 GND.n8150 GND.n5853 4.65
R7865 GND.n7400 GND.n7399 4.65
R7866 GND.n7200 GND.n6529 4.65
R7867 GND.n7184 GND.n7183 4.65
R7868 GND.n7162 GND.n7161 4.65
R7869 GND.n7378 GND.n7377 4.65
R7870 GND.n7429 GND.n7428 4.65
R7871 GND.n7416 GND.n7415 4.65
R7872 GND.n7403 GND.n7402 4.65
R7873 GND.n7397 GND.n7396 4.65
R7874 GND.n7382 GND.n7381 4.65
R7875 GND.n7586 GND.n7585 4.65
R7876 GND.n7592 GND.n7591 4.65
R7877 GND.n7595 GND.n7594 4.65
R7878 GND.n7618 GND.n7617 4.65
R7879 GND.n7613 GND.n7612 4.65
R7880 GND.n7610 GND.n7609 4.65
R7881 GND.n7607 GND.n7606 4.65
R7882 GND.n7604 GND.n7603 4.65
R7883 GND.n7601 GND.n7600 4.65
R7884 GND.n7598 GND.n7597 4.65
R7885 GND.n11744 GND.n11743 4.65
R7886 GND.n12123 GND.n12122 4.65
R7887 GND.n12120 GND.n12119 4.65
R7888 GND.n12114 GND.n12113 4.65
R7889 GND.n12111 GND.n12110 4.65
R7890 GND.n12108 GND.n12107 4.65
R7891 GND.n12105 GND.n12104 4.65
R7892 GND.n12102 GND.n12101 4.65
R7893 GND.n12099 GND.n12098 4.65
R7894 GND.n11729 GND.n11728 4.65
R7895 GND.n13201 GND.n13200 4.65
R7896 GND.n13204 GND.n13203 4.65
R7897 GND.n13336 GND.n13335 4.65
R7898 GND.n13333 GND.n13332 4.65
R7899 GND.n13328 GND.n13327 4.65
R7900 GND.n11123 GND.n11122 4.65
R7901 GND.n11129 GND.n11128 4.65
R7902 GND.n11144 GND.n11143 4.65
R7903 GND.n11318 GND.n11317 4.65
R7904 GND.n11315 GND.n11314 4.65
R7905 GND.n13549 GND.n13548 4.65
R7906 GND.n13722 GND.n13721 4.65
R7907 GND.n14016 GND.n14015 4.65
R7908 GND.n14019 GND.n14018 4.65
R7909 GND.n14022 GND.n14021 4.65
R7910 GND.n14013 GND.n14012 4.65
R7911 GND.n14028 GND.n14027 4.65
R7912 GND.n8387 GND.n8386 4.65
R7913 GND.n8380 GND.n8379 4.65
R7914 GND.n5827 GND.n5826 4.65
R7915 GND.n6043 GND.n6042 4.65
R7916 GND.n6050 GND.n6049 4.65
R7917 GND.n6111 GND.n6110 4.65
R7918 GND.n6120 GND.n6119 4.65
R7919 GND.n7972 GND.n7971 4.65
R7920 GND.n7967 GND.n7966 4.65
R7921 GND.n6143 GND.n6142 4.65
R7922 GND.n6138 GND.n6137 4.65
R7923 GND.n6135 GND.n6134 4.65
R7924 GND.n6132 GND.n6131 4.65
R7925 GND.n6129 GND.n6128 4.65
R7926 GND.n6126 GND.n6125 4.65
R7927 GND.n6123 GND.n6122 4.65
R7928 GND.n12485 GND.n12484 4.65
R7929 GND.n12489 GND.n12488 4.65
R7930 GND.n12494 GND.n12493 4.65
R7931 GND.n12498 GND.n12497 4.65
R7932 GND.n12501 GND.n12500 4.65
R7933 GND.n12504 GND.n12503 4.65
R7934 GND.n12507 GND.n12506 4.65
R7935 GND.n12510 GND.n12509 4.65
R7936 GND.n12513 GND.n12512 4.65
R7937 GND.n12516 GND.n12515 4.65
R7938 GND.n12844 GND.n12843 4.65
R7939 GND.n12839 GND.n12838 4.65
R7940 GND.n12835 GND.n12834 4.65
R7941 GND.n12832 GND.n12831 4.65
R7942 GND.n12527 GND.n12526 4.65
R7943 GND.n10890 GND.n10889 4.65
R7944 GND.n10901 GND.n10900 4.65
R7945 GND.n13999 GND.n13998 4.65
R7946 GND.n14004 GND.n14003 4.65
R7947 GND.n14009 GND.n14008 4.65
R7948 GND.n8406 GND.n8405 4.65
R7949 GND.n8403 GND.n8402 4.65
R7950 GND.n8400 GND.n8399 4.65
R7951 GND.n8397 GND.n8396 4.65
R7952 GND.n8394 GND.n8393 4.65
R7953 GND.n1697 GND.n1696 4.65
R7954 GND.n9278 GND.n9277 4.65
R7955 GND.n2490 GND.n2489 4.65
R7956 GND.n3382 GND.n3381 4.65
R7957 GND.n4787 GND.n4786 4.65
R7958 GND.n4907 GND.n4906 4.65
R7959 GND.n4757 GND.n4756 4.65
R7960 GND.n4760 GND.n4759 4.65
R7961 GND.n4769 GND.n4768 4.65
R7962 GND.n4784 GND.n4783 4.65
R7963 GND.n3500 GND.n3499 4.65
R7964 GND.n1957 GND.n1956 4.65
R7965 GND.n2972 GND.n2971 4.65
R7966 GND.n2978 GND.n2977 4.65
R7967 GND.n15880 GND.n15879 4.65
R7968 GND.n15875 GND.n15874 4.65
R7969 GND.n14082 GND.n14081 4.65
R7970 GND.n14097 GND.n14096 4.65
R7971 GND.n14103 GND.n14102 4.65
R7972 GND.n14116 GND.n14115 4.65
R7973 GND.n15539 GND.n15538 4.65
R7974 GND.n15544 GND.n15543 4.65
R7975 GND.n14100 GND.n14099 4.65
R7976 GND.n15739 GND.n15738 4.65
R7977 GND.n15429 GND.n15428 4.65
R7978 GND.n15312 GND.n15311 4.65
R7979 GND.n9962 GND.n9961 4.65
R7980 GND.n15282 GND.n15281 4.65
R7981 GND.n15285 GND.n15284 4.65
R7982 GND.n15294 GND.n15293 4.65
R7983 GND.n15308 GND.n15307 4.65
R7984 GND.n14379 GND.n14378 4.65
R7985 GND.n14722 GND.n14721 4.65
R7986 GND.n14731 GND.n14730 4.65
R7987 GND.n14736 GND.n14735 4.65
R7988 GND.n14417 GND.n14416 4.65
R7989 GND.n812 GND.n811 4.65
R7990 GND.n16236 GND.n16235 4.65
R7991 GND.n807 GND.n806 4.65
R7992 GND.n826 GND.n825 4.65
R7993 GND.n829 GND.n828 4.65
R7994 GND.n823 GND.n822 4.65
R7995 GND.n9589 GND.n9588 4.65
R7996 GND.n9938 GND.n9937 4.65
R7997 GND.n9941 GND.n9940 4.65
R7998 GND.n9944 GND.n9943 4.65
R7999 GND.n9948 GND.n9947 4.65
R8000 GND.n9953 GND.n9952 4.65
R8001 GND.n9957 GND.n9956 4.65
R8002 GND.n9244 GND.n9243 4.65
R8003 GND.n9249 GND.n9248 4.65
R8004 GND.n9262 GND.n9261 4.65
R8005 GND.n9275 GND.n9274 4.65
R8006 GND.n9281 GND.n9280 4.65
R8007 GND.n9417 GND.n9416 4.65
R8008 GND.n1185 GND.n1184 4.65
R8009 GND.n3352 GND.n3351 4.65
R8010 GND.n3355 GND.n3354 4.65
R8011 GND.n3364 GND.n3363 4.65
R8012 GND.n3379 GND.n3378 4.65
R8013 GND.n3385 GND.n3384 4.65
R8014 GND.n3398 GND.n3397 4.65
R8015 GND.n5220 GND.n5219 4.65
R8016 GND.n5225 GND.n5224 4.65
R8017 GND.n5303 GND.n5302 4.65
R8018 GND.n5306 GND.n5305 4.65
R8019 GND.n1904 GND.n1903 4.65
R8020 GND.n9235 GND.n9234 4.65
R8021 GND.n9240 GND.n9239 4.65
R8022 GND.n10330 GND.n10329 4.65
R8023 GND.n10333 GND.n10332 4.65
R8024 GND.n10339 GND.n10338 4.65
R8025 GND.n10342 GND.n10341 4.65
R8026 GND.n10345 GND.n10344 4.65
R8027 GND.n10348 GND.n10347 4.65
R8028 GND.n10351 GND.n10350 4.65
R8029 GND.n10354 GND.n10353 4.65
R8030 GND.n10357 GND.n10356 4.65
R8031 GND.n10362 GND.n10361 4.65
R8032 GND.n10366 GND.n10365 4.65
R8033 GND.n10371 GND.n10370 4.65
R8034 GND.n10375 GND.n10374 4.65
R8035 GND.n10378 GND.n10377 4.65
R8036 GND.n10381 GND.n10380 4.65
R8037 GND.n10384 GND.n10383 4.65
R8038 GND.n10387 GND.n10386 4.65
R8039 GND.n10390 GND.n10389 4.65
R8040 GND.n10393 GND.n10392 4.65
R8041 GND.n15889 GND.n15888 4.65
R8042 GND.n15884 GND.n15883 4.65
R8043 GND.n10324 GND.n10323 4.65
R8044 GND.n10321 GND.n10320 4.65
R8045 GND.n10318 GND.n10317 4.65
R8046 GND.n10315 GND.n10314 4.65
R8047 GND.n10312 GND.n10311 4.65
R8048 GND.n8875 GND.n8874 4.65
R8049 GND.n8878 GND.n8877 4.65
R8050 GND.n8885 GND.n8884 4.65
R8051 GND.n8888 GND.n8887 4.65
R8052 GND.n5820 GND.n5819 4.65
R8053 GND.n5815 GND.n5814 4.65
R8054 GND.n5812 GND.n5811 4.65
R8055 GND.n5809 GND.n5808 4.65
R8056 GND.n5806 GND.n5805 4.65
R8057 GND.n5803 GND.n5802 4.65
R8058 GND.n5800 GND.n5799 4.65
R8059 GND.n5797 GND.n5796 4.65
R8060 GND.n1910 GND.n1909 4.65
R8061 GND.n4543 GND.n4542 4.65
R8062 GND.n4547 GND.n4546 4.65
R8063 GND.n4550 GND.n4549 4.65
R8064 GND.n4553 GND.n4552 4.65
R8065 GND.n4558 GND.n4557 4.65
R8066 GND.n4562 GND.n4561 4.65
R8067 GND.n4565 GND.n4564 4.65
R8068 GND.n4568 GND.n4567 4.65
R8069 GND.n4574 GND.n4573 4.65
R8070 GND.n4577 GND.n4576 4.65
R8071 GND.n5431 GND.n5430 4.65
R8072 GND.n5437 GND.n5436 4.65
R8073 GND.n5440 GND.n5439 4.65
R8074 GND.n5448 GND.n5447 4.65
R8075 GND.n5443 GND.n5442 4.65
R8076 GND.n5294 GND.n5293 4.65
R8077 GND.n5297 GND.n5296 4.65
R8078 GND.n5300 GND.n5299 4.65
R8079 GND.n5229 GND.n5228 4.65
R8080 GND.n5234 GND.n5233 4.65
R8081 GND.n5238 GND.n5237 4.65
R8082 GND.n5241 GND.n5240 4.65
R8083 GND.n5244 GND.n5243 4.65
R8084 GND.n5427 GND.n5426 4.65
R8085 GND.n14314 GND.n14312 4.574
R8086 GND.n14278 GND.n14216 4.574
R8087 GND.n10769 GND.n10733 4.574
R8088 GND.n13932 GND.n10729 4.574
R8089 GND.n13805 GND.n13804 4.574
R8090 GND.n13789 GND.n13788 4.574
R8091 GND.n12778 GND.n12777 4.574
R8092 GND.n11658 GND.n11657 4.574
R8093 GND.n11554 GND.n11443 4.574
R8094 GND.n11047 GND.n11046 4.574
R8095 GND.n13260 GND.n13259 4.574
R8096 GND.n11385 GND.n11384 4.574
R8097 GND.n8226 GND.n8225 4.574
R8098 GND.n8317 GND.n8316 4.574
R8099 GND.n5968 GND.n5967 4.574
R8100 GND.n6366 GND.n6365 4.574
R8101 GND.n6472 GND.n6342 4.574
R8102 GND.n6880 GND.n6879 4.574
R8103 GND.n6645 GND.n6644 4.574
R8104 GND.n6776 GND.n6775 4.574
R8105 GND.n7499 GND.n7498 4.574
R8106 GND.n7521 GND.n6159 4.574
R8107 GND.n9483 GND.n1641 4.574
R8108 GND.n1833 GND.n1832 4.574
R8109 GND.n9359 GND.n9358 4.574
R8110 GND.n1766 GND.n1765 4.574
R8111 GND.n8635 GND.n8585 4.574
R8112 GND.n5166 GND.n5165 4.574
R8113 GND.n2558 GND.n2557 4.574
R8114 GND.n2295 GND.n2294 4.574
R8115 GND.n2416 GND.n2414 4.574
R8116 GND.n3464 GND.n2272 4.574
R8117 GND.n2157 GND.n2155 4.574
R8118 GND.n2121 GND.n2059 4.574
R8119 GND.n4855 GND.n4854 4.574
R8120 GND.n3555 GND.n3554 4.574
R8121 GND.n2902 GND.n2901 4.574
R8122 GND.n15469 GND.n15468 4.574
R8123 GND.n10644 GND.n10643 4.574
R8124 GND.n15810 GND.n15809 4.574
R8125 GND.n14589 GND.n14587 4.574
R8126 GND.n14654 GND.n14653 4.574
R8127 GND.n15365 GND.n15364 4.574
R8128 GND.n14987 GND.n14986 4.574
R8129 GND.n15051 GND.n14408 4.574
R8130 GND.n16391 GND.n16390 4.574
R8131 GND.n16451 GND.n16450 4.574
R8132 GND.n16565 GND.n16564 4.574
R8133 GND.n16652 GND.n16651 4.574
R8134 GND.n16712 GND.n16711 4.574
R8135 GND.n16826 GND.n16825 4.574
R8136 GND.n16913 GND.n16912 4.574
R8137 GND.n16973 GND.n16972 4.574
R8138 GND.n17087 GND.n17086 4.574
R8139 GND.n17174 GND.n17173 4.574
R8140 GND.n17234 GND.n17233 4.574
R8141 GND.n17348 GND.n17347 4.574
R8142 GND.n17435 GND.n17434 4.574
R8143 GND.n17495 GND.n17494 4.574
R8144 GND.n17609 GND.n17608 4.574
R8145 GND.n612 GND.n611 4.574
R8146 GND.n678 GND.n677 4.574
R8147 GND.n781 GND.n780 4.574
R8148 GND.n354 GND.n353 4.574
R8149 GND.n420 GND.n419 4.574
R8150 GND.n523 GND.n522 4.574
R8151 GND.n96 GND.n95 4.574
R8152 GND.n162 GND.n161 4.574
R8153 GND.n265 GND.n264 4.574
R8154 GND.n17932 GND.n17931 4.574
R8155 GND.n17777 GND.n17776 4.574
R8156 GND.n17854 GND.n17853 4.574
R8157 GND.n15601 GND.n15600 4.517
R8158 GND.n15660 GND.n15659 4.517
R8159 GND.n11254 GND.n11253 4.517
R8160 GND.n11198 GND.n11197 4.517
R8161 GND.n13661 GND.n13660 4.517
R8162 GND.n13605 GND.n13604 4.517
R8163 GND.n13389 GND.n13388 4.517
R8164 GND.n13448 GND.n13447 4.517
R8165 GND.n12641 GND.n12640 4.517
R8166 GND.n12582 GND.n12581 4.517
R8167 GND.n13082 GND.n13081 4.517
R8168 GND.n13150 GND.n13149 4.517
R8169 GND.n12887 GND.n12886 4.517
R8170 GND.n12963 GND.n12962 4.517
R8171 GND.n11976 GND.n11975 4.517
R8172 GND.n12055 GND.n12054 4.517
R8173 GND.n11769 GND.n11768 4.517
R8174 GND.n11859 GND.n11858 4.517
R8175 GND.n12239 GND.n12238 4.517
R8176 GND.n12159 GND.n12158 4.517
R8177 GND.n12444 GND.n12443 4.517
R8178 GND.n12358 GND.n12357 4.517
R8179 GND.n7728 GND.n7727 4.517
R8180 GND.n7645 GND.n7644 4.517
R8181 GND.n7914 GND.n7913 4.517
R8182 GND.n7846 GND.n7845 4.517
R8183 GND.n7315 GND.n7314 4.517
R8184 GND.n7256 GND.n7255 4.517
R8185 GND.n6273 GND.n6272 4.517
R8186 GND.n6217 GND.n6216 4.517
R8187 GND.n7039 GND.n7038 4.517
R8188 GND.n7098 GND.n7097 4.517
R8189 GND.n8089 GND.n8088 4.517
R8190 GND.n8030 GND.n8029 4.517
R8191 GND.n15982 GND.n15981 4.517
R8192 GND.n16027 GND.n16026 4.517
R8193 GND.n16132 GND.n16131 4.517
R8194 GND.n1081 GND.n1080 4.517
R8195 GND.n1041 GND.n1040 4.517
R8196 GND.n930 GND.n929 4.517
R8197 GND.n9682 GND.n9681 4.517
R8198 GND.n9727 GND.n9726 4.517
R8199 GND.n9832 GND.n9831 4.517
R8200 GND.n1273 GND.n1272 4.517
R8201 GND.n1317 GND.n1316 4.517
R8202 GND.n1424 GND.n1423 4.517
R8203 GND.n10249 GND.n10248 4.517
R8204 GND.n10190 GND.n10189 4.517
R8205 GND.n10075 GND.n10074 4.517
R8206 GND.n10019 GND.n10018 4.517
R8207 GND.n8814 GND.n8813 4.517
R8208 GND.n8758 GND.n8757 4.517
R8209 GND.n8519 GND.n8518 4.517
R8210 GND.n8460 GND.n8459 4.517
R8211 GND.n8981 GND.n8980 4.517
R8212 GND.n9026 GND.n9025 4.517
R8213 GND.n9131 GND.n9130 4.517
R8214 GND.n5700 GND.n5699 4.517
R8215 GND.n5660 GND.n5659 4.517
R8216 GND.n5549 GND.n5548 4.517
R8217 GND.n4441 GND.n4440 4.517
R8218 GND.n4401 GND.n4400 4.517
R8219 GND.n4290 GND.n4289 4.517
R8220 GND.n4691 GND.n4690 4.517
R8221 GND.n4632 GND.n4631 4.517
R8222 GND.n5037 GND.n5036 4.517
R8223 GND.n4978 GND.n4977 4.517
R8224 GND.n3033 GND.n3032 4.517
R8225 GND.n3089 GND.n3088 4.517
R8226 GND.n3233 GND.n3232 4.517
R8227 GND.n3289 GND.n3288 4.517
R8228 GND.n10457 GND.n10456 4.517
R8229 GND.n10513 GND.n10512 4.517
R8230 GND.n14853 GND.n14852 4.517
R8231 GND.n14794 GND.n14793 4.517
R8232 GND.n15164 GND.n15163 4.517
R8233 GND.n15220 GND.n15219 4.517
R8234 GND.n3862 GND.n3861 4.517
R8235 GND.n3822 GND.n3821 4.517
R8236 GND.n3713 GND.n3712 4.517
R8237 GND.n6154 GND.n6153 4.142
R8238 GND.n6116 GND.n6115 4.142
R8239 GND.n9414 GND.n9413 4.142
R8240 GND.n14727 GND.n14726 4.142
R8241 GND.n15291 GND.n15290 4.142
R8242 GND.n10400 GND.n10399 4.142
R8243 GND.n15535 GND.n15534 4.142
R8244 GND.n2968 GND.n2967 4.142
R8245 GND.n4766 GND.n4765 4.142
R8246 GND.n12532 GND.n12531 4.142
R8247 GND.n14000 GND.n10722 4.142
R8248 GND.n13329 GND.n13325 4.142
R8249 GND.n11145 GND.n11015 4.142
R8250 GND.n3361 GND.n3360 4.142
R8251 GND.n1924 GND.n1923 4.142
R8252 GND.n15569 GND.n15563 4.141
R8253 GND.n15703 GND.n15697 4.141
R8254 GND.n11295 GND.n11290 4.141
R8255 GND.n11167 GND.n11162 4.141
R8256 GND.n13702 GND.n13697 4.141
R8257 GND.n13574 GND.n13569 4.141
R8258 GND.n13357 GND.n13351 4.141
R8259 GND.n13491 GND.n13485 4.141
R8260 GND.n12684 GND.n12678 4.141
R8261 GND.n12550 GND.n12544 4.141
R8262 GND.n13123 GND.n13118 4.141
R8263 GND.n13172 GND.n13171 4.141
R8264 GND.n12866 GND.n12865 4.141
R8265 GND.n12931 GND.n12925 4.141
R8266 GND.n12019 GND.n12014 4.141
R8267 GND.n12078 GND.n12077 4.141
R8268 GND.n11805 GND.n11804 4.141
R8269 GND.n11827 GND.n11822 4.141
R8270 GND.n12207 GND.n12202 4.141
R8271 GND.n12182 GND.n12181 4.141
R8272 GND.n12423 GND.n12422 4.141
R8273 GND.n12401 GND.n12395 4.141
R8274 GND.n7697 GND.n7692 4.141
R8275 GND.n7667 GND.n7666 4.141
R8276 GND.n7950 GND.n7949 4.141
R8277 GND.n7888 GND.n7883 4.141
R8278 GND.n7358 GND.n7353 4.141
R8279 GND.n7224 GND.n7219 4.141
R8280 GND.n6314 GND.n6309 4.141
R8281 GND.n6186 GND.n6180 4.141
R8282 GND.n7007 GND.n7001 4.141
R8283 GND.n7141 GND.n7135 4.141
R8284 GND.n8132 GND.n8126 4.141
R8285 GND.n7998 GND.n7992 4.141
R8286 GND.n15950 GND.n15945 4.141
R8287 GND.n16052 GND.n16051 4.141
R8288 GND.n16219 GND.n16218 4.141
R8289 GND.n16174 GND.n16168 4.141
R8290 GND.n1122 GND.n1117 4.141
R8291 GND.n1018 GND.n1017 4.141
R8292 GND.n851 GND.n850 4.141
R8293 GND.n898 GND.n892 4.141
R8294 GND.n9650 GND.n9645 4.141
R8295 GND.n9752 GND.n9751 4.141
R8296 GND.n9919 GND.n9918 4.141
R8297 GND.n9874 GND.n9868 4.141
R8298 GND.n1242 GND.n1237 4.141
R8299 GND.n1342 GND.n1341 4.141
R8300 GND.n1489 GND.n1488 4.141
R8301 GND.n1467 GND.n1461 4.141
R8302 GND.n10292 GND.n10287 4.141
R8303 GND.n10158 GND.n10153 4.141
R8304 GND.n10116 GND.n10111 4.141
R8305 GND.n9988 GND.n9982 4.141
R8306 GND.n8855 GND.n8850 4.141
R8307 GND.n8727 GND.n8722 4.141
R8308 GND.n8562 GND.n8557 4.141
R8309 GND.n8428 GND.n8423 4.141
R8310 GND.n8949 GND.n8944 4.141
R8311 GND.n9051 GND.n9050 4.141
R8312 GND.n9218 GND.n9217 4.141
R8313 GND.n9173 GND.n9167 4.141
R8314 GND.n5741 GND.n5736 4.141
R8315 GND.n5637 GND.n5636 4.141
R8316 GND.n5470 GND.n5469 4.141
R8317 GND.n5517 GND.n5511 4.141
R8318 GND.n4484 GND.n4479 4.141
R8319 GND.n4378 GND.n4377 4.141
R8320 GND.n4211 GND.n4210 4.141
R8321 GND.n4258 GND.n4252 4.141
R8322 GND.n4734 GND.n4728 4.141
R8323 GND.n4600 GND.n4594 4.141
R8324 GND.n5080 GND.n5074 4.141
R8325 GND.n4946 GND.n4940 4.141
R8326 GND.n3002 GND.n2997 4.141
R8327 GND.n3131 GND.n3125 4.141
R8328 GND.n3202 GND.n3197 4.141
R8329 GND.n3331 GND.n3325 4.141
R8330 GND.n10426 GND.n10421 4.141
R8331 GND.n10554 GND.n10549 4.141
R8332 GND.n14896 GND.n14890 4.141
R8333 GND.n14762 GND.n14756 4.141
R8334 GND.n15133 GND.n15128 4.141
R8335 GND.n15262 GND.n15257 4.141
R8336 GND.n3903 GND.n3898 4.141
R8337 GND.n3799 GND.n3798 4.141
R8338 GND.n3659 GND.n3658 4.141
R8339 GND.n3682 GND.n3676 4.141
R8340 GND.n14919 GND.n14918 4.139
R8341 GND.n15444 GND.n15443 4.139
R8342 GND.n15757 GND.n15756 4.139
R8343 GND.n15723 GND.n15722 4.139
R8344 GND.n2672 GND.n2635 4.139
R8345 GND.n4921 GND.n1939 4.139
R8346 GND.n7198 GND.n6580 4.139
R8347 GND.n7168 GND.n7167 4.139
R8348 GND.n12709 GND.n12708 4.139
R8349 GND.n11004 GND.n11003 4.139
R8350 GND.n13515 GND.n13514 4.139
R8351 GND.n13545 GND.n11438 4.139
R8352 GND.n6522 GND.n6521 4.139
R8353 GND.n8156 GND.n8155 4.139
R8354 GND.n8701 GND.n8700 4.139
R8355 GND.n1181 GND.n1180 4.139
R8356 GND.n3178 GND.n3159 4.139
R8357 GND.n1932 GND.n1931 4.139
R8358 GND.n14725 GND.n14724 4.131
R8359 GND.n15289 GND.n15288 4.131
R8360 GND.n14917 GND.n14916 4.131
R8361 GND.n15442 GND.n15441 4.131
R8362 GND.n15755 GND.n15754 4.131
R8363 GND.n15721 GND.n15720 4.131
R8364 GND.n10398 GND.n10397 4.131
R8365 GND.n15533 GND.n15532 4.131
R8366 GND.n2634 GND.n2633 4.131
R8367 GND.n1938 GND.n1937 4.131
R8368 GND.n2966 GND.n2965 4.131
R8369 GND.n4764 GND.n4763 4.131
R8370 GND.n6579 GND.n6578 4.131
R8371 GND.n7166 GND.n7165 4.131
R8372 GND.n7421 GND.n7420 4.131
R8373 GND.n6152 GND.n6151 4.131
R8374 GND.n12707 GND.n12706 4.131
R8375 GND.n11002 GND.n11001 4.131
R8376 GND.n12530 GND.n12529 4.131
R8377 GND.n10721 GND.n10720 4.131
R8378 GND.n13324 GND.n13323 4.131
R8379 GND.n11014 GND.n11013 4.131
R8380 GND.n13513 GND.n13512 4.131
R8381 GND.n11437 GND.n11436 4.131
R8382 GND.n8372 GND.n8371 4.131
R8383 GND.n6114 GND.n6113 4.131
R8384 GND.n6520 GND.n6519 4.131
R8385 GND.n8154 GND.n8153 4.131
R8386 GND.n9254 GND.n9253 4.131
R8387 GND.n9412 GND.n9411 4.131
R8388 GND.n8699 GND.n8698 4.131
R8389 GND.n1179 GND.n1178 4.131
R8390 GND.n3359 GND.n3358 4.131
R8391 GND.n1922 GND.n1921 4.131
R8392 GND.n3158 GND.n3157 4.131
R8393 GND.n1930 GND.n1929 4.131
R8394 GND.n15588 GND.n15587 3.764
R8395 GND.n15672 GND.n15671 3.764
R8396 GND.n11266 GND.n11265 3.764
R8397 GND.n11186 GND.n11185 3.764
R8398 GND.n13673 GND.n13672 3.764
R8399 GND.n13593 GND.n13592 3.764
R8400 GND.n13376 GND.n13375 3.764
R8401 GND.n13460 GND.n13459 3.764
R8402 GND.n12653 GND.n12652 3.764
R8403 GND.n12569 GND.n12568 3.764
R8404 GND.n13094 GND.n13093 3.764
R8405 GND.n13178 GND.n13177 3.764
R8406 GND.n12881 GND.n12880 3.764
R8407 GND.n12950 GND.n12949 3.764
R8408 GND.n11989 GND.n11988 3.764
R8409 GND.n12062 GND.n12061 3.764
R8410 GND.n11797 GND.n11796 3.764
R8411 GND.n11847 GND.n11846 3.764
R8412 GND.n12227 GND.n12226 3.764
R8413 GND.n12166 GND.n12165 3.764
R8414 GND.n12438 GND.n12437 3.764
R8415 GND.n12370 GND.n12369 3.764
R8416 GND.n7716 GND.n7715 3.764
R8417 GND.n7673 GND.n7672 3.764
R8418 GND.n7942 GND.n7941 3.764
R8419 GND.n7858 GND.n7857 3.764
R8420 GND.n7328 GND.n7327 3.764
R8421 GND.n7244 GND.n7243 3.764
R8422 GND.n6285 GND.n6284 3.764
R8423 GND.n6205 GND.n6204 3.764
R8424 GND.n7026 GND.n7025 3.764
R8425 GND.n7110 GND.n7109 3.764
R8426 GND.n8101 GND.n8100 3.764
R8427 GND.n8017 GND.n8016 3.764
R8428 GND.n15970 GND.n15969 3.764
R8429 GND.n16035 GND.n16034 3.764
R8430 GND.n16211 GND.n16210 3.764
R8431 GND.n16144 GND.n16143 3.764
R8432 GND.n1093 GND.n1092 3.764
R8433 GND.n1033 GND.n1032 3.764
R8434 GND.n866 GND.n865 3.764
R8435 GND.n917 GND.n916 3.764
R8436 GND.n9670 GND.n9669 3.764
R8437 GND.n9735 GND.n9734 3.764
R8438 GND.n9911 GND.n9910 3.764
R8439 GND.n9844 GND.n9843 3.764
R8440 GND.n1261 GND.n1260 3.764
R8441 GND.n1325 GND.n1324 3.764
R8442 GND.n1504 GND.n1503 3.764
R8443 GND.n1436 GND.n1435 3.764
R8444 GND.n10262 GND.n10261 3.764
R8445 GND.n10178 GND.n10177 3.764
R8446 GND.n10087 GND.n10086 3.764
R8447 GND.n10007 GND.n10006 3.764
R8448 GND.n8826 GND.n8825 3.764
R8449 GND.n8746 GND.n8745 3.764
R8450 GND.n8532 GND.n8531 3.764
R8451 GND.n8448 GND.n8447 3.764
R8452 GND.n8969 GND.n8968 3.764
R8453 GND.n9034 GND.n9033 3.764
R8454 GND.n9210 GND.n9209 3.764
R8455 GND.n9143 GND.n9142 3.764
R8456 GND.n5712 GND.n5711 3.764
R8457 GND.n5652 GND.n5651 3.764
R8458 GND.n5485 GND.n5484 3.764
R8459 GND.n5536 GND.n5535 3.764
R8460 GND.n4454 GND.n4453 3.764
R8461 GND.n4393 GND.n4392 3.764
R8462 GND.n4226 GND.n4225 3.764
R8463 GND.n4277 GND.n4276 3.764
R8464 GND.n4703 GND.n4702 3.764
R8465 GND.n4619 GND.n4618 3.764
R8466 GND.n5049 GND.n5048 3.764
R8467 GND.n4965 GND.n4964 3.764
R8468 GND.n3021 GND.n3020 3.764
R8469 GND.n3101 GND.n3100 3.764
R8470 GND.n3221 GND.n3220 3.764
R8471 GND.n3301 GND.n3300 3.764
R8472 GND.n10445 GND.n10444 3.764
R8473 GND.n10525 GND.n10524 3.764
R8474 GND.n14865 GND.n14864 3.764
R8475 GND.n14781 GND.n14780 3.764
R8476 GND.n15152 GND.n15151 3.764
R8477 GND.n15232 GND.n15231 3.764
R8478 GND.n3874 GND.n3873 3.764
R8479 GND.n3814 GND.n3813 3.764
R8480 GND.n3651 GND.n3650 3.764
R8481 GND.n3701 GND.n3700 3.764
R8482 GND.n4046 GND.n4045 3.584
R8483 GND.n4115 GND.n4112 3.584
R8484 GND.n2732 GND.n2731 3.584
R8485 GND.n5249 GND.n5246 3.487
R8486 GND.n5249 GND.n5248 3.487
R8487 GND.n3269 GND.n3268 3.396
R8488 GND.n3921 GND.n3920 3.396
R8489 GND.n3741 GND.n3740 3.396
R8490 GND.n3069 GND.n3068 3.396
R8491 GND.n7640 GND.n7635 3.396
R8492 GND.n7931 GND.n7930 3.396
R8493 GND.n13145 GND.n13140 3.396
R8494 GND.n12032 GND.n12031 3.396
R8495 GND.n12041 GND.n12036 3.396
R8496 GND.n11786 GND.n11785 3.396
R8497 GND.n12136 GND.n12135 3.396
R8498 GND.n12145 GND.n12140 3.396
R8499 GND.n7295 GND.n7293 3.396
R8500 GND.n7286 GND.n7284 3.396
R8501 GND.n6245 GND.n6244 3.396
R8502 GND.n11226 GND.n11225 3.396
R8503 GND.n13633 GND.n13632 3.396
R8504 GND.n10493 GND.n10492 3.396
R8505 GND.n8902 GND.n8901 3.396
R8506 GND.n8907 GND.n8906 3.396
R8507 GND.n9111 GND.n9110 3.396
R8508 GND.n9603 GND.n9602 3.396
R8509 GND.n9608 GND.n9607 3.396
R8510 GND.n9812 GND.n9811 3.396
R8511 GND.n15903 GND.n15902 3.396
R8512 GND.n15908 GND.n15907 3.396
R8513 GND.n16112 GND.n16111 3.396
R8514 GND.n1140 GND.n1139 3.396
R8515 GND.n1203 GND.n1202 3.396
R8516 GND.n10229 GND.n10227 3.396
R8517 GND.n10220 GND.n10218 3.396
R8518 GND.n10047 GND.n10046 3.396
R8519 GND.n8786 GND.n8785 3.396
R8520 GND.n8499 GND.n8497 3.396
R8521 GND.n8490 GND.n8488 3.396
R8522 GND.n5759 GND.n5758 3.396
R8523 GND.n4498 GND.n4497 3.396
R8524 GND.n4503 GND.n4502 3.396
R8525 GND.n15200 GND.n15199 3.396
R8526 GND.n14408 GND.n14405 3.388
R8527 GND.n14986 GND.n14982 3.388
R8528 GND.n14653 GND.n14652 3.388
R8529 GND.n14587 GND.n14586 3.388
R8530 GND.n15809 GND.n15805 3.388
R8531 GND.n10643 GND.n10638 3.388
R8532 GND.n15468 GND.n15465 3.388
R8533 GND.n14216 GND.n14215 3.388
R8534 GND.n14312 GND.n14311 3.388
R8535 GND.n2901 GND.n2897 3.388
R8536 GND.n3554 GND.n3551 3.388
R8537 GND.n4854 GND.n4850 3.388
R8538 GND.n5165 GND.n5162 3.388
R8539 GND.n15581 GND.n15576 3.388
R8540 GND.n15690 GND.n15685 3.388
R8541 GND.n6159 GND.n6156 3.388
R8542 GND.n12777 GND.n12773 3.388
R8543 GND.n10729 GND.n10728 3.388
R8544 GND.n10733 GND.n10732 3.388
R8545 GND.n13788 GND.n13785 3.388
R8546 GND.n13804 GND.n13800 3.388
R8547 GND.n11283 GND.n11278 3.388
R8548 GND.n11179 GND.n11174 3.388
R8549 GND.n13690 GND.n13685 3.388
R8550 GND.n13586 GND.n13581 3.388
R8551 GND.n13369 GND.n13364 3.388
R8552 GND.n13478 GND.n13473 3.388
R8553 GND.n12671 GND.n12666 3.388
R8554 GND.n12562 GND.n12557 3.388
R8555 GND.n11443 GND.n11442 3.388
R8556 GND.n11657 GND.n11656 3.388
R8557 GND.n11384 GND.n11381 3.388
R8558 GND.n11046 GND.n11042 3.388
R8559 GND.n13259 GND.n13255 3.388
R8560 GND.n13111 GND.n13106 3.388
R8561 GND.n13158 GND.n13157 3.388
R8562 GND.n12871 GND.n12870 3.388
R8563 GND.n12943 GND.n12938 3.388
R8564 GND.n12007 GND.n12001 3.388
R8565 GND.n12071 GND.n12070 3.388
R8566 GND.n11762 GND.n11761 3.388
R8567 GND.n11840 GND.n11834 3.388
R8568 GND.n12220 GND.n12214 3.388
R8569 GND.n12175 GND.n12174 3.388
R8570 GND.n12428 GND.n12427 3.388
R8571 GND.n12388 GND.n12383 3.388
R8572 GND.n7709 GND.n7704 3.388
R8573 GND.n7653 GND.n7652 3.388
R8574 GND.n7907 GND.n7906 3.388
R8575 GND.n7876 GND.n7870 3.388
R8576 GND.n7346 GND.n7340 3.388
R8577 GND.n7237 GND.n7231 3.388
R8578 GND.n6302 GND.n6297 3.388
R8579 GND.n6198 GND.n6193 3.388
R8580 GND.n8225 GND.n8222 3.388
R8581 GND.n8316 GND.n8311 3.388
R8582 GND.n6342 GND.n6339 3.388
R8583 GND.n6365 GND.n6364 3.388
R8584 GND.n5967 GND.n5966 3.388
R8585 GND.n7019 GND.n7014 3.388
R8586 GND.n7128 GND.n7123 3.388
R8587 GND.n8119 GND.n8114 3.388
R8588 GND.n8010 GND.n8005 3.388
R8589 GND.n6644 GND.n6643 3.388
R8590 GND.n6879 GND.n6878 3.388
R8591 GND.n6775 GND.n6770 3.388
R8592 GND.n7498 GND.n7494 3.388
R8593 GND.n15963 GND.n15957 3.388
R8594 GND.n16044 GND.n16043 3.388
R8595 GND.n16193 GND.n16192 3.388
R8596 GND.n16161 GND.n16156 3.388
R8597 GND.n1110 GND.n1105 3.388
R8598 GND.n1026 GND.n1025 3.388
R8599 GND.n856 GND.n855 3.388
R8600 GND.n910 GND.n905 3.388
R8601 GND.n9663 GND.n9657 3.388
R8602 GND.n9744 GND.n9743 3.388
R8603 GND.n9893 GND.n9892 3.388
R8604 GND.n9861 GND.n9856 3.388
R8605 GND.n1254 GND.n1249 3.388
R8606 GND.n1334 GND.n1333 3.388
R8607 GND.n1494 GND.n1493 3.388
R8608 GND.n1454 GND.n1449 3.388
R8609 GND.n10280 GND.n10274 3.388
R8610 GND.n10171 GND.n10165 3.388
R8611 GND.n10104 GND.n10099 3.388
R8612 GND.n10000 GND.n9995 3.388
R8613 GND.n8843 GND.n8838 3.388
R8614 GND.n8739 GND.n8734 3.388
R8615 GND.n8550 GND.n8544 3.388
R8616 GND.n8441 GND.n8435 3.388
R8617 GND.n8585 GND.n8581 3.388
R8618 GND.n9358 GND.n9355 3.388
R8619 GND.n1765 GND.n1760 3.388
R8620 GND.n1641 GND.n1640 3.388
R8621 GND.n1832 GND.n1831 3.388
R8622 GND.n8962 GND.n8956 3.388
R8623 GND.n9043 GND.n9042 3.388
R8624 GND.n9192 GND.n9191 3.388
R8625 GND.n9160 GND.n9155 3.388
R8626 GND.n5729 GND.n5724 3.388
R8627 GND.n5645 GND.n5644 3.388
R8628 GND.n5475 GND.n5474 3.388
R8629 GND.n5529 GND.n5524 3.388
R8630 GND.n4472 GND.n4466 3.388
R8631 GND.n4386 GND.n4385 3.388
R8632 GND.n4216 GND.n4215 3.388
R8633 GND.n4270 GND.n4265 3.388
R8634 GND.n4721 GND.n4716 3.388
R8635 GND.n4612 GND.n4607 3.388
R8636 GND.n5067 GND.n5062 3.388
R8637 GND.n4958 GND.n4953 3.388
R8638 GND.n2557 GND.n2553 3.388
R8639 GND.n2272 GND.n2271 3.388
R8640 GND.n2414 GND.n2413 3.388
R8641 GND.n2294 GND.n2291 3.388
R8642 GND.n2059 GND.n2058 3.388
R8643 GND.n2155 GND.n2154 3.388
R8644 GND.n3014 GND.n3009 3.388
R8645 GND.n3118 GND.n3113 3.388
R8646 GND.n3214 GND.n3209 3.388
R8647 GND.n3318 GND.n3313 3.388
R8648 GND.n10438 GND.n10433 3.388
R8649 GND.n10542 GND.n10537 3.388
R8650 GND.n14883 GND.n14878 3.388
R8651 GND.n14774 GND.n14769 3.388
R8652 GND.n15364 GND.n15359 3.388
R8653 GND.n15145 GND.n15140 3.388
R8654 GND.n15250 GND.n15244 3.388
R8655 GND.n3891 GND.n3886 3.388
R8656 GND.n3807 GND.n3806 3.388
R8657 GND.n3633 GND.n3632 3.388
R8658 GND.n3694 GND.n3689 3.388
R8659 GND.n16450 GND.n16448 3.388
R8660 GND.n16564 GND.n16562 3.388
R8661 GND.n16390 GND.n16388 3.388
R8662 GND.n16711 GND.n16709 3.388
R8663 GND.n16825 GND.n16823 3.388
R8664 GND.n16651 GND.n16649 3.388
R8665 GND.n16972 GND.n16970 3.388
R8666 GND.n17086 GND.n17084 3.388
R8667 GND.n16912 GND.n16910 3.388
R8668 GND.n17233 GND.n17231 3.388
R8669 GND.n17347 GND.n17345 3.388
R8670 GND.n17173 GND.n17171 3.388
R8671 GND.n17494 GND.n17492 3.388
R8672 GND.n17608 GND.n17606 3.388
R8673 GND.n17434 GND.n17432 3.388
R8674 GND.n677 GND.n675 3.388
R8675 GND.n780 GND.n778 3.388
R8676 GND.n611 GND.n609 3.388
R8677 GND.n419 GND.n417 3.388
R8678 GND.n522 GND.n520 3.388
R8679 GND.n353 GND.n351 3.388
R8680 GND.n161 GND.n159 3.388
R8681 GND.n264 GND.n262 3.388
R8682 GND.n95 GND.n93 3.388
R8683 GND.n17776 GND.n17774 3.388
R8684 GND.n17853 GND.n17851 3.388
R8685 GND.n17931 GND.n17929 3.388
R8686 GND.n4069 GND.n4062 3.328
R8687 GND.n2750 GND.n2745 3.328
R8688 GND.n14406 GND.t192 3.326
R8689 GND.n14984 GND.n14983 3.326
R8690 GND.n14584 GND.t191 3.326
R8691 GND.n15807 GND.n15806 3.326
R8692 GND.n10641 GND.n10639 3.326
R8693 GND.n10641 GND.n10640 3.326
R8694 GND.n15466 GND.t174 3.326
R8695 GND.n14309 GND.t173 3.326
R8696 GND.n2899 GND.n2898 3.326
R8697 GND.n3552 GND.t178 3.326
R8698 GND.n4852 GND.n4851 3.326
R8699 GND.n5163 GND.t206 3.326
R8700 GND.n6157 GND.t160 3.326
R8701 GND.n12775 GND.n12774 3.326
R8702 GND.n10726 GND.n10725 3.326
R8703 GND.n10726 GND.t71 3.326
R8704 GND.n13786 GND.t72 3.326
R8705 GND.n13802 GND.n13801 3.326
R8706 GND.n11440 GND.n11439 3.326
R8707 GND.n11440 GND.t228 3.326
R8708 GND.n11382 GND.t229 3.326
R8709 GND.n11044 GND.n11043 3.326
R8710 GND.n13257 GND.n13256 3.326
R8711 GND.n8223 GND.t115 3.326
R8712 GND.n8314 GND.n8312 3.326
R8713 GND.n8314 GND.n8313 3.326
R8714 GND.n6362 GND.t116 3.326
R8715 GND.n5964 GND.n5963 3.326
R8716 GND.n6876 GND.t159 3.326
R8717 GND.n6773 GND.n6771 3.326
R8718 GND.n6773 GND.n6772 3.326
R8719 GND.n7496 GND.n7495 3.326
R8720 GND.n8583 GND.n8582 3.326
R8721 GND.n9356 GND.t210 3.326
R8722 GND.n1763 GND.n1761 3.326
R8723 GND.n1763 GND.n1762 3.326
R8724 GND.n1638 GND.t209 3.326
R8725 GND.n2555 GND.n2554 3.326
R8726 GND.n2269 GND.n2268 3.326
R8727 GND.n2269 GND.t205 3.326
R8728 GND.n2411 GND.n2410 3.326
R8729 GND.n2056 GND.n2055 3.326
R8730 GND.n2056 GND.t177 3.326
R8731 GND.n15362 GND.n15360 3.326
R8732 GND.n15362 GND.n15361 3.326
R8733 GND.n16407 GND.t39 3.326
R8734 GND.n16554 GND.t238 3.326
R8735 GND.n16554 GND.t23 3.326
R8736 GND.n16380 GND.t21 3.326
R8737 GND.n16668 GND.t15 3.326
R8738 GND.n16815 GND.t242 3.326
R8739 GND.n16815 GND.t1 3.326
R8740 GND.n16641 GND.t17 3.326
R8741 GND.n16929 GND.t43 3.326
R8742 GND.n17076 GND.t253 3.326
R8743 GND.n17076 GND.t255 3.326
R8744 GND.n16902 GND.t258 3.326
R8745 GND.n17190 GND.t41 3.326
R8746 GND.n17337 GND.t55 3.326
R8747 GND.n17337 GND.t5 3.326
R8748 GND.n17163 GND.t27 3.326
R8749 GND.n17451 GND.t19 3.326
R8750 GND.n17598 GND.t236 3.326
R8751 GND.n17598 GND.t234 3.326
R8752 GND.n17424 GND.t37 3.326
R8753 GND.n667 GND.t45 3.326
R8754 GND.n770 GND.t240 3.326
R8755 GND.n770 GND.t13 3.326
R8756 GND.n601 GND.t51 3.326
R8757 GND.n409 GND.t25 3.326
R8758 GND.n512 GND.t246 3.326
R8759 GND.n512 GND.t49 3.326
R8760 GND.n343 GND.t47 3.326
R8761 GND.n151 GND.t33 3.326
R8762 GND.n254 GND.t244 3.326
R8763 GND.n254 GND.t3 3.326
R8764 GND.n85 GND.t35 3.326
R8765 GND.n17766 GND.t29 3.326
R8766 GND.n17843 GND.t250 3.326
R8767 GND.n17843 GND.t248 3.326
R8768 GND.n17921 GND.t31 3.326
R8769 GND.n3260 GND.n3259 3.324
R8770 GND.n3917 GND.n3916 3.324
R8771 GND.n3748 GND.n3747 3.324
R8772 GND.n3060 GND.n3059 3.324
R8773 GND.n7076 GND.n7075 3.324
R8774 GND.n8058 GND.n8057 3.324
R8775 GND.n7632 GND.n7631 3.324
R8776 GND.n7927 GND.n7926 3.324
R8777 GND.n13426 GND.n13425 3.324
R8778 GND.n12611 GND.n12610 3.324
R8779 GND.n12619 GND.n12618 3.324
R8780 GND.n13417 GND.n13416 3.324
R8781 GND.n13137 GND.n13136 3.324
R8782 GND.n12914 GND.n12912 3.324
R8783 GND.n12910 GND.n12909 3.324
R8784 GND.n11782 GND.n11781 3.324
R8785 GND.n12471 GND.n12469 3.324
R8786 GND.n12467 GND.n12466 3.324
R8787 GND.n7067 GND.n7066 3.324
R8788 GND.n8067 GND.n8066 3.324
R8789 GND.n6252 GND.n6251 3.324
R8790 GND.n11233 GND.n11232 3.324
R8791 GND.n13640 GND.n13639 3.324
R8792 GND.n10484 GND.n10483 3.324
R8793 GND.n14823 GND.n14822 3.324
R8794 GND.n9102 GND.n9101 3.324
R8795 GND.n9803 GND.n9802 3.324
R8796 GND.n16103 GND.n16102 3.324
R8797 GND.n1136 GND.n1135 3.324
R8798 GND.n959 GND.n958 3.324
R8799 GND.n967 GND.n966 3.324
R8800 GND.n1199 GND.n1198 3.324
R8801 GND.n1402 GND.n1401 3.324
R8802 GND.n1393 GND.n1392 3.324
R8803 GND.n10054 GND.n10053 3.324
R8804 GND.n8793 GND.n8792 3.324
R8805 GND.n5755 GND.n5754 3.324
R8806 GND.n5578 GND.n5577 3.324
R8807 GND.n5586 GND.n5585 3.324
R8808 GND.n4319 GND.n4318 3.324
R8809 GND.n4327 GND.n4326 3.324
R8810 GND.n15638 GND.n15637 3.324
R8811 GND.n15191 GND.n15190 3.324
R8812 GND.n15629 GND.n15628 3.324
R8813 GND.n4661 GND.n4660 3.324
R8814 GND.n5007 GND.n5006 3.324
R8815 GND.n4669 GND.n4668 3.324
R8816 GND.n5015 GND.n5014 3.324
R8817 GND.n14831 GND.n14830 3.324
R8818 GND.n2680 GND.n2679 3.1
R8819 GND.n2685 GND.n2684 3.1
R8820 GND.n2690 GND.n2689 3.1
R8821 GND.n2695 GND.n2694 3.1
R8822 GND.n2700 GND.n2699 3.1
R8823 GND.n2705 GND.n2704 3.1
R8824 GND.n2708 GND.n2707 3.1
R8825 GND.n2713 GND.n2712 3.1
R8826 GND.n2718 GND.n2717 3.1
R8827 GND.n2723 GND.n2722 3.1
R8828 GND.n2730 GND.n2729 3.1
R8829 GND.n2754 GND.n2753 3.1
R8830 GND.n2759 GND.n2758 3.1
R8831 GND.n2764 GND.n2763 3.1
R8832 GND.n2769 GND.n2768 3.1
R8833 GND.n2774 GND.n2773 3.1
R8834 GND.n2777 GND.n2776 3.1
R8835 GND.n2782 GND.n2781 3.1
R8836 GND.n2787 GND.n2786 3.1
R8837 GND.n2792 GND.n2791 3.1
R8838 GND.n2797 GND.n2796 3.1
R8839 GND.n2804 GND.n2803 3.1
R8840 GND.n3964 GND.n3963 3.1
R8841 GND.n3971 GND.n3970 3.1
R8842 GND.n3978 GND.n3977 3.1
R8843 GND.n3985 GND.n3984 3.1
R8844 GND.n3992 GND.n3991 3.1
R8845 GND.n4006 GND.n4005 3.1
R8846 GND.n4013 GND.n4012 3.1
R8847 GND.n4020 GND.n4019 3.1
R8848 GND.n4027 GND.n4026 3.1
R8849 GND.n4034 GND.n4033 3.1
R8850 GND.n4044 GND.n4043 3.1
R8851 GND.n4074 GND.n4073 3.1
R8852 GND.n4081 GND.n4080 3.1
R8853 GND.n4088 GND.n4087 3.1
R8854 GND.n4095 GND.n4094 3.1
R8855 GND.n4102 GND.n4101 3.1
R8856 GND.n4116 GND.n4115 3.1
R8857 GND.n4123 GND.n4122 3.1
R8858 GND.n4130 GND.n4129 3.1
R8859 GND.n4137 GND.n4136 3.1
R8860 GND.n4144 GND.n4143 3.1
R8861 GND.n4154 GND.n4153 3.1
R8862 GND.n16240 GND.n16239 3.099
R8863 GND.n9580 GND.n9579 3.099
R8864 GND.n9585 GND.n9584 3.099
R8865 GND.n16245 GND.n16244 3.099
R8866 GND.n15576 GND.n15575 3.011
R8867 GND.n15685 GND.n15684 3.011
R8868 GND.n11278 GND.n11277 3.011
R8869 GND.n11174 GND.n11173 3.011
R8870 GND.n13685 GND.n13684 3.011
R8871 GND.n13581 GND.n13580 3.011
R8872 GND.n13364 GND.n13363 3.011
R8873 GND.n13473 GND.n13472 3.011
R8874 GND.n12666 GND.n12665 3.011
R8875 GND.n12557 GND.n12556 3.011
R8876 GND.n13106 GND.n13105 3.011
R8877 GND.n13157 GND.n13156 3.011
R8878 GND.n12870 GND.n12869 3.011
R8879 GND.n12938 GND.n12937 3.011
R8880 GND.n12001 GND.n12000 3.011
R8881 GND.n12070 GND.n12069 3.011
R8882 GND.n11761 GND.n11760 3.011
R8883 GND.n11834 GND.n11833 3.011
R8884 GND.n12214 GND.n12213 3.011
R8885 GND.n12174 GND.n12173 3.011
R8886 GND.n12427 GND.n12426 3.011
R8887 GND.n12383 GND.n12382 3.011
R8888 GND.n7704 GND.n7703 3.011
R8889 GND.n7652 GND.n7651 3.011
R8890 GND.n7906 GND.n7905 3.011
R8891 GND.n7870 GND.n7869 3.011
R8892 GND.n7340 GND.n7339 3.011
R8893 GND.n7231 GND.n7230 3.011
R8894 GND.n6297 GND.n6296 3.011
R8895 GND.n6193 GND.n6192 3.011
R8896 GND.n7014 GND.n7013 3.011
R8897 GND.n7123 GND.n7122 3.011
R8898 GND.n8114 GND.n8113 3.011
R8899 GND.n8005 GND.n8004 3.011
R8900 GND.n15957 GND.n15956 3.011
R8901 GND.n16043 GND.n16042 3.011
R8902 GND.n16192 GND.n16191 3.011
R8903 GND.n16156 GND.n16155 3.011
R8904 GND.n1105 GND.n1104 3.011
R8905 GND.n1025 GND.n1024 3.011
R8906 GND.n855 GND.n854 3.011
R8907 GND.n905 GND.n904 3.011
R8908 GND.n9657 GND.n9656 3.011
R8909 GND.n9743 GND.n9742 3.011
R8910 GND.n9892 GND.n9891 3.011
R8911 GND.n9856 GND.n9855 3.011
R8912 GND.n1249 GND.n1248 3.011
R8913 GND.n1333 GND.n1332 3.011
R8914 GND.n1493 GND.n1492 3.011
R8915 GND.n1449 GND.n1448 3.011
R8916 GND.n10274 GND.n10273 3.011
R8917 GND.n10165 GND.n10164 3.011
R8918 GND.n10099 GND.n10098 3.011
R8919 GND.n9995 GND.n9994 3.011
R8920 GND.n8838 GND.n8837 3.011
R8921 GND.n8734 GND.n8733 3.011
R8922 GND.n8544 GND.n8543 3.011
R8923 GND.n8435 GND.n8434 3.011
R8924 GND.n8956 GND.n8955 3.011
R8925 GND.n9042 GND.n9041 3.011
R8926 GND.n9191 GND.n9190 3.011
R8927 GND.n9155 GND.n9154 3.011
R8928 GND.n5724 GND.n5723 3.011
R8929 GND.n5644 GND.n5643 3.011
R8930 GND.n5474 GND.n5473 3.011
R8931 GND.n5524 GND.n5523 3.011
R8932 GND.n4466 GND.n4465 3.011
R8933 GND.n4385 GND.n4384 3.011
R8934 GND.n4215 GND.n4214 3.011
R8935 GND.n4265 GND.n4264 3.011
R8936 GND.n4716 GND.n4715 3.011
R8937 GND.n4607 GND.n4606 3.011
R8938 GND.n5062 GND.n5061 3.011
R8939 GND.n4953 GND.n4952 3.011
R8940 GND.n3009 GND.n3008 3.011
R8941 GND.n3113 GND.n3112 3.011
R8942 GND.n3209 GND.n3208 3.011
R8943 GND.n3313 GND.n3312 3.011
R8944 GND.n4542 GND.n4539 3.011
R8945 GND.n10433 GND.n10432 3.011
R8946 GND.n10537 GND.n10536 3.011
R8947 GND.n14878 GND.n14877 3.011
R8948 GND.n14769 GND.n14768 3.011
R8949 GND.n15140 GND.n15139 3.011
R8950 GND.n15244 GND.n15243 3.011
R8951 GND.n5436 GND.n5433 3.011
R8952 GND.n3886 GND.n3885 3.011
R8953 GND.n3806 GND.n3805 3.011
R8954 GND.n3632 GND.n3631 3.011
R8955 GND.n3689 GND.n3688 3.011
R8956 GND.n14358 GND.n14357 3
R8957 GND.n14315 GND.n14314 3
R8958 GND.n14306 GND.n14305 3
R8959 GND.n14299 GND.n14298 3
R8960 GND.n2457 GND.n2456 3
R8961 GND.n2417 GND.n2416 3
R8962 GND.n2407 GND.n2406 3
R8963 GND.n2400 GND.n2399 3
R8964 GND.n2198 GND.n2197 3
R8965 GND.n2158 GND.n2157 3
R8966 GND.n2149 GND.n2148 3
R8967 GND.n2142 GND.n2141 3
R8968 GND.n14630 GND.n14628 3
R8969 GND.n14631 GND.n14589 3
R8970 GND.n14633 GND.n14582 3
R8971 GND.n14634 GND.n14576 3
R8972 GND.n6402 GND.n6383 2.989
R8973 GND.n2386 GND.n2296 2.989
R8974 GND.n6402 GND.n6359 2.987
R8975 GND.n6467 GND.n6412 2.987
R8976 GND.n6651 GND.n6590 2.987
R8977 GND.n2386 GND.n2385 2.987
R8978 GND.n16412 GND.n16409 2.987
R8979 GND.n16673 GND.n16670 2.987
R8980 GND.n16934 GND.n16931 2.987
R8981 GND.n17195 GND.n17192 2.987
R8982 GND.n17456 GND.n17453 2.987
R8983 GND.n2386 GND.n2329 2.979
R8984 GND.n6402 GND.n6401 2.979
R8985 GND.n15594 GND.n15588 2.635
R8986 GND.n15678 GND.n15672 2.635
R8987 GND.n11271 GND.n11266 2.635
R8988 GND.n11191 GND.n11186 2.635
R8989 GND.n13678 GND.n13673 2.635
R8990 GND.n13598 GND.n13593 2.635
R8991 GND.n13382 GND.n13376 2.635
R8992 GND.n13466 GND.n13460 2.635
R8993 GND.n12659 GND.n12653 2.635
R8994 GND.n12575 GND.n12569 2.635
R8995 GND.n13099 GND.n13094 2.635
R8996 GND.n13179 GND.n13178 2.635
R8997 GND.n12882 GND.n12879 2.635
R8998 GND.n12882 GND.n12881 2.635
R8999 GND.n12956 GND.n12950 2.635
R9000 GND.n11994 GND.n11989 2.635
R9001 GND.n12063 GND.n12062 2.635
R9002 GND.n11798 GND.n11795 2.635
R9003 GND.n11798 GND.n11797 2.635
R9004 GND.n11852 GND.n11847 2.635
R9005 GND.n12232 GND.n12227 2.635
R9006 GND.n12167 GND.n12166 2.635
R9007 GND.n12439 GND.n12436 2.635
R9008 GND.n12439 GND.n12438 2.635
R9009 GND.n12376 GND.n12370 2.635
R9010 GND.n7721 GND.n7716 2.635
R9011 GND.n7674 GND.n7673 2.635
R9012 GND.n7943 GND.n7940 2.635
R9013 GND.n7943 GND.n7942 2.635
R9014 GND.n7863 GND.n7858 2.635
R9015 GND.n7333 GND.n7328 2.635
R9016 GND.n7249 GND.n7244 2.635
R9017 GND.n6290 GND.n6285 2.635
R9018 GND.n6210 GND.n6205 2.635
R9019 GND.n7032 GND.n7026 2.635
R9020 GND.n7116 GND.n7110 2.635
R9021 GND.n8107 GND.n8101 2.635
R9022 GND.n8023 GND.n8017 2.635
R9023 GND.n15975 GND.n15970 2.635
R9024 GND.n16036 GND.n16035 2.635
R9025 GND.n16212 GND.n16209 2.635
R9026 GND.n16212 GND.n16211 2.635
R9027 GND.n16149 GND.n16144 2.635
R9028 GND.n1098 GND.n1093 2.635
R9029 GND.n1034 GND.n1033 2.635
R9030 GND.n867 GND.n864 2.635
R9031 GND.n867 GND.n866 2.635
R9032 GND.n923 GND.n917 2.635
R9033 GND.n9675 GND.n9670 2.635
R9034 GND.n9736 GND.n9735 2.635
R9035 GND.n9912 GND.n9909 2.635
R9036 GND.n9912 GND.n9911 2.635
R9037 GND.n9849 GND.n9844 2.635
R9038 GND.n1266 GND.n1261 2.635
R9039 GND.n1326 GND.n1325 2.635
R9040 GND.n1505 GND.n1502 2.635
R9041 GND.n1505 GND.n1504 2.635
R9042 GND.n1442 GND.n1436 2.635
R9043 GND.n10267 GND.n10262 2.635
R9044 GND.n10183 GND.n10178 2.635
R9045 GND.n10092 GND.n10087 2.635
R9046 GND.n10012 GND.n10007 2.635
R9047 GND.n8831 GND.n8826 2.635
R9048 GND.n8751 GND.n8746 2.635
R9049 GND.n8537 GND.n8532 2.635
R9050 GND.n8453 GND.n8448 2.635
R9051 GND.n8974 GND.n8969 2.635
R9052 GND.n9035 GND.n9034 2.635
R9053 GND.n9211 GND.n9208 2.635
R9054 GND.n9211 GND.n9210 2.635
R9055 GND.n9148 GND.n9143 2.635
R9056 GND.n5717 GND.n5712 2.635
R9057 GND.n5653 GND.n5652 2.635
R9058 GND.n5486 GND.n5483 2.635
R9059 GND.n5486 GND.n5485 2.635
R9060 GND.n5542 GND.n5536 2.635
R9061 GND.n4459 GND.n4454 2.635
R9062 GND.n4394 GND.n4393 2.635
R9063 GND.n4227 GND.n4224 2.635
R9064 GND.n4227 GND.n4226 2.635
R9065 GND.n4283 GND.n4277 2.635
R9066 GND.n4709 GND.n4703 2.635
R9067 GND.n4625 GND.n4619 2.635
R9068 GND.n5055 GND.n5049 2.635
R9069 GND.n4971 GND.n4965 2.635
R9070 GND.n3026 GND.n3021 2.635
R9071 GND.n3106 GND.n3101 2.635
R9072 GND.n3226 GND.n3221 2.635
R9073 GND.n3306 GND.n3301 2.635
R9074 GND.n10450 GND.n10445 2.635
R9075 GND.n10530 GND.n10525 2.635
R9076 GND.n14871 GND.n14865 2.635
R9077 GND.n14787 GND.n14781 2.635
R9078 GND.n15157 GND.n15152 2.635
R9079 GND.n15237 GND.n15232 2.635
R9080 GND.n3879 GND.n3874 2.635
R9081 GND.n3815 GND.n3814 2.635
R9082 GND.n3652 GND.n3649 2.635
R9083 GND.n3652 GND.n3651 2.635
R9084 GND.n3706 GND.n3701 2.635
R9085 GND.n4057 GND.n4056 2.56
R9086 GND.n2740 GND.n2739 2.56
R9087 GND.n16569 GND.n16511 2.469
R9088 GND.n16830 GND.n16772 2.469
R9089 GND.n17091 GND.n17033 2.469
R9090 GND.n17352 GND.n17294 2.469
R9091 GND.n17613 GND.n17555 2.469
R9092 GND.n785 GND.n732 2.469
R9093 GND.n702 GND.n701 2.469
R9094 GND.n527 GND.n474 2.469
R9095 GND.n444 GND.n443 2.469
R9096 GND.n269 GND.n216 2.469
R9097 GND.n186 GND.n185 2.469
R9098 GND.n17804 GND.n17726 2.469
R9099 GND.n17801 GND.n17800 2.469
R9100 GND.n16569 GND.n16529 2.468
R9101 GND.n16483 GND.n16482 2.468
R9102 GND.n16830 GND.n16790 2.468
R9103 GND.n16744 GND.n16743 2.468
R9104 GND.n17091 GND.n17051 2.468
R9105 GND.n17005 GND.n17004 2.468
R9106 GND.n17352 GND.n17312 2.468
R9107 GND.n17266 GND.n17265 2.468
R9108 GND.n17613 GND.n17573 2.468
R9109 GND.n17527 GND.n17526 2.468
R9110 GND.n15563 GND.n15562 2.258
R9111 GND.n15697 GND.n15696 2.258
R9112 GND.n11290 GND.n11289 2.258
R9113 GND.n11162 GND.n11161 2.258
R9114 GND.n13697 GND.n13696 2.258
R9115 GND.n13569 GND.n13568 2.258
R9116 GND.n13351 GND.n13350 2.258
R9117 GND.n13485 GND.n13484 2.258
R9118 GND.n12678 GND.n12677 2.258
R9119 GND.n12544 GND.n12543 2.258
R9120 GND.n13118 GND.n13117 2.258
R9121 GND.n13171 GND.n13170 2.258
R9122 GND.n12865 GND.n12864 2.258
R9123 GND.n12925 GND.n12924 2.258
R9124 GND.n12014 GND.n12013 2.258
R9125 GND.n12077 GND.n12076 2.258
R9126 GND.n11804 GND.n11803 2.258
R9127 GND.n11822 GND.n11821 2.258
R9128 GND.n12202 GND.n12201 2.258
R9129 GND.n12181 GND.n12180 2.258
R9130 GND.n12422 GND.n12421 2.258
R9131 GND.n12395 GND.n12394 2.258
R9132 GND.n7692 GND.n7691 2.258
R9133 GND.n7666 GND.n7665 2.258
R9134 GND.n7949 GND.n7948 2.258
R9135 GND.n7883 GND.n7882 2.258
R9136 GND.n7591 GND.n7588 2.258
R9137 GND.n7353 GND.n7352 2.258
R9138 GND.n7219 GND.n7218 2.258
R9139 GND.n6309 GND.n6308 2.258
R9140 GND.n6180 GND.n6179 2.258
R9141 GND.n7971 GND.n7968 2.258
R9142 GND.n7001 GND.n7000 2.258
R9143 GND.n7135 GND.n7134 2.258
R9144 GND.n8126 GND.n8125 2.258
R9145 GND.n7992 GND.n7991 2.258
R9146 GND.n15945 GND.n15944 2.258
R9147 GND.n16051 GND.n16050 2.258
R9148 GND.n16218 GND.n16217 2.258
R9149 GND.n16168 GND.n16167 2.258
R9150 GND.n1117 GND.n1116 2.258
R9151 GND.n1017 GND.n1016 2.258
R9152 GND.n850 GND.n849 2.258
R9153 GND.n892 GND.n891 2.258
R9154 GND.n9645 GND.n9644 2.258
R9155 GND.n9751 GND.n9750 2.258
R9156 GND.n9918 GND.n9917 2.258
R9157 GND.n9868 GND.n9867 2.258
R9158 GND.n1237 GND.n1236 2.258
R9159 GND.n1341 GND.n1340 2.258
R9160 GND.n1488 GND.n1487 2.258
R9161 GND.n1461 GND.n1460 2.258
R9162 GND.n10287 GND.n10286 2.258
R9163 GND.n10153 GND.n10152 2.258
R9164 GND.n10111 GND.n10110 2.258
R9165 GND.n9982 GND.n9981 2.258
R9166 GND.n8850 GND.n8849 2.258
R9167 GND.n8722 GND.n8721 2.258
R9168 GND.n8557 GND.n8556 2.258
R9169 GND.n8423 GND.n8422 2.258
R9170 GND.n8944 GND.n8943 2.258
R9171 GND.n9050 GND.n9049 2.258
R9172 GND.n9217 GND.n9216 2.258
R9173 GND.n9167 GND.n9166 2.258
R9174 GND.n5736 GND.n5735 2.258
R9175 GND.n5636 GND.n5635 2.258
R9176 GND.n5469 GND.n5468 2.258
R9177 GND.n5511 GND.n5510 2.258
R9178 GND.n4479 GND.n4478 2.258
R9179 GND.n4377 GND.n4376 2.258
R9180 GND.n4210 GND.n4209 2.258
R9181 GND.n4252 GND.n4251 2.258
R9182 GND.n4728 GND.n4727 2.258
R9183 GND.n4594 GND.n4593 2.258
R9184 GND.n5074 GND.n5073 2.258
R9185 GND.n4940 GND.n4939 2.258
R9186 GND.n2997 GND.n2996 2.258
R9187 GND.n3125 GND.n3124 2.258
R9188 GND.n3197 GND.n3196 2.258
R9189 GND.n3325 GND.n3324 2.258
R9190 GND.n10329 GND.n10326 2.258
R9191 GND.n10421 GND.n10420 2.258
R9192 GND.n10549 GND.n10548 2.258
R9193 GND.n14890 GND.n14889 2.258
R9194 GND.n14756 GND.n14755 2.258
R9195 GND.n15128 GND.n15127 2.258
R9196 GND.n15257 GND.n15256 2.258
R9197 GND.n9961 GND.n9958 2.258
R9198 GND.n3898 GND.n3897 2.258
R9199 GND.n3798 GND.n3797 2.258
R9200 GND.n3658 GND.n3657 2.258
R9201 GND.n3676 GND.n3675 2.258
R9202 GND.n2682 GND.n2681 2.25
R9203 GND.n2687 GND.n2686 2.25
R9204 GND.n2692 GND.n2691 2.25
R9205 GND.n2697 GND.n2696 2.25
R9206 GND.n2702 GND.n2701 2.25
R9207 GND.n3997 GND.n3996 2.25
R9208 GND.n2710 GND.n2709 2.25
R9209 GND.n2715 GND.n2714 2.25
R9210 GND.n2720 GND.n2719 2.25
R9211 GND.n2725 GND.n2724 2.25
R9212 GND.n2727 GND.n2726 2.25
R9213 GND.n2747 GND.n2746 2.25
R9214 GND.n2756 GND.n2755 2.25
R9215 GND.n2761 GND.n2760 2.25
R9216 GND.n2766 GND.n2765 2.25
R9217 GND.n2771 GND.n2770 2.25
R9218 GND.n4107 GND.n4106 2.25
R9219 GND.n2779 GND.n2778 2.25
R9220 GND.n2784 GND.n2783 2.25
R9221 GND.n2789 GND.n2788 2.25
R9222 GND.n2794 GND.n2793 2.25
R9223 GND.n2799 GND.n2798 2.25
R9224 GND.n4040 GND.n4039 2.25
R9225 GND.n4039 GND.n4038 2.25
R9226 GND.n4030 GND.n4029 2.25
R9227 GND.n4029 GND.n4028 2.25
R9228 GND.n4016 GND.n4015 2.25
R9229 GND.n4015 GND.n4014 2.25
R9230 GND.n3995 GND.n3994 2.25
R9231 GND.n3994 GND.n3993 2.25
R9232 GND.n3981 GND.n3980 2.25
R9233 GND.n3980 GND.n3979 2.25
R9234 GND.n3967 GND.n3966 2.25
R9235 GND.n3966 GND.n3965 2.25
R9236 GND.n3974 GND.n3973 2.25
R9237 GND.n3973 GND.n3972 2.25
R9238 GND.n3988 GND.n3987 2.25
R9239 GND.n3987 GND.n3986 2.25
R9240 GND.n4009 GND.n4008 2.25
R9241 GND.n4008 GND.n4007 2.25
R9242 GND.n4023 GND.n4022 2.25
R9243 GND.n4022 GND.n4021 2.25
R9244 GND.n4037 GND.n4036 2.25
R9245 GND.n4036 GND.n4035 2.25
R9246 GND.n4147 GND.n4146 2.25
R9247 GND.n4146 GND.n4145 2.25
R9248 GND.n4140 GND.n4139 2.25
R9249 GND.n4139 GND.n4138 2.25
R9250 GND.n4133 GND.n4132 2.25
R9251 GND.n4132 GND.n4131 2.25
R9252 GND.n4126 GND.n4125 2.25
R9253 GND.n4125 GND.n4124 2.25
R9254 GND.n4119 GND.n4118 2.25
R9255 GND.n4118 GND.n4117 2.25
R9256 GND.n4105 GND.n4104 2.25
R9257 GND.n4104 GND.n4103 2.25
R9258 GND.n4098 GND.n4097 2.25
R9259 GND.n4097 GND.n4096 2.25
R9260 GND.n4091 GND.n4090 2.25
R9261 GND.n4090 GND.n4089 2.25
R9262 GND.n4084 GND.n4083 2.25
R9263 GND.n4083 GND.n4082 2.25
R9264 GND.n4077 GND.n4076 2.25
R9265 GND.n4076 GND.n4075 2.25
R9266 GND.n4065 GND.n4064 2.25
R9267 GND.n4064 GND.n4063 2.25
R9268 GND.n3488 GND.n2204 2.249
R9269 GND.n15454 GND.n15453 2.249
R9270 GND.n14185 GND.n14184 2.248
R9271 GND.n3485 GND.n2205 2.248
R9272 GND.n2027 GND.n2026 2.248
R9273 GND.n14530 GND.n14528 2.248
R9274 GND.n1606 GND.n1605 2.248
R9275 GND.n10835 GND.n10832 2.231
R9276 GND.n11496 GND.n11493 2.231
R9277 GND.n16393 GND.n16392 2.231
R9278 GND.n16567 GND.n16566 2.231
R9279 GND.n16654 GND.n16653 2.231
R9280 GND.n16828 GND.n16827 2.231
R9281 GND.n16915 GND.n16914 2.231
R9282 GND.n17089 GND.n17088 2.231
R9283 GND.n17176 GND.n17175 2.231
R9284 GND.n17350 GND.n17349 2.231
R9285 GND.n17437 GND.n17436 2.231
R9286 GND.n17611 GND.n17610 2.231
R9287 GND.n614 GND.n613 2.231
R9288 GND.n680 GND.n679 2.231
R9289 GND.n783 GND.n782 2.231
R9290 GND.n356 GND.n355 2.231
R9291 GND.n422 GND.n421 2.231
R9292 GND.n525 GND.n524 2.231
R9293 GND.n98 GND.n97 2.231
R9294 GND.n164 GND.n163 2.231
R9295 GND.n267 GND.n266 2.231
R9296 GND.n17934 GND.n17933 2.231
R9297 GND.n17779 GND.n17778 2.231
R9298 GND.n17856 GND.n17855 2.231
R9299 GND.n13799 GND.n13798 2.231
R9300 GND.n12779 GND.n12538 2.231
R9301 GND.n11041 GND.n11040 2.231
R9302 GND.n8230 GND.n8227 2.231
R9303 GND.n8318 GND.n8235 2.231
R9304 GND.n7501 GND.n7500 2.231
R9305 GND.n7520 GND.n7513 2.231
R9306 GND.n5167 GND.n1927 2.231
R9307 GND.n2559 GND.n2461 2.231
R9308 GND.n4856 GND.n3497 2.231
R9309 GND.n15464 GND.n15463 2.231
R9310 GND.n15050 GND.n15001 2.231
R9311 GND.n13931 GND.n10842 2.231
R9312 GND.n13793 GND.n13790 2.231
R9313 GND.n11553 GND.n11503 2.231
R9314 GND.n11386 GND.n11010 2.231
R9315 GND.n2896 GND.n2846 2.231
R9316 GND.n14989 GND.n14988 2.231
R9317 GND.n7090 GND.n7089 2.163
R9318 GND.n7115 GND.n7114 2.163
R9319 GND.n7140 GND.n7139 2.163
R9320 GND.n8047 GND.n8046 2.163
R9321 GND.n8022 GND.n8021 2.163
R9322 GND.n7997 GND.n7996 2.163
R9323 GND.n7875 GND.n7874 2.163
R9324 GND.n13440 GND.n13439 2.163
R9325 GND.n13465 GND.n13464 2.163
R9326 GND.n13490 GND.n13489 2.163
R9327 GND.n12599 GND.n12598 2.163
R9328 GND.n12574 GND.n12573 2.163
R9329 GND.n12549 GND.n12548 2.163
R9330 GND.n12633 GND.n12632 2.163
R9331 GND.n12658 GND.n12657 2.163
R9332 GND.n12683 GND.n12682 2.163
R9333 GND.n13356 GND.n13355 2.163
R9334 GND.n13381 GND.n13380 2.163
R9335 GND.n13406 GND.n13405 2.163
R9336 GND.n12979 GND.n12978 2.163
R9337 GND.n12955 GND.n12954 2.163
R9338 GND.n12930 GND.n12929 2.163
R9339 GND.n12042 GND.n12041 2.163
R9340 GND.n12058 GND.n12057 2.163
R9341 GND.n12073 GND.n12072 2.163
R9342 GND.n12006 GND.n12005 2.163
R9343 GND.n11981 GND.n11980 2.163
R9344 GND.n12033 GND.n12032 2.163
R9345 GND.n11839 GND.n11838 2.163
R9346 GND.n11826 GND.n11825 2.163
R9347 GND.n12146 GND.n12145 2.163
R9348 GND.n12162 GND.n12161 2.163
R9349 GND.n12177 GND.n12176 2.163
R9350 GND.n12350 GND.n12349 2.163
R9351 GND.n12375 GND.n12374 2.163
R9352 GND.n12400 GND.n12399 2.163
R9353 GND.n12219 GND.n12218 2.163
R9354 GND.n12244 GND.n12243 2.163
R9355 GND.n12137 GND.n12136 2.163
R9356 GND.n12425 GND.n12424 2.163
R9357 GND.n12441 GND.n12440 2.163
R9358 GND.n12458 GND.n12457 2.163
R9359 GND.n12868 GND.n12867 2.163
R9360 GND.n12884 GND.n12883 2.163
R9361 GND.n12901 GND.n12900 2.163
R9362 GND.n8131 GND.n8130 2.163
R9363 GND.n8106 GND.n8105 2.163
R9364 GND.n8081 GND.n8080 2.163
R9365 GND.n7006 GND.n7005 2.163
R9366 GND.n7031 GND.n7030 2.163
R9367 GND.n7056 GND.n7055 2.163
R9368 GND.n7286 GND.n7285 2.163
R9369 GND.n7261 GND.n7260 2.163
R9370 GND.n7236 GND.n7235 2.163
R9371 GND.n6185 GND.n6184 2.163
R9372 GND.n7295 GND.n7294 2.163
R9373 GND.n7320 GND.n7319 2.163
R9374 GND.n7345 GND.n7344 2.163
R9375 GND.n14811 GND.n14810 2.163
R9376 GND.n14786 GND.n14785 2.163
R9377 GND.n14761 GND.n14760 2.163
R9378 GND.n8908 GND.n8907 2.163
R9379 GND.n8917 GND.n8916 2.163
R9380 GND.n8926 GND.n8925 2.163
R9381 GND.n9609 GND.n9608 2.163
R9382 GND.n9618 GND.n9617 2.163
R9383 GND.n9627 GND.n9626 2.163
R9384 GND.n15909 GND.n15908 2.163
R9385 GND.n15918 GND.n15917 2.163
R9386 GND.n15927 GND.n15926 2.163
R9387 GND.n15904 GND.n15903 2.163
R9388 GND.n15987 GND.n15986 2.163
R9389 GND.n15962 GND.n15961 2.163
R9390 GND.n16173 GND.n16172 2.163
R9391 GND.n947 GND.n946 2.163
R9392 GND.n922 GND.n921 2.163
R9393 GND.n897 GND.n896 2.163
R9394 GND.n881 GND.n880 2.163
R9395 GND.n869 GND.n868 2.163
R9396 GND.n853 GND.n852 2.163
R9397 GND.n9604 GND.n9603 2.163
R9398 GND.n9687 GND.n9686 2.163
R9399 GND.n9662 GND.n9661 2.163
R9400 GND.n9873 GND.n9872 2.163
R9401 GND.n1416 GND.n1415 2.163
R9402 GND.n1441 GND.n1440 2.163
R9403 GND.n1466 GND.n1465 2.163
R9404 GND.n1519 GND.n1518 2.163
R9405 GND.n1507 GND.n1506 2.163
R9406 GND.n1491 GND.n1490 2.163
R9407 GND.n10220 GND.n10219 2.163
R9408 GND.n10195 GND.n10194 2.163
R9409 GND.n10170 GND.n10169 2.163
R9410 GND.n10229 GND.n10228 2.163
R9411 GND.n10254 GND.n10253 2.163
R9412 GND.n10279 GND.n10278 2.163
R9413 GND.n8490 GND.n8489 2.163
R9414 GND.n8465 GND.n8464 2.163
R9415 GND.n8440 GND.n8439 2.163
R9416 GND.n8549 GND.n8548 2.163
R9417 GND.n8524 GND.n8523 2.163
R9418 GND.n8499 GND.n8498 2.163
R9419 GND.n9987 GND.n9986 2.163
R9420 GND.n8903 GND.n8902 2.163
R9421 GND.n8986 GND.n8985 2.163
R9422 GND.n8961 GND.n8960 2.163
R9423 GND.n9172 GND.n9171 2.163
R9424 GND.n5566 GND.n5565 2.163
R9425 GND.n5541 GND.n5540 2.163
R9426 GND.n5516 GND.n5515 2.163
R9427 GND.n4504 GND.n4503 2.163
R9428 GND.n4513 GND.n4512 2.163
R9429 GND.n4522 GND.n4521 2.163
R9430 GND.n4307 GND.n4306 2.163
R9431 GND.n4282 GND.n4281 2.163
R9432 GND.n4257 GND.n4256 2.163
R9433 GND.n4241 GND.n4240 2.163
R9434 GND.n4229 GND.n4228 2.163
R9435 GND.n4213 GND.n4212 2.163
R9436 GND.n4499 GND.n4498 2.163
R9437 GND.n4446 GND.n4445 2.163
R9438 GND.n4471 GND.n4470 2.163
R9439 GND.n15652 GND.n15651 2.163
R9440 GND.n15677 GND.n15676 2.163
R9441 GND.n15702 GND.n15701 2.163
R9442 GND.n4649 GND.n4648 2.163
R9443 GND.n4624 GND.n4623 2.163
R9444 GND.n4599 GND.n4598 2.163
R9445 GND.n4995 GND.n4994 2.163
R9446 GND.n4970 GND.n4969 2.163
R9447 GND.n4945 GND.n4944 2.163
R9448 GND.n5029 GND.n5028 2.163
R9449 GND.n5054 GND.n5053 2.163
R9450 GND.n5079 GND.n5078 2.163
R9451 GND.n4683 GND.n4682 2.163
R9452 GND.n4708 GND.n4707 2.163
R9453 GND.n4733 GND.n4732 2.163
R9454 GND.n3130 GND.n3129 2.163
R9455 GND.n3330 GND.n3329 2.163
R9456 GND.n14845 GND.n14844 2.163
R9457 GND.n14870 GND.n14869 2.163
R9458 GND.n14895 GND.n14894 2.163
R9459 GND.n15618 GND.n15617 2.163
R9460 GND.n15593 GND.n15592 2.163
R9461 GND.n15568 GND.n15567 2.163
R9462 GND.n15249 GND.n15248 2.163
R9463 GND.n15261 GND.n15260 2.163
R9464 GND.n3681 GND.n3680 2.163
R9465 GND.n5500 GND.n5499 2.163
R9466 GND.n5488 GND.n5487 2.163
R9467 GND.n5472 GND.n5471 2.163
R9468 GND.n15606 GND.n15601 1.882
R9469 GND.n15665 GND.n15660 1.882
R9470 GND.n11259 GND.n11254 1.882
R9471 GND.n11203 GND.n11198 1.882
R9472 GND.n13666 GND.n13661 1.882
R9473 GND.n13610 GND.n13605 1.882
R9474 GND.n13394 GND.n13389 1.882
R9475 GND.n13453 GND.n13448 1.882
R9476 GND.n12646 GND.n12641 1.882
R9477 GND.n12587 GND.n12582 1.882
R9478 GND.n13087 GND.n13082 1.882
R9479 GND.n13151 GND.n13150 1.882
R9480 GND.n12888 GND.n12885 1.882
R9481 GND.n12888 GND.n12887 1.882
R9482 GND.n12968 GND.n12963 1.882
R9483 GND.n11982 GND.n11976 1.882
R9484 GND.n12056 GND.n12055 1.882
R9485 GND.n11770 GND.n11767 1.882
R9486 GND.n11770 GND.n11769 1.882
R9487 GND.n11864 GND.n11859 1.882
R9488 GND.n12245 GND.n12239 1.882
R9489 GND.n12160 GND.n12159 1.882
R9490 GND.n12445 GND.n12442 1.882
R9491 GND.n12445 GND.n12444 1.882
R9492 GND.n12363 GND.n12358 1.882
R9493 GND.n7733 GND.n7728 1.882
R9494 GND.n7646 GND.n7645 1.882
R9495 GND.n7915 GND.n7912 1.882
R9496 GND.n7915 GND.n7914 1.882
R9497 GND.n7851 GND.n7846 1.882
R9498 GND.n7321 GND.n7315 1.882
R9499 GND.n7262 GND.n7256 1.882
R9500 GND.n6278 GND.n6273 1.882
R9501 GND.n6222 GND.n6217 1.882
R9502 GND.n7044 GND.n7039 1.882
R9503 GND.n7103 GND.n7098 1.882
R9504 GND.n8094 GND.n8089 1.882
R9505 GND.n8035 GND.n8030 1.882
R9506 GND.n15988 GND.n15982 1.882
R9507 GND.n16028 GND.n16027 1.882
R9508 GND.n16200 GND.n16198 1.882
R9509 GND.n16200 GND.n16199 1.882
R9510 GND.n16137 GND.n16132 1.882
R9511 GND.n1086 GND.n1081 1.882
R9512 GND.n1042 GND.n1041 1.882
R9513 GND.n872 GND.n870 1.882
R9514 GND.n872 GND.n871 1.882
R9515 GND.n935 GND.n930 1.882
R9516 GND.n9688 GND.n9682 1.882
R9517 GND.n9728 GND.n9727 1.882
R9518 GND.n9900 GND.n9898 1.882
R9519 GND.n9900 GND.n9899 1.882
R9520 GND.n9837 GND.n9832 1.882
R9521 GND.n1278 GND.n1273 1.882
R9522 GND.n1318 GND.n1317 1.882
R9523 GND.n1510 GND.n1508 1.882
R9524 GND.n1510 GND.n1509 1.882
R9525 GND.n1429 GND.n1424 1.882
R9526 GND.n10255 GND.n10249 1.882
R9527 GND.n10196 GND.n10190 1.882
R9528 GND.n10080 GND.n10075 1.882
R9529 GND.n10024 GND.n10019 1.882
R9530 GND.n8819 GND.n8814 1.882
R9531 GND.n8763 GND.n8758 1.882
R9532 GND.n8525 GND.n8519 1.882
R9533 GND.n8466 GND.n8460 1.882
R9534 GND.n8987 GND.n8981 1.882
R9535 GND.n9027 GND.n9026 1.882
R9536 GND.n9199 GND.n9197 1.882
R9537 GND.n9199 GND.n9198 1.882
R9538 GND.n9136 GND.n9131 1.882
R9539 GND.n5705 GND.n5700 1.882
R9540 GND.n5661 GND.n5660 1.882
R9541 GND.n5491 GND.n5489 1.882
R9542 GND.n5491 GND.n5490 1.882
R9543 GND.n5554 GND.n5549 1.882
R9544 GND.n4447 GND.n4441 1.882
R9545 GND.n4402 GND.n4401 1.882
R9546 GND.n4232 GND.n4230 1.882
R9547 GND.n4232 GND.n4231 1.882
R9548 GND.n4295 GND.n4290 1.882
R9549 GND.n4696 GND.n4691 1.882
R9550 GND.n4637 GND.n4632 1.882
R9551 GND.n5042 GND.n5037 1.882
R9552 GND.n4983 GND.n4978 1.882
R9553 GND.n3038 GND.n3033 1.882
R9554 GND.n3094 GND.n3089 1.882
R9555 GND.n3238 GND.n3233 1.882
R9556 GND.n3294 GND.n3289 1.882
R9557 GND.n10462 GND.n10457 1.882
R9558 GND.n10518 GND.n10513 1.882
R9559 GND.n14858 GND.n14853 1.882
R9560 GND.n14799 GND.n14794 1.882
R9561 GND.n15169 GND.n15164 1.882
R9562 GND.n15225 GND.n15220 1.882
R9563 GND.n3867 GND.n3862 1.882
R9564 GND.n3823 GND.n3822 1.882
R9565 GND.n3640 GND.n3638 1.882
R9566 GND.n3640 GND.n3639 1.882
R9567 GND.n3718 GND.n3713 1.882
R9568 GND.n3998 GND.n3997 1.536
R9569 GND.n15551 GND.n15550 1.505
R9570 GND.n15710 GND.n15709 1.505
R9571 GND.n11302 GND.n11301 1.505
R9572 GND.n11149 GND.n11148 1.505
R9573 GND.n13709 GND.n13708 1.505
R9574 GND.n13556 GND.n13555 1.505
R9575 GND.n13339 GND.n13338 1.505
R9576 GND.n13498 GND.n13497 1.505
R9577 GND.n12691 GND.n12690 1.505
R9578 GND.n12518 GND.n12517 1.505
R9579 GND.n13130 GND.n13129 1.505
R9580 GND.n13164 GND.n13163 1.505
R9581 GND.n12855 GND.n12854 1.505
R9582 GND.n12851 GND.n12850 1.505
R9583 GND.n12026 GND.n12025 1.505
R9584 GND.n12085 GND.n12084 1.505
R9585 GND.n11754 GND.n11753 1.505
R9586 GND.n11752 GND.n11751 1.505
R9587 GND.n12130 GND.n12129 1.505
R9588 GND.n12189 GND.n12188 1.505
R9589 GND.n12412 GND.n12411 1.505
R9590 GND.n12408 GND.n12407 1.505
R9591 GND.n7625 GND.n7624 1.505
R9592 GND.n7659 GND.n7658 1.505
R9593 GND.n7899 GND.n7898 1.505
R9594 GND.n7895 GND.n7894 1.505
R9595 GND.n13200 GND.n13197 1.505
R9596 GND.n7365 GND.n7364 1.505
R9597 GND.n7206 GND.n7205 1.505
R9598 GND.n6321 GND.n6320 1.505
R9599 GND.n6167 GND.n6166 1.505
R9600 GND.n12843 GND.n12840 1.505
R9601 GND.n6989 GND.n6988 1.505
R9602 GND.n7148 GND.n7147 1.505
R9603 GND.n8139 GND.n8138 1.505
R9604 GND.n7979 GND.n7978 1.505
R9605 GND.n15896 GND.n15895 1.505
R9606 GND.n16059 GND.n16058 1.505
R9607 GND.n16185 GND.n16184 1.505
R9608 GND.n16181 GND.n16180 1.505
R9609 GND.n1129 GND.n1128 1.505
R9610 GND.n1009 GND.n1008 1.505
R9611 GND.n840 GND.n839 1.505
R9612 GND.n836 GND.n835 1.505
R9613 GND.n9596 GND.n9595 1.505
R9614 GND.n9759 GND.n9758 1.505
R9615 GND.n9885 GND.n9884 1.505
R9616 GND.n9881 GND.n9880 1.505
R9617 GND.n1192 GND.n1191 1.505
R9618 GND.n1349 GND.n1348 1.505
R9619 GND.n1478 GND.n1477 1.505
R9620 GND.n1474 GND.n1473 1.505
R9621 GND.n10299 GND.n10298 1.505
R9622 GND.n10140 GND.n10139 1.505
R9623 GND.n10123 GND.n10122 1.505
R9624 GND.n9969 GND.n9968 1.505
R9625 GND.n8862 GND.n8861 1.505
R9626 GND.n8709 GND.n8708 1.505
R9627 GND.n8569 GND.n8568 1.505
R9628 GND.n8410 GND.n8409 1.505
R9629 GND.n8895 GND.n8894 1.505
R9630 GND.n9058 GND.n9057 1.505
R9631 GND.n9184 GND.n9183 1.505
R9632 GND.n9180 GND.n9179 1.505
R9633 GND.n5748 GND.n5747 1.505
R9634 GND.n5628 GND.n5627 1.505
R9635 GND.n5459 GND.n5458 1.505
R9636 GND.n5455 GND.n5454 1.505
R9637 GND.n4491 GND.n4490 1.505
R9638 GND.n4369 GND.n4368 1.505
R9639 GND.n4200 GND.n4199 1.505
R9640 GND.n4196 GND.n4195 1.505
R9641 GND.n4741 GND.n4740 1.505
R9642 GND.n4581 GND.n4580 1.505
R9643 GND.n5087 GND.n5086 1.505
R9644 GND.n4927 GND.n4926 1.505
R9645 GND.n2985 GND.n2984 1.505
R9646 GND.n3138 GND.n3137 1.505
R9647 GND.n3186 GND.n3185 1.505
R9648 GND.n3338 GND.n3337 1.505
R9649 GND.n15888 GND.n15885 1.505
R9650 GND.n10409 GND.n10408 1.505
R9651 GND.n10561 GND.n10560 1.505
R9652 GND.n14903 GND.n14902 1.505
R9653 GND.n14743 GND.n14742 1.505
R9654 GND.n15115 GND.n15114 1.505
R9655 GND.n15269 GND.n15268 1.505
R9656 GND.n811 GND.n808 1.505
R9657 GND.n3910 GND.n3909 1.505
R9658 GND.n3790 GND.n3789 1.505
R9659 GND.n3625 GND.n3624 1.505
R9660 GND.n3623 GND.n3622 1.505
R9661 GND.n14470 GND.n14469 1.377
R9662 GND.n15303 GND.n15302 1.377
R9663 GND.n14484 GND.n14483 1.377
R9664 GND.n15435 GND.n15434 1.377
R9665 GND.n15745 GND.n15744 1.377
R9666 GND.n15734 GND.n15733 1.377
R9667 GND.n14092 GND.n14091 1.377
R9668 GND.n14109 GND.n14108 1.377
R9669 GND.n2664 GND.n2663 1.377
R9670 GND.n4913 GND.n4912 1.377
R9671 GND.n1950 GND.n1949 1.377
R9672 GND.n4779 GND.n4778 1.377
R9673 GND.n7190 GND.n7189 1.377
R9674 GND.n7179 GND.n7178 1.377
R9675 GND.n7409 GND.n7408 1.377
R9676 GND.n7392 GND.n7391 1.377
R9677 GND.n10777 GND.n10776 1.377
R9678 GND.n13875 GND.n13874 1.377
R9679 GND.n10885 GND.n10884 1.377
R9680 GND.n10896 GND.n10895 1.377
R9681 GND.n11118 GND.n11117 1.377
R9682 GND.n11135 GND.n11134 1.377
R9683 GND.n13526 GND.n13525 1.377
R9684 GND.n13537 GND.n13536 1.377
R9685 GND.n6038 GND.n6037 1.377
R9686 GND.n6055 GND.n6054 1.377
R9687 GND.n8243 GND.n8242 1.377
R9688 GND.n5907 GND.n5906 1.377
R9689 GND.n9270 GND.n9269 1.377
R9690 GND.n9287 GND.n9286 1.377
R9691 GND.n1576 GND.n1575 1.377
R9692 GND.n1692 GND.n1691 1.377
R9693 GND.n3374 GND.n3373 1.377
R9694 GND.n3391 GND.n3390 1.377
R9695 GND.n3170 GND.n3169 1.377
R9696 GND.n2485 GND.n2484 1.377
R9697 GND.n16555 GND.n16554 1.155
R9698 GND.n16816 GND.n16815 1.155
R9699 GND.n17077 GND.n17076 1.155
R9700 GND.n17338 GND.n17337 1.155
R9701 GND.n17599 GND.n17598 1.155
R9702 GND.n771 GND.n770 1.155
R9703 GND.n513 GND.n512 1.155
R9704 GND.n255 GND.n254 1.155
R9705 GND.n17844 GND.n17843 1.155
R9706 GND.n16408 GND.n16407 1.155
R9707 GND.n16381 GND.n16380 1.155
R9708 GND.n16669 GND.n16668 1.155
R9709 GND.n16642 GND.n16641 1.155
R9710 GND.n16930 GND.n16929 1.155
R9711 GND.n16903 GND.n16902 1.155
R9712 GND.n17191 GND.n17190 1.155
R9713 GND.n17164 GND.n17163 1.155
R9714 GND.n17452 GND.n17451 1.155
R9715 GND.n17425 GND.n17424 1.155
R9716 GND.n668 GND.n667 1.155
R9717 GND.n602 GND.n601 1.155
R9718 GND.n410 GND.n409 1.155
R9719 GND.n344 GND.n343 1.155
R9720 GND.n152 GND.n151 1.155
R9721 GND.n86 GND.n85 1.155
R9722 GND.n17767 GND.n17766 1.155
R9723 GND.n17922 GND.n17921 1.155
R9724 GND.n15619 GND.n15613 1.129
R9725 GND.n15653 GND.n15647 1.129
R9726 GND.n11247 GND.n11242 1.129
R9727 GND.n11215 GND.n11210 1.129
R9728 GND.n13654 GND.n13649 1.129
R9729 GND.n13622 GND.n13617 1.129
R9730 GND.n13407 GND.n13401 1.129
R9731 GND.n13441 GND.n13435 1.129
R9732 GND.n12634 GND.n12628 1.129
R9733 GND.n12600 GND.n12594 1.129
R9734 GND.n13075 GND.n13070 1.129
R9735 GND.n13186 GND.n13185 1.129
R9736 GND.n12899 GND.n12896 1.129
R9737 GND.n12899 GND.n12898 1.129
R9738 GND.n12981 GND.n12980 1.129
R9739 GND.n11969 GND.n11964 1.129
R9740 GND.n12048 GND.n12046 1.129
R9741 GND.n12048 GND.n12047 1.129
R9742 GND.n11790 GND.n11787 1.129
R9743 GND.n11790 GND.n11789 1.129
R9744 GND.n11876 GND.n11875 1.129
R9745 GND.n12262 GND.n12257 1.129
R9746 GND.n12152 GND.n12150 1.129
R9747 GND.n12152 GND.n12151 1.129
R9748 GND.n12456 GND.n12453 1.129
R9749 GND.n12456 GND.n12455 1.129
R9750 GND.n12351 GND.n12345 1.129
R9751 GND.n7750 GND.n7745 1.129
R9752 GND.n7681 GND.n7680 1.129
R9753 GND.n7935 GND.n7932 1.129
R9754 GND.n7935 GND.n7934 1.129
R9755 GND.n7839 GND.n7834 1.129
R9756 GND.n7308 GND.n7303 1.129
R9757 GND.n7274 GND.n7269 1.129
R9758 GND.n6266 GND.n6261 1.129
R9759 GND.n6234 GND.n6229 1.129
R9760 GND.n7057 GND.n7051 1.129
R9761 GND.n7091 GND.n7085 1.129
R9762 GND.n8082 GND.n8076 1.129
R9763 GND.n8048 GND.n8042 1.129
R9764 GND.n16005 GND.n16000 1.129
R9765 GND.n16020 GND.n16019 1.129
R9766 GND.n16092 GND.n815 1.129
R9767 GND.n16093 GND.n16092 1.129
R9768 GND.n16125 GND.n16120 1.129
R9769 GND.n1074 GND.n1069 1.129
R9770 GND.n1050 GND.n1049 1.129
R9771 GND.n977 GND.n818 1.129
R9772 GND.n977 GND.n976 1.129
R9773 GND.n948 GND.n942 1.129
R9774 GND.n9705 GND.n9700 1.129
R9775 GND.n9720 GND.n9719 1.129
R9776 GND.n9792 GND.n9592 1.129
R9777 GND.n9793 GND.n9792 1.129
R9778 GND.n9825 GND.n9820 1.129
R9779 GND.n1295 GND.n1290 1.129
R9780 GND.n1310 GND.n1309 1.129
R9781 GND.n1382 GND.n1188 1.129
R9782 GND.n1383 GND.n1382 1.129
R9783 GND.n1417 GND.n1411 1.129
R9784 GND.n10242 GND.n10237 1.129
R9785 GND.n10208 GND.n10203 1.129
R9786 GND.n10068 GND.n10063 1.129
R9787 GND.n10036 GND.n10031 1.129
R9788 GND.n8807 GND.n8802 1.129
R9789 GND.n8775 GND.n8770 1.129
R9790 GND.n8512 GND.n8507 1.129
R9791 GND.n8478 GND.n8473 1.129
R9792 GND.n9004 GND.n8999 1.129
R9793 GND.n9019 GND.n9018 1.129
R9794 GND.n9091 GND.n1907 1.129
R9795 GND.n9092 GND.n9091 1.129
R9796 GND.n9124 GND.n9119 1.129
R9797 GND.n5693 GND.n5688 1.129
R9798 GND.n5669 GND.n5668 1.129
R9799 GND.n5596 GND.n1913 1.129
R9800 GND.n5596 GND.n5595 1.129
R9801 GND.n5567 GND.n5561 1.129
R9802 GND.n4434 GND.n4429 1.129
R9803 GND.n4410 GND.n4409 1.129
R9804 GND.n4337 GND.n4192 1.129
R9805 GND.n4337 GND.n4336 1.129
R9806 GND.n4308 GND.n4302 1.129
R9807 GND.n4684 GND.n4678 1.129
R9808 GND.n4650 GND.n4644 1.129
R9809 GND.n5030 GND.n5024 1.129
R9810 GND.n4996 GND.n4990 1.129
R9811 GND.n3050 GND.n3045 1.129
R9812 GND.n3082 GND.n3077 1.129
R9813 GND.n3250 GND.n3245 1.129
R9814 GND.n3282 GND.n3277 1.129
R9815 GND.n10474 GND.n10469 1.129
R9816 GND.n10506 GND.n10501 1.129
R9817 GND.n14846 GND.n14840 1.129
R9818 GND.n14812 GND.n14806 1.129
R9819 GND.n15181 GND.n15176 1.129
R9820 GND.n15213 GND.n15208 1.129
R9821 GND.n3855 GND.n3850 1.129
R9822 GND.n3831 GND.n3830 1.129
R9823 GND.n3758 GND.n3619 1.129
R9824 GND.n3758 GND.n3757 1.129
R9825 GND.n3730 GND.n3725 1.129
R9826 GND.n9586 GND.n9580 1.035
R9827 GND.n16246 GND.n16240 1.035
R9828 GND.n16246 GND.n16245 1.035
R9829 GND.n9586 GND.n9585 1.035
R9830 GND.n4062 GND.n4061 1.024
R9831 GND.n2745 GND.n2744 1.024
R9832 GND.n16409 GND.n16408 0.921
R9833 GND.n16382 GND.n16381 0.921
R9834 GND.n16670 GND.n16669 0.921
R9835 GND.n16643 GND.n16642 0.921
R9836 GND.n16931 GND.n16930 0.921
R9837 GND.n16904 GND.n16903 0.921
R9838 GND.n17192 GND.n17191 0.921
R9839 GND.n17165 GND.n17164 0.921
R9840 GND.n17453 GND.n17452 0.921
R9841 GND.n17426 GND.n17425 0.921
R9842 GND.n669 GND.n668 0.921
R9843 GND.n603 GND.n602 0.921
R9844 GND.n411 GND.n410 0.921
R9845 GND.n345 GND.n344 0.921
R9846 GND.n153 GND.n152 0.921
R9847 GND.n87 GND.n86 0.921
R9848 GND.n17768 GND.n17767 0.921
R9849 GND.n17923 GND.n17922 0.921
R9850 GND.n16556 GND.n16555 0.903
R9851 GND.n16817 GND.n16816 0.903
R9852 GND.n17078 GND.n17077 0.903
R9853 GND.n17339 GND.n17338 0.903
R9854 GND.n17600 GND.n17599 0.903
R9855 GND.n772 GND.n771 0.903
R9856 GND.n514 GND.n513 0.903
R9857 GND.n256 GND.n255 0.903
R9858 GND.n17845 GND.n17844 0.903
R9859 GND.n16067 GND.n16065 0.818
R9860 GND.n1005 GND.n1003 0.818
R9861 GND.n9767 GND.n9765 0.818
R9862 GND.n1357 GND.n1355 0.818
R9863 GND.n9066 GND.n9064 0.818
R9864 GND.n4365 GND.n4363 0.818
R9865 GND.n3786 GND.n3784 0.818
R9866 GND.n5624 GND.n5622 0.818
R9867 GND.n4049 GND.n4046 0.768
R9868 GND.n2735 GND.n2732 0.768
R9869 GND.n14471 GND.n14466 0.752
R9870 GND.n15304 GND.n15300 0.752
R9871 GND.n14485 GND.n14480 0.752
R9872 GND.n15436 GND.n15431 0.752
R9873 GND.n15746 GND.n15741 0.752
R9874 GND.n15735 GND.n15730 0.752
R9875 GND.n14093 GND.n14088 0.752
R9876 GND.n14110 GND.n14105 0.752
R9877 GND.n2665 GND.n2660 0.752
R9878 GND.n4914 GND.n4909 0.752
R9879 GND.n1951 GND.n1946 0.752
R9880 GND.n4780 GND.n4775 0.752
R9881 GND.n7191 GND.n7186 0.752
R9882 GND.n7180 GND.n7175 0.752
R9883 GND.n7410 GND.n7405 0.752
R9884 GND.n7393 GND.n7388 0.752
R9885 GND.n10778 GND.n10773 0.752
R9886 GND.n13876 GND.n13871 0.752
R9887 GND.n10886 GND.n10881 0.752
R9888 GND.n10897 GND.n10892 0.752
R9889 GND.n11119 GND.n11114 0.752
R9890 GND.n11136 GND.n11131 0.752
R9891 GND.n13527 GND.n13522 0.752
R9892 GND.n13538 GND.n13533 0.752
R9893 GND.n6039 GND.n6034 0.752
R9894 GND.n6056 GND.n6052 0.752
R9895 GND.n8244 GND.n8239 0.752
R9896 GND.n5908 GND.n5903 0.752
R9897 GND.n9271 GND.n9266 0.752
R9898 GND.n9288 GND.n9283 0.752
R9899 GND.n1577 GND.n1572 0.752
R9900 GND.n1693 GND.n1688 0.752
R9901 GND.n3375 GND.n3370 0.752
R9902 GND.n3392 GND.n3387 0.752
R9903 GND.n3171 GND.n3166 0.752
R9904 GND.n2486 GND.n2481 0.752
R9905 GND.n3343 GND.n3342 0.644
R9906 GND.n6993 GND.n6992 0.644
R9907 GND.n7153 GND.n7152 0.644
R9908 GND.n8143 GND.n8142 0.644
R9909 GND.n7957 GND.n7956 0.644
R9910 GND.n13502 GND.n13501 0.644
R9911 GND.n12695 GND.n12694 0.644
R9912 GND.n12860 GND.n12857 0.644
R9913 GND.n12090 GND.n12089 0.644
R9914 GND.n11814 GND.n11813 0.644
R9915 GND.n11759 GND.n11756 0.644
R9916 GND.n12194 GND.n12193 0.644
R9917 GND.n12417 GND.n12414 0.644
R9918 GND.n12474 GND.n12473 0.644
R9919 GND.n12917 GND.n12916 0.644
R9920 GND.n7904 GND.n7901 0.644
R9921 GND.n7984 GND.n7983 0.644
R9922 GND.n7369 GND.n7368 0.644
R9923 GND.n6172 GND.n6171 0.644
R9924 GND.n6325 GND.n6324 0.644
R9925 GND.n11306 GND.n11305 0.644
R9926 GND.n13713 GND.n13712 0.644
R9927 GND.n14907 GND.n14906 0.644
R9928 GND.n9225 GND.n9224 0.644
R9929 GND.n9926 GND.n9925 0.644
R9930 GND.n16226 GND.n16225 0.644
R9931 GND.n16190 GND.n16187 0.644
R9932 GND.n845 GND.n842 0.644
R9933 GND.n884 GND.n883 0.644
R9934 GND.n9890 GND.n9887 0.644
R9935 GND.n1483 GND.n1480 0.644
R9936 GND.n1522 GND.n1521 0.644
R9937 GND.n8573 GND.n8572 0.644
R9938 GND.n9974 GND.n9973 0.644
R9939 GND.n9189 GND.n9186 0.644
R9940 GND.n5464 GND.n5461 0.644
R9941 GND.n4205 GND.n4202 0.644
R9942 GND.n4244 GND.n4243 0.644
R9943 GND.n15555 GND.n15554 0.644
R9944 GND.n15273 GND.n15272 0.644
R9945 GND.n4745 GND.n4744 0.644
R9946 GND.n5091 GND.n5090 0.644
R9947 GND.n4932 GND.n4931 0.644
R9948 GND.n4586 GND.n4585 0.644
R9949 GND.n2989 GND.n2988 0.644
R9950 GND.n14748 GND.n14747 0.644
R9951 GND.n15715 GND.n15714 0.644
R9952 GND.n15120 GND.n15119 0.644
R9953 GND.n3630 GND.n3627 0.644
R9954 GND.n3668 GND.n3667 0.644
R9955 GND.n5503 GND.n5502 0.644
R9956 GND.n5427 GND.n5249 0.583
R9957 GND.n12018 GND.n12017 0.551
R9958 GND.n12080 GND.n12079 0.551
R9959 GND.n11809 GND.n11806 0.551
R9960 GND.n12206 GND.n12205 0.551
R9961 GND.n12184 GND.n12183 0.551
R9962 GND.n13122 GND.n13121 0.551
R9963 GND.n7696 GND.n7695 0.551
R9964 GND.n7954 GND.n7951 0.551
R9965 GND.n7887 GND.n7886 0.551
R9966 GND.n7357 GND.n7356 0.551
R9967 GND.n6313 GND.n6312 0.551
R9968 GND.n7223 GND.n7222 0.551
R9969 GND.n11294 GND.n11293 0.551
R9970 GND.n13701 GND.n13700 0.551
R9971 GND.n8948 GND.n8947 0.551
R9972 GND.n9649 GND.n9648 0.551
R9973 GND.n15949 GND.n15948 0.551
R9974 GND.n15931 GND.n15930 0.551
R9975 GND.n16223 GND.n16220 0.551
R9976 GND.n1121 GND.n1120 0.551
R9977 GND.n9631 GND.n9630 0.551
R9978 GND.n9923 GND.n9920 0.551
R9979 GND.n1241 GND.n1240 0.551
R9980 GND.n10291 GND.n10290 0.551
R9981 GND.n10157 GND.n10156 0.551
R9982 GND.n8561 GND.n8560 0.551
R9983 GND.n8854 GND.n8853 0.551
R9984 GND.n8427 GND.n8426 0.551
R9985 GND.n10115 GND.n10114 0.551
R9986 GND.n8930 GND.n8929 0.551
R9987 GND.n9222 GND.n9219 0.551
R9988 GND.n4483 GND.n4482 0.551
R9989 GND.n4526 GND.n4525 0.551
R9990 GND.n3001 GND.n3000 0.551
R9991 GND.n3201 GND.n3200 0.551
R9992 GND.n10425 GND.n10424 0.551
R9993 GND.n15132 GND.n15131 0.551
R9994 GND.n3663 GND.n3660 0.551
R9995 GND.n3902 GND.n3901 0.551
R9996 GND.n5740 GND.n5739 0.551
R9997 GND.n10136 GND.n10134 0.549
R9998 GND.n8705 GND.n8703 0.549
R9999 GND.n15058 GND.n15057 0.536
R10000 GND.n14975 GND.n14974 0.536
R10001 GND.n14663 GND.n14662 0.536
R10002 GND.n14675 GND.n14674 0.536
R10003 GND.n14624 GND.n14623 0.536
R10004 GND.n14612 GND.n14611 0.536
R10005 GND.n15817 GND.n15816 0.536
R10006 GND.n10618 GND.n10617 0.536
R10007 GND.n10630 GND.n10629 0.536
R10008 GND.n15476 GND.n15475 0.536
R10009 GND.n14269 GND.n14268 0.536
R10010 GND.n14257 GND.n14256 0.536
R10011 GND.n14352 GND.n14351 0.536
R10012 GND.n14340 GND.n14339 0.536
R10013 GND.n2909 GND.n2908 0.536
R10014 GND.n3562 GND.n3561 0.536
R10015 GND.n4830 GND.n4829 0.536
R10016 GND.n4842 GND.n4841 0.536
R10017 GND.n5154 GND.n5153 0.536
R10018 GND.n7528 GND.n7527 0.536
R10019 GND.n12765 GND.n12764 0.536
R10020 GND.n13940 GND.n13939 0.536
R10021 GND.n13952 GND.n13951 0.536
R10022 GND.n10762 GND.n10761 0.536
R10023 GND.n10750 GND.n10749 0.536
R10024 GND.n13778 GND.n13777 0.536
R10025 GND.n13824 GND.n13823 0.536
R10026 GND.n13812 GND.n13811 0.536
R10027 GND.n11562 GND.n11561 0.536
R10028 GND.n11574 GND.n11573 0.536
R10029 GND.n11666 GND.n11665 0.536
R10030 GND.n11678 GND.n11677 0.536
R10031 GND.n11374 GND.n11373 0.536
R10032 GND.n11066 GND.n11065 0.536
R10033 GND.n11054 GND.n11053 0.536
R10034 GND.n13267 GND.n13266 0.536
R10035 GND.n8202 GND.n8201 0.536
R10036 GND.n8214 GND.n8213 0.536
R10037 GND.n8291 GND.n8290 0.536
R10038 GND.n8303 GND.n8302 0.536
R10039 GND.n6453 GND.n6452 0.536
R10040 GND.n5859 GND.n5858 0.536
R10041 GND.n5976 GND.n5975 0.536
R10042 GND.n5988 GND.n5987 0.536
R10043 GND.n6653 GND.n6652 0.536
R10044 GND.n6665 GND.n6664 0.536
R10045 GND.n6888 GND.n6887 0.536
R10046 GND.n6900 GND.n6899 0.536
R10047 GND.n6750 GND.n6749 0.536
R10048 GND.n6762 GND.n6761 0.536
R10049 GND.n7486 GND.n7485 0.536
R10050 GND.n8642 GND.n8641 0.536
R10051 GND.n9347 GND.n9346 0.536
R10052 GND.n1740 GND.n1739 0.536
R10053 GND.n1752 GND.n1751 0.536
R10054 GND.n9474 GND.n9473 0.536
R10055 GND.n9462 GND.n9461 0.536
R10056 GND.n1842 GND.n1841 0.536
R10057 GND.n1854 GND.n1853 0.536
R10058 GND.n2533 GND.n2532 0.536
R10059 GND.n2545 GND.n2544 0.536
R10060 GND.n3455 GND.n3454 0.536
R10061 GND.n3443 GND.n3442 0.536
R10062 GND.n2451 GND.n2450 0.536
R10063 GND.n2439 GND.n2438 0.536
R10064 GND.n2383 GND.n2382 0.536
R10065 GND.n2112 GND.n2111 0.536
R10066 GND.n2100 GND.n2099 0.536
R10067 GND.n2192 GND.n2191 0.536
R10068 GND.n2180 GND.n2179 0.536
R10069 GND.n15384 GND.n15383 0.536
R10070 GND.n15372 GND.n15371 0.536
R10071 GND.n15488 GND.n15487 0.536
R10072 GND.n3574 GND.n3573 0.536
R10073 GND.n13766 GND.n13765 0.536
R10074 GND.n12753 GND.n12752 0.536
R10075 GND.n13279 GND.n13278 0.536
R10076 GND.n11362 GND.n11361 0.536
R10077 GND.n6352 GND.n6351 0.536
R10078 GND.n6465 GND.n6464 0.536
R10079 GND.n7474 GND.n7473 0.536
R10080 GND.n7540 GND.n7539 0.536
R10081 GND.n9335 GND.n9334 0.536
R10082 GND.n8654 GND.n8653 0.536
R10083 GND.n2371 GND.n2370 0.536
R10084 GND.n5142 GND.n5141 0.536
R10085 GND.n2921 GND.n2920 0.536
R10086 GND.n15829 GND.n15828 0.536
R10087 GND.n14963 GND.n14962 0.536
R10088 GND.n15070 GND.n15069 0.536
R10089 GND.n14408 GND.n14407 0.506
R10090 GND.n14986 GND.n14985 0.506
R10091 GND.n14653 GND.n14651 0.506
R10092 GND.n14682 GND.n14681 0.506
R10093 GND.n14587 GND.n14585 0.506
R10094 GND.n14605 GND.n14604 0.506
R10095 GND.n15809 GND.n15808 0.506
R10096 GND.n10611 GND.n10610 0.506
R10097 GND.n10643 GND.n10642 0.506
R10098 GND.n15468 GND.n15467 0.506
R10099 GND.n14216 GND.n14214 0.506
R10100 GND.n14250 GND.n14249 0.506
R10101 GND.n14312 GND.n14310 0.506
R10102 GND.n14333 GND.n14332 0.506
R10103 GND.n2901 GND.n2900 0.506
R10104 GND.n3554 GND.n3553 0.506
R10105 GND.n4823 GND.n4822 0.506
R10106 GND.n4854 GND.n4853 0.506
R10107 GND.n5165 GND.n5164 0.506
R10108 GND.n6159 GND.n6158 0.506
R10109 GND.n12777 GND.n12776 0.506
R10110 GND.n10729 GND.n10727 0.506
R10111 GND.n13959 GND.n13958 0.506
R10112 GND.n10733 GND.n10731 0.506
R10113 GND.n10743 GND.n10742 0.506
R10114 GND.n13788 GND.n13787 0.506
R10115 GND.n13831 GND.n13830 0.506
R10116 GND.n13804 GND.n13803 0.506
R10117 GND.n11443 GND.n11441 0.506
R10118 GND.n11581 GND.n11580 0.506
R10119 GND.n11657 GND.n11655 0.506
R10120 GND.n11685 GND.n11684 0.506
R10121 GND.n11384 GND.n11383 0.506
R10122 GND.n11073 GND.n11072 0.506
R10123 GND.n11046 GND.n11045 0.506
R10124 GND.n13259 GND.n13258 0.506
R10125 GND.n8195 GND.n8194 0.506
R10126 GND.n8225 GND.n8224 0.506
R10127 GND.n8284 GND.n8283 0.506
R10128 GND.n8316 GND.n8315 0.506
R10129 GND.n6446 GND.n6445 0.506
R10130 GND.n5866 GND.n5865 0.506
R10131 GND.n5967 GND.n5965 0.506
R10132 GND.n5995 GND.n5994 0.506
R10133 GND.n6644 GND.n6642 0.506
R10134 GND.n6672 GND.n6671 0.506
R10135 GND.n6879 GND.n6877 0.506
R10136 GND.n6907 GND.n6906 0.506
R10137 GND.n6743 GND.n6742 0.506
R10138 GND.n6775 GND.n6774 0.506
R10139 GND.n7498 GND.n7497 0.506
R10140 GND.n8585 GND.n8584 0.506
R10141 GND.n9358 GND.n9357 0.506
R10142 GND.n1733 GND.n1732 0.506
R10143 GND.n1765 GND.n1764 0.506
R10144 GND.n1641 GND.n1639 0.506
R10145 GND.n9455 GND.n9454 0.506
R10146 GND.n1832 GND.n1830 0.506
R10147 GND.n1861 GND.n1860 0.506
R10148 GND.n2526 GND.n2525 0.506
R10149 GND.n2557 GND.n2556 0.506
R10150 GND.n2272 GND.n2270 0.506
R10151 GND.n3436 GND.n3435 0.506
R10152 GND.n2414 GND.n2412 0.506
R10153 GND.n2432 GND.n2431 0.506
R10154 GND.n2294 GND.n2293 0.506
R10155 GND.n2059 GND.n2057 0.506
R10156 GND.n2093 GND.n2092 0.506
R10157 GND.n2155 GND.n2153 0.506
R10158 GND.n2173 GND.n2172 0.506
R10159 GND.n15391 GND.n15390 0.506
R10160 GND.n15364 GND.n15363 0.506
R10161 GND.n16450 GND.n16449 0.506
R10162 GND.n16564 GND.n16563 0.506
R10163 GND.n16390 GND.n16389 0.506
R10164 GND.n16711 GND.n16710 0.506
R10165 GND.n16825 GND.n16824 0.506
R10166 GND.n16651 GND.n16650 0.506
R10167 GND.n16972 GND.n16971 0.506
R10168 GND.n17086 GND.n17085 0.506
R10169 GND.n16912 GND.n16911 0.506
R10170 GND.n17233 GND.n17232 0.506
R10171 GND.n17347 GND.n17346 0.506
R10172 GND.n17173 GND.n17172 0.506
R10173 GND.n17494 GND.n17493 0.506
R10174 GND.n17608 GND.n17607 0.506
R10175 GND.n17434 GND.n17433 0.506
R10176 GND.n677 GND.n676 0.506
R10177 GND.n780 GND.n779 0.506
R10178 GND.n611 GND.n610 0.506
R10179 GND.n419 GND.n418 0.506
R10180 GND.n522 GND.n521 0.506
R10181 GND.n353 GND.n352 0.506
R10182 GND.n161 GND.n160 0.506
R10183 GND.n264 GND.n263 0.506
R10184 GND.n95 GND.n94 0.506
R10185 GND.n17776 GND.n17775 0.506
R10186 GND.n17853 GND.n17852 0.506
R10187 GND.n17931 GND.n17930 0.506
R10188 GND.n15495 GND.n15494 0.506
R10189 GND.n3581 GND.n3580 0.506
R10190 GND.n13759 GND.n13758 0.506
R10191 GND.n12746 GND.n12745 0.506
R10192 GND.n13286 GND.n13285 0.506
R10193 GND.n11355 GND.n11354 0.506
R10194 GND.n6365 GND.n6363 0.506
R10195 GND.n6342 GND.n6341 0.506
R10196 GND.n7467 GND.n7466 0.506
R10197 GND.n7547 GND.n7546 0.506
R10198 GND.n9328 GND.n9327 0.506
R10199 GND.n8661 GND.n8660 0.506
R10200 GND.n2364 GND.n2363 0.506
R10201 GND.n5135 GND.n5134 0.506
R10202 GND.n2928 GND.n2927 0.506
R10203 GND.n15836 GND.n15835 0.506
R10204 GND.n14956 GND.n14955 0.506
R10205 GND.n15077 GND.n15076 0.506
R10206 GND.n15041 GND.n15040 0.476
R10207 GND.n14426 GND.n14425 0.476
R10208 GND.n14639 GND.n14638 0.476
R10209 GND.n14689 GND.n14688 0.476
R10210 GND.n14573 GND.n14572 0.476
R10211 GND.n14598 GND.n14597 0.476
R10212 GND.n15795 GND.n15794 0.476
R10213 GND.n10604 GND.n10603 0.476
R10214 GND.n10655 GND.n10654 0.476
R10215 GND.n14069 GND.n14068 0.476
R10216 GND.n14288 GND.n14287 0.476
R10217 GND.n14243 GND.n14242 0.476
R10218 GND.n14295 GND.n14294 0.476
R10219 GND.n14326 GND.n14325 0.476
R10220 GND.n2887 GND.n2886 0.476
R10221 GND.n3541 GND.n3540 0.476
R10222 GND.n4816 GND.n4815 0.476
R10223 GND.n4866 GND.n4865 0.476
R10224 GND.n5177 GND.n5176 0.476
R10225 GND.n6946 GND.n6945 0.476
R10226 GND.n12789 GND.n12788 0.476
R10227 GND.n13921 GND.n13920 0.476
R10228 GND.n13966 GND.n13965 0.476
R10229 GND.n10822 GND.n10821 0.476
R10230 GND.n10736 GND.n10735 0.476
R10231 GND.n10990 GND.n10989 0.476
R10232 GND.n13838 GND.n13837 0.476
R10233 GND.n10941 GND.n10940 0.476
R10234 GND.n11543 GND.n11542 0.476
R10235 GND.n11588 GND.n11587 0.476
R10236 GND.n11483 GND.n11482 0.476
R10237 GND.n11692 GND.n11691 0.476
R10238 GND.n11396 GND.n11395 0.476
R10239 GND.n11080 GND.n11079 0.476
R10240 GND.n11020 GND.n11019 0.476
R10241 GND.n13245 GND.n13244 0.476
R10242 GND.n8188 GND.n8187 0.476
R10243 GND.n6067 GND.n6066 0.476
R10244 GND.n8277 GND.n8276 0.476
R10245 GND.n8328 GND.n8327 0.476
R10246 GND.n6439 GND.n6438 0.476
R10247 GND.n5873 GND.n5872 0.476
R10248 GND.n5952 GND.n5951 0.476
R10249 GND.n6002 GND.n6001 0.476
R10250 GND.n6630 GND.n6629 0.476
R10251 GND.n6679 GND.n6678 0.476
R10252 GND.n6865 GND.n6864 0.476
R10253 GND.n6914 GND.n6913 0.476
R10254 GND.n6736 GND.n6735 0.476
R10255 GND.n6787 GND.n6786 0.476
R10256 GND.n6537 GND.n6536 0.476
R10257 GND.n8625 GND.n8624 0.476
R10258 GND.n9370 GND.n9369 0.476
R10259 GND.n1726 GND.n1725 0.476
R10260 GND.n1777 GND.n1776 0.476
R10261 GND.n9493 GND.n9492 0.476
R10262 GND.n9448 GND.n9447 0.476
R10263 GND.n1818 GND.n1817 0.476
R10264 GND.n1868 GND.n1867 0.476
R10265 GND.n2519 GND.n2518 0.476
R10266 GND.n2569 GND.n2568 0.476
R10267 GND.n3474 GND.n3473 0.476
R10268 GND.n3429 GND.n3428 0.476
R10269 GND.n2396 GND.n2395 0.476
R10270 GND.n2425 GND.n2424 0.476
R10271 GND.n2283 GND.n2282 0.476
R10272 GND.n2131 GND.n2130 0.476
R10273 GND.n2086 GND.n2085 0.476
R10274 GND.n2138 GND.n2137 0.476
R10275 GND.n2166 GND.n2165 0.476
R10276 GND.n15398 GND.n15397 0.476
R10277 GND.n15349 GND.n15348 0.476
R10278 GND.n16462 GND.n16461 0.476
R10279 GND.n16545 GND.n16544 0.476
R10280 GND.n16370 GND.n16369 0.476
R10281 GND.n16723 GND.n16722 0.476
R10282 GND.n16806 GND.n16805 0.476
R10283 GND.n16631 GND.n16630 0.476
R10284 GND.n16984 GND.n16983 0.476
R10285 GND.n17067 GND.n17066 0.476
R10286 GND.n16892 GND.n16891 0.476
R10287 GND.n17245 GND.n17244 0.476
R10288 GND.n17328 GND.n17327 0.476
R10289 GND.n17153 GND.n17152 0.476
R10290 GND.n17506 GND.n17505 0.476
R10291 GND.n17589 GND.n17588 0.476
R10292 GND.n17414 GND.n17413 0.476
R10293 GND.n658 GND.n657 0.476
R10294 GND.n761 GND.n760 0.476
R10295 GND.n593 GND.n592 0.476
R10296 GND.n400 GND.n399 0.476
R10297 GND.n503 GND.n502 0.476
R10298 GND.n335 GND.n334 0.476
R10299 GND.n142 GND.n141 0.476
R10300 GND.n245 GND.n244 0.476
R10301 GND.n77 GND.n76 0.476
R10302 GND.n17757 GND.n17756 0.476
R10303 GND.n17834 GND.n17833 0.476
R10304 GND.n17913 GND.n17912 0.476
R10305 GND.n15502 GND.n15501 0.475
R10306 GND.n3588 GND.n3587 0.475
R10307 GND.n13752 GND.n13751 0.475
R10308 GND.n12739 GND.n12738 0.475
R10309 GND.n13293 GND.n13292 0.475
R10310 GND.n11348 GND.n11347 0.475
R10311 GND.n6373 GND.n6372 0.475
R10312 GND.n6482 GND.n6481 0.475
R10313 GND.n7460 GND.n7459 0.475
R10314 GND.n7554 GND.n7553 0.475
R10315 GND.n9321 GND.n9320 0.475
R10316 GND.n8668 GND.n8667 0.475
R10317 GND.n2357 GND.n2356 0.475
R10318 GND.n5128 GND.n5127 0.475
R10319 GND.n2935 GND.n2934 0.475
R10320 GND.n15843 GND.n15842 0.475
R10321 GND.n14949 GND.n14948 0.475
R10322 GND.n15084 GND.n15083 0.475
R10323 GND.n7018 GND.n7017 0.455
R10324 GND.n8118 GND.n8117 0.455
R10325 GND.n13368 GND.n13367 0.455
R10326 GND.n12670 GND.n12669 0.455
R10327 GND.n12561 GND.n12560 0.455
R10328 GND.n13477 GND.n13476 0.455
R10329 GND.n12875 GND.n12872 0.455
R10330 GND.n11766 GND.n11763 0.455
R10331 GND.n12432 GND.n12429 0.455
R10332 GND.n12387 GND.n12386 0.455
R10333 GND.n13110 GND.n13109 0.455
R10334 GND.n12942 GND.n12941 0.455
R10335 GND.n7708 GND.n7707 0.455
R10336 GND.n7911 GND.n7908 0.455
R10337 GND.n8009 GND.n8008 0.455
R10338 GND.n7127 GND.n7126 0.455
R10339 GND.n6301 GND.n6300 0.455
R10340 GND.n11282 GND.n11281 0.455
R10341 GND.n13689 GND.n13688 0.455
R10342 GND.n14882 GND.n14881 0.455
R10343 GND.n16197 GND.n16194 0.455
R10344 GND.n860 GND.n857 0.455
R10345 GND.n909 GND.n908 0.455
R10346 GND.n1109 GND.n1108 0.455
R10347 GND.n9897 GND.n9894 0.455
R10348 GND.n1498 GND.n1495 0.455
R10349 GND.n1453 GND.n1452 0.455
R10350 GND.n1253 GND.n1252 0.455
R10351 GND.n8842 GND.n8841 0.455
R10352 GND.n10103 GND.n10102 0.455
R10353 GND.n9196 GND.n9193 0.455
R10354 GND.n5479 GND.n5476 0.455
R10355 GND.n4220 GND.n4217 0.455
R10356 GND.n4269 GND.n4268 0.455
R10357 GND.n15580 GND.n15579 0.455
R10358 GND.n4720 GND.n4719 0.455
R10359 GND.n5066 GND.n5065 0.455
R10360 GND.n4957 GND.n4956 0.455
R10361 GND.n4611 GND.n4610 0.455
R10362 GND.n3013 GND.n3012 0.455
R10363 GND.n3213 GND.n3212 0.455
R10364 GND.n14773 GND.n14772 0.455
R10365 GND.n10437 GND.n10436 0.455
R10366 GND.n15689 GND.n15688 0.455
R10367 GND.n15144 GND.n15143 0.455
R10368 GND.n3637 GND.n3634 0.455
R10369 GND.n3890 GND.n3889 0.455
R10370 GND.n5528 GND.n5527 0.455
R10371 GND.n5728 GND.n5727 0.455
R10372 GND.n15031 GND.n15030 0.445
R10373 GND.n14436 GND.n14435 0.445
R10374 GND.n14510 GND.n14509 0.445
R10375 GND.n14696 GND.n14695 0.445
R10376 GND.n14562 GND.n14561 0.445
R10377 GND.n14381 GND.n14380 0.445
R10378 GND.n15785 GND.n15784 0.445
R10379 GND.n10597 GND.n10596 0.445
R10380 GND.n10665 GND.n10664 0.445
R10381 GND.n14059 GND.n14058 0.445
R10382 GND.n14204 GND.n14203 0.445
R10383 GND.n14236 GND.n14235 0.445
R10384 GND.n14151 GND.n14150 0.445
R10385 GND.n14319 GND.n14318 0.445
R10386 GND.n4809 GND.n4808 0.445
R10387 GND.n4876 GND.n4875 0.445
R10388 GND.n5187 GND.n5186 0.445
R10389 GND.n6956 GND.n6955 0.445
R10390 GND.n12799 GND.n12798 0.445
R10391 GND.n13911 GND.n13910 0.445
R10392 GND.n13973 GND.n13972 0.445
R10393 GND.n10812 GND.n10811 0.445
R10394 GND.n10854 GND.n10853 0.445
R10395 GND.n10980 GND.n10979 0.445
R10396 GND.n13845 GND.n13844 0.445
R10397 GND.n10931 GND.n10930 0.445
R10398 GND.n11533 GND.n11532 0.445
R10399 GND.n11595 GND.n11594 0.445
R10400 GND.n11473 GND.n11472 0.445
R10401 GND.n11699 GND.n11698 0.445
R10402 GND.n11406 GND.n11405 0.445
R10403 GND.n11087 GND.n11086 0.445
R10404 GND.n11624 GND.n11623 0.445
R10405 GND.n13235 GND.n13234 0.445
R10406 GND.n8181 GND.n8180 0.445
R10407 GND.n6077 GND.n6076 0.445
R10408 GND.n8270 GND.n8269 0.445
R10409 GND.n8338 GND.n8337 0.445
R10410 GND.n6432 GND.n6431 0.445
R10411 GND.n5880 GND.n5879 0.445
R10412 GND.n5942 GND.n5941 0.445
R10413 GND.n6009 GND.n6008 0.445
R10414 GND.n6620 GND.n6619 0.445
R10415 GND.n6686 GND.n6685 0.445
R10416 GND.n6855 GND.n6854 0.445
R10417 GND.n6921 GND.n6920 0.445
R10418 GND.n6729 GND.n6728 0.445
R10419 GND.n6797 GND.n6796 0.445
R10420 GND.n6547 GND.n6546 0.445
R10421 GND.n8615 GND.n8614 0.445
R10422 GND.n9380 GND.n9379 0.445
R10423 GND.n1719 GND.n1718 0.445
R10424 GND.n1787 GND.n1786 0.445
R10425 GND.n1651 GND.n1650 0.445
R10426 GND.n9441 GND.n9440 0.445
R10427 GND.n1626 GND.n1625 0.445
R10428 GND.n1875 GND.n1874 0.445
R10429 GND.n2512 GND.n2511 0.445
R10430 GND.n2579 GND.n2578 0.445
R10431 GND.n2259 GND.n2258 0.445
R10432 GND.n3422 GND.n3421 0.445
R10433 GND.n2230 GND.n2229 0.445
R10434 GND.n2610 GND.n2609 0.445
R10435 GND.n2317 GND.n2316 0.445
R10436 GND.n2046 GND.n2045 0.445
R10437 GND.n2079 GND.n2078 0.445
R10438 GND.n1993 GND.n1992 0.445
R10439 GND.n2637 GND.n2636 0.445
R10440 GND.n15405 GND.n15404 0.445
R10441 GND.n15339 GND.n15338 0.445
R10442 GND.n16474 GND.n16473 0.445
R10443 GND.n16534 GND.n16533 0.445
R10444 GND.n16359 GND.n16358 0.445
R10445 GND.n16735 GND.n16734 0.445
R10446 GND.n16795 GND.n16794 0.445
R10447 GND.n16620 GND.n16619 0.445
R10448 GND.n16996 GND.n16995 0.445
R10449 GND.n17056 GND.n17055 0.445
R10450 GND.n16881 GND.n16880 0.445
R10451 GND.n17257 GND.n17256 0.445
R10452 GND.n17317 GND.n17316 0.445
R10453 GND.n17142 GND.n17141 0.445
R10454 GND.n17518 GND.n17517 0.445
R10455 GND.n17578 GND.n17577 0.445
R10456 GND.n17403 GND.n17402 0.445
R10457 GND.n647 GND.n646 0.445
R10458 GND.n749 GND.n748 0.445
R10459 GND.n581 GND.n580 0.445
R10460 GND.n389 GND.n388 0.445
R10461 GND.n491 GND.n490 0.445
R10462 GND.n323 GND.n322 0.445
R10463 GND.n131 GND.n130 0.445
R10464 GND.n233 GND.n232 0.445
R10465 GND.n65 GND.n64 0.445
R10466 GND.n17746 GND.n17745 0.445
R10467 GND.n17822 GND.n17821 0.445
R10468 GND.n17901 GND.n17900 0.445
R10469 GND.n15509 GND.n15508 0.445
R10470 GND.n3531 GND.n3530 0.445
R10471 GND.n3595 GND.n3594 0.445
R10472 GND.n13745 GND.n13744 0.445
R10473 GND.n12732 GND.n12731 0.445
R10474 GND.n13300 GND.n13299 0.445
R10475 GND.n11341 GND.n11340 0.445
R10476 GND.n6388 GND.n6387 0.445
R10477 GND.n6491 GND.n6490 0.445
R10478 GND.n7453 GND.n7452 0.445
R10479 GND.n7561 GND.n7560 0.445
R10480 GND.n9314 GND.n9313 0.445
R10481 GND.n8675 GND.n8674 0.445
R10482 GND.n2350 GND.n2349 0.445
R10483 GND.n5121 GND.n5120 0.445
R10484 GND.n2877 GND.n2876 0.445
R10485 GND.n2942 GND.n2941 0.445
R10486 GND.n15850 GND.n15849 0.445
R10487 GND.n14942 GND.n14941 0.445
R10488 GND.n15091 GND.n15090 0.445
R10489 GND.n15022 GND.n15021 0.414
R10490 GND.n14446 GND.n14445 0.414
R10491 GND.n14520 GND.n14519 0.414
R10492 GND.n14703 GND.n14702 0.414
R10493 GND.n14551 GND.n14550 0.414
R10494 GND.n14388 GND.n14387 0.414
R10495 GND.n15776 GND.n15775 0.414
R10496 GND.n10590 GND.n10589 0.414
R10497 GND.n10675 GND.n10674 0.414
R10498 GND.n14050 GND.n14049 0.414
R10499 GND.n14193 GND.n14192 0.414
R10500 GND.n14229 GND.n14228 0.414
R10501 GND.n14140 GND.n14139 0.414
R10502 GND.n10700 GND.n10699 0.414
R10503 GND.n2867 GND.n2866 0.414
R10504 GND.n3521 GND.n3520 0.414
R10505 GND.n4802 GND.n4801 0.414
R10506 GND.n4886 GND.n4885 0.414
R10507 GND.n5197 GND.n5196 0.414
R10508 GND.n6966 GND.n6965 0.414
R10509 GND.n12809 GND.n12808 0.414
R10510 GND.n13901 GND.n13900 0.414
R10511 GND.n13980 GND.n13979 0.414
R10512 GND.n10802 GND.n10801 0.414
R10513 GND.n10861 GND.n10860 0.414
R10514 GND.n10971 GND.n10970 0.414
R10515 GND.n13852 GND.n13851 0.414
R10516 GND.n10922 GND.n10921 0.414
R10517 GND.n11523 GND.n11522 0.414
R10518 GND.n11602 GND.n11601 0.414
R10519 GND.n11463 GND.n11462 0.414
R10520 GND.n11706 GND.n11705 0.414
R10521 GND.n11416 GND.n11415 0.414
R10522 GND.n11094 GND.n11093 0.414
R10523 GND.n11634 GND.n11633 0.414
R10524 GND.n13226 GND.n13225 0.414
R10525 GND.n8174 GND.n8173 0.414
R10526 GND.n6087 GND.n6086 0.414
R10527 GND.n8263 GND.n8262 0.414
R10528 GND.n8348 GND.n8347 0.414
R10529 GND.n6425 GND.n6424 0.414
R10530 GND.n5887 GND.n5886 0.414
R10531 GND.n5932 GND.n5931 0.414
R10532 GND.n6016 GND.n6015 0.414
R10533 GND.n6610 GND.n6609 0.414
R10534 GND.n6693 GND.n6692 0.414
R10535 GND.n6845 GND.n6844 0.414
R10536 GND.n6928 GND.n6927 0.414
R10537 GND.n6722 GND.n6721 0.414
R10538 GND.n6807 GND.n6806 0.414
R10539 GND.n6557 GND.n6556 0.414
R10540 GND.n8605 GND.n8604 0.414
R10541 GND.n9390 GND.n9389 0.414
R10542 GND.n1712 GND.n1711 0.414
R10543 GND.n1797 GND.n1796 0.414
R10544 GND.n1661 GND.n1660 0.414
R10545 GND.n9434 GND.n9433 0.414
R10546 GND.n1615 GND.n1614 0.414
R10547 GND.n1882 GND.n1881 0.414
R10548 GND.n2505 GND.n2504 0.414
R10549 GND.n2589 GND.n2588 0.414
R10550 GND.n2248 GND.n2247 0.414
R10551 GND.n3415 GND.n3414 0.414
R10552 GND.n2219 GND.n2218 0.414
R10553 GND.n2617 GND.n2616 0.414
R10554 GND.n2327 GND.n2326 0.414
R10555 GND.n2035 GND.n2034 0.414
R10556 GND.n2072 GND.n2071 0.414
R10557 GND.n1982 GND.n1981 0.414
R10558 GND.n2644 GND.n2643 0.414
R10559 GND.n15412 GND.n15411 0.414
R10560 GND.n15330 GND.n15329 0.414
R10561 GND.n16439 GND.n16438 0.414
R10562 GND.n16525 GND.n16524 0.414
R10563 GND.n16348 GND.n16347 0.414
R10564 GND.n16700 GND.n16699 0.414
R10565 GND.n16786 GND.n16785 0.414
R10566 GND.n16609 GND.n16608 0.414
R10567 GND.n16961 GND.n16960 0.414
R10568 GND.n17047 GND.n17046 0.414
R10569 GND.n16870 GND.n16869 0.414
R10570 GND.n17222 GND.n17221 0.414
R10571 GND.n17308 GND.n17307 0.414
R10572 GND.n17131 GND.n17130 0.414
R10573 GND.n17483 GND.n17482 0.414
R10574 GND.n17569 GND.n17568 0.414
R10575 GND.n17392 GND.n17391 0.414
R10576 GND.n635 GND.n634 0.414
R10577 GND.n737 GND.n736 0.414
R10578 GND.n569 GND.n568 0.414
R10579 GND.n377 GND.n376 0.414
R10580 GND.n479 GND.n478 0.414
R10581 GND.n311 GND.n310 0.414
R10582 GND.n119 GND.n118 0.414
R10583 GND.n221 GND.n220 0.414
R10584 GND.n53 GND.n52 0.414
R10585 GND.n17734 GND.n17733 0.414
R10586 GND.n17810 GND.n17809 0.414
R10587 GND.n17889 GND.n17888 0.414
R10588 GND.n15516 GND.n15515 0.413
R10589 GND.n3602 GND.n3601 0.413
R10590 GND.n13738 GND.n13737 0.413
R10591 GND.n12725 GND.n12724 0.413
R10592 GND.n13307 GND.n13306 0.413
R10593 GND.n11334 GND.n11333 0.413
R10594 GND.n6397 GND.n6396 0.413
R10595 GND.n6500 GND.n6499 0.413
R10596 GND.n7446 GND.n7445 0.413
R10597 GND.n7568 GND.n7567 0.413
R10598 GND.n9307 GND.n9306 0.413
R10599 GND.n8682 GND.n8681 0.413
R10600 GND.n2343 GND.n2342 0.413
R10601 GND.n5114 GND.n5113 0.413
R10602 GND.n2949 GND.n2948 0.413
R10603 GND.n15857 GND.n15856 0.413
R10604 GND.n14935 GND.n14934 0.413
R10605 GND.n15098 GND.n15097 0.413
R10606 GND.n15014 GND.n15013 0.382
R10607 GND.n14455 GND.n14454 0.382
R10608 GND.n14501 GND.n14500 0.382
R10609 GND.n14710 GND.n14709 0.382
R10610 GND.n14540 GND.n14539 0.382
R10611 GND.n14395 GND.n14394 0.382
R10612 GND.n15768 GND.n15767 0.382
R10613 GND.n10583 GND.n10582 0.382
R10614 GND.n10684 GND.n10683 0.382
R10615 GND.n14042 GND.n14041 0.382
R10616 GND.n14172 GND.n14171 0.382
R10617 GND.n14222 GND.n14221 0.382
R10618 GND.n14130 GND.n14129 0.382
R10619 GND.n10707 GND.n10706 0.382
R10620 GND.n4795 GND.n4794 0.382
R10621 GND.n4895 GND.n4894 0.382
R10622 GND.n5206 GND.n5205 0.382
R10623 GND.n6975 GND.n6974 0.382
R10624 GND.n12818 GND.n12817 0.382
R10625 GND.n13893 GND.n13892 0.382
R10626 GND.n13987 GND.n13986 0.382
R10627 GND.n10793 GND.n10792 0.382
R10628 GND.n10868 GND.n10867 0.382
R10629 GND.n10963 GND.n10962 0.382
R10630 GND.n13859 GND.n13858 0.382
R10631 GND.n10914 GND.n10913 0.382
R10632 GND.n11515 GND.n11514 0.382
R10633 GND.n11609 GND.n11608 0.382
R10634 GND.n11454 GND.n11453 0.382
R10635 GND.n11713 GND.n11712 0.382
R10636 GND.n11425 GND.n11424 0.382
R10637 GND.n11101 GND.n11100 0.382
R10638 GND.n11643 GND.n11642 0.382
R10639 GND.n13218 GND.n13217 0.382
R10640 GND.n8167 GND.n8166 0.382
R10641 GND.n6096 GND.n6095 0.382
R10642 GND.n8256 GND.n8255 0.382
R10643 GND.n8357 GND.n8356 0.382
R10644 GND.n6418 GND.n6417 0.382
R10645 GND.n5894 GND.n5893 0.382
R10646 GND.n5923 GND.n5922 0.382
R10647 GND.n6023 GND.n6022 0.382
R10648 GND.n6601 GND.n6600 0.382
R10649 GND.n6700 GND.n6699 0.382
R10650 GND.n6836 GND.n6835 0.382
R10651 GND.n6935 GND.n6934 0.382
R10652 GND.n6715 GND.n6714 0.382
R10653 GND.n6816 GND.n6815 0.382
R10654 GND.n6566 GND.n6565 0.382
R10655 GND.n8597 GND.n8596 0.382
R10656 GND.n9399 GND.n9398 0.382
R10657 GND.n1705 GND.n1704 0.382
R10658 GND.n1806 GND.n1805 0.382
R10659 GND.n1671 GND.n1670 0.382
R10660 GND.n9427 GND.n9426 0.382
R10661 GND.n1593 GND.n1592 0.382
R10662 GND.n1889 GND.n1888 0.382
R10663 GND.n2498 GND.n2497 0.382
R10664 GND.n2598 GND.n2597 0.382
R10665 GND.n2464 GND.n2463 0.382
R10666 GND.n3408 GND.n3407 0.382
R10667 GND.n2208 GND.n2207 0.382
R10668 GND.n2624 GND.n2623 0.382
R10669 GND.n2308 GND.n2307 0.382
R10670 GND.n2014 GND.n2013 0.382
R10671 GND.n2065 GND.n2064 0.382
R10672 GND.n1971 GND.n1970 0.382
R10673 GND.n2651 GND.n2650 0.382
R10674 GND.n15419 GND.n15418 0.382
R10675 GND.n15322 GND.n15321 0.382
R10676 GND.n16428 GND.n16427 0.382
R10677 GND.n16499 GND.n16498 0.382
R10678 GND.n16337 GND.n16336 0.382
R10679 GND.n16689 GND.n16688 0.382
R10680 GND.n16760 GND.n16759 0.382
R10681 GND.n16598 GND.n16597 0.382
R10682 GND.n16950 GND.n16949 0.382
R10683 GND.n17021 GND.n17020 0.382
R10684 GND.n16859 GND.n16858 0.382
R10685 GND.n17211 GND.n17210 0.382
R10686 GND.n17282 GND.n17281 0.382
R10687 GND.n17120 GND.n17119 0.382
R10688 GND.n17472 GND.n17471 0.382
R10689 GND.n17543 GND.n17542 0.382
R10690 GND.n17381 GND.n17380 0.382
R10691 GND.n693 GND.n692 0.382
R10692 GND.n720 GND.n719 0.382
R10693 GND.n560 GND.n559 0.382
R10694 GND.n435 GND.n434 0.382
R10695 GND.n462 GND.n461 0.382
R10696 GND.n302 GND.n301 0.382
R10697 GND.n177 GND.n176 0.382
R10698 GND.n204 GND.n203 0.382
R10699 GND.n44 GND.n43 0.382
R10700 GND.n17792 GND.n17791 0.382
R10701 GND.n17714 GND.n17713 0.382
R10702 GND.n17880 GND.n17879 0.382
R10703 GND.n15523 GND.n15522 0.382
R10704 GND.n3513 GND.n3512 0.382
R10705 GND.n3609 GND.n3608 0.382
R10706 GND.n13731 GND.n13730 0.382
R10707 GND.n12718 GND.n12717 0.382
R10708 GND.n13314 GND.n13313 0.382
R10709 GND.n11327 GND.n11326 0.382
R10710 GND.n5839 GND.n5838 0.382
R10711 GND.n6508 GND.n6507 0.382
R10712 GND.n7439 GND.n7438 0.382
R10713 GND.n7575 GND.n7574 0.382
R10714 GND.n9300 GND.n9299 0.382
R10715 GND.n8689 GND.n8688 0.382
R10716 GND.n2336 GND.n2335 0.382
R10717 GND.n5107 GND.n5106 0.382
R10718 GND.n2859 GND.n2858 0.382
R10719 GND.n2956 GND.n2955 0.382
R10720 GND.n15864 GND.n15863 0.382
R10721 GND.n14928 GND.n14927 0.382
R10722 GND.n15105 GND.n15104 0.382
R10723 GND.n15631 GND.n15626 0.376
R10724 GND.n15640 GND.n15634 0.376
R10725 GND.n11235 GND.n11230 0.376
R10726 GND.n11227 GND.n11222 0.376
R10727 GND.n13642 GND.n13637 0.376
R10728 GND.n13634 GND.n13629 0.376
R10729 GND.n13419 GND.n13414 0.376
R10730 GND.n13428 GND.n13422 0.376
R10731 GND.n12621 GND.n12616 0.376
R10732 GND.n12613 GND.n12607 0.376
R10733 GND.n13067 GND.n13066 0.376
R10734 GND.n13066 GND.n13065 0.376
R10735 GND.n13144 GND.n13142 0.376
R10736 GND.n13144 GND.n13143 0.376
R10737 GND.n12905 GND.n12902 0.376
R10738 GND.n12905 GND.n12904 0.376
R10739 GND.n11732 GND.n11731 0.376
R10740 GND.n11733 GND.n11732 0.376
R10741 GND.n11961 GND.n11960 0.376
R10742 GND.n11960 GND.n11959 0.376
R10743 GND.n12040 GND.n12038 0.376
R10744 GND.n12040 GND.n12039 0.376
R10745 GND.n11778 GND.n11775 0.376
R10746 GND.n11778 GND.n11777 0.376
R10747 GND.n11747 GND.n11746 0.376
R10748 GND.n11748 GND.n11747 0.376
R10749 GND.n12254 GND.n12253 0.376
R10750 GND.n12253 GND.n12252 0.376
R10751 GND.n12144 GND.n12142 0.376
R10752 GND.n12144 GND.n12143 0.376
R10753 GND.n12462 GND.n12459 0.376
R10754 GND.n12462 GND.n12461 0.376
R10755 GND.n11738 GND.n11737 0.376
R10756 GND.n11739 GND.n11738 0.376
R10757 GND.n7742 GND.n7741 0.376
R10758 GND.n7741 GND.n7740 0.376
R10759 GND.n7639 GND.n7637 0.376
R10760 GND.n7639 GND.n7638 0.376
R10761 GND.n7923 GND.n7920 0.376
R10762 GND.n7923 GND.n7922 0.376
R10763 GND.n6146 GND.n6145 0.376
R10764 GND.n6147 GND.n6146 0.376
R10765 GND.n7296 GND.n7290 0.376
R10766 GND.n7287 GND.n7281 0.376
R10767 GND.n6254 GND.n6249 0.376
R10768 GND.n6246 GND.n6241 0.376
R10769 GND.n7069 GND.n7064 0.376
R10770 GND.n7078 GND.n7072 0.376
R10771 GND.n8069 GND.n8063 0.376
R10772 GND.n8060 GND.n8055 0.376
R10773 GND.n15997 GND.n15996 0.376
R10774 GND.n15996 GND.n15995 0.376
R10775 GND.n16012 GND.n16011 0.376
R10776 GND.n16105 GND.n16100 0.376
R10777 GND.n16113 GND.n16108 0.376
R10778 GND.n1066 GND.n1065 0.376
R10779 GND.n1065 GND.n1064 0.376
R10780 GND.n1058 GND.n1057 0.376
R10781 GND.n969 GND.n964 0.376
R10782 GND.n961 GND.n955 0.376
R10783 GND.n9697 GND.n9696 0.376
R10784 GND.n9696 GND.n9695 0.376
R10785 GND.n9712 GND.n9711 0.376
R10786 GND.n9805 GND.n9800 0.376
R10787 GND.n9813 GND.n9808 0.376
R10788 GND.n1287 GND.n1286 0.376
R10789 GND.n1286 GND.n1285 0.376
R10790 GND.n1302 GND.n1301 0.376
R10791 GND.n1395 GND.n1390 0.376
R10792 GND.n1404 GND.n1398 0.376
R10793 GND.n10230 GND.n10224 0.376
R10794 GND.n10221 GND.n10215 0.376
R10795 GND.n10056 GND.n10051 0.376
R10796 GND.n10048 GND.n10043 0.376
R10797 GND.n8795 GND.n8790 0.376
R10798 GND.n8787 GND.n8782 0.376
R10799 GND.n8500 GND.n8494 0.376
R10800 GND.n8491 GND.n8485 0.376
R10801 GND.n8996 GND.n8995 0.376
R10802 GND.n8995 GND.n8994 0.376
R10803 GND.n9011 GND.n9010 0.376
R10804 GND.n9104 GND.n9099 0.376
R10805 GND.n9112 GND.n9107 0.376
R10806 GND.n5685 GND.n5684 0.376
R10807 GND.n5684 GND.n5683 0.376
R10808 GND.n5677 GND.n5676 0.376
R10809 GND.n5588 GND.n5583 0.376
R10810 GND.n5580 GND.n5574 0.376
R10811 GND.n4426 GND.n4425 0.376
R10812 GND.n4425 GND.n4424 0.376
R10813 GND.n4418 GND.n4417 0.376
R10814 GND.n4329 GND.n4324 0.376
R10815 GND.n4321 GND.n4315 0.376
R10816 GND.n4671 GND.n4666 0.376
R10817 GND.n4663 GND.n4657 0.376
R10818 GND.n5017 GND.n5012 0.376
R10819 GND.n5009 GND.n5003 0.376
R10820 GND.n3062 GND.n3057 0.376
R10821 GND.n3070 GND.n3065 0.376
R10822 GND.n3262 GND.n3257 0.376
R10823 GND.n3270 GND.n3265 0.376
R10824 GND.n8881 GND.n8880 0.376
R10825 GND.n10486 GND.n10481 0.376
R10826 GND.n10494 GND.n10489 0.376
R10827 GND.n14833 GND.n14828 0.376
R10828 GND.n14825 GND.n14819 0.376
R10829 GND.n15193 GND.n15188 0.376
R10830 GND.n15201 GND.n15196 0.376
R10831 GND.n3847 GND.n3846 0.376
R10832 GND.n3846 GND.n3845 0.376
R10833 GND.n3839 GND.n3838 0.376
R10834 GND.n3750 GND.n3745 0.376
R10835 GND.n3742 GND.n3737 0.376
R10836 GND.n15718 GND.n15717 0.359
R10837 GND.n15122 GND.n15113 0.359
R10838 GND.n11993 GND.n11992 0.358
R10839 GND.n12065 GND.n12064 0.358
R10840 GND.n11802 GND.n11799 0.358
R10841 GND.n12231 GND.n12230 0.358
R10842 GND.n12169 GND.n12168 0.358
R10843 GND.n13098 GND.n13097 0.358
R10844 GND.n7720 GND.n7719 0.358
R10845 GND.n7947 GND.n7944 0.358
R10846 GND.n7332 GND.n7331 0.358
R10847 GND.n6289 GND.n6288 0.358
R10848 GND.n7248 GND.n7247 0.358
R10849 GND.n11270 GND.n11269 0.358
R10850 GND.n13677 GND.n13676 0.358
R10851 GND.n8973 GND.n8972 0.358
R10852 GND.n9674 GND.n9673 0.358
R10853 GND.n15974 GND.n15973 0.358
R10854 GND.n15922 GND.n15921 0.358
R10855 GND.n16216 GND.n16213 0.358
R10856 GND.n1097 GND.n1096 0.358
R10857 GND.n9622 GND.n9621 0.358
R10858 GND.n9916 GND.n9913 0.358
R10859 GND.n1265 GND.n1264 0.358
R10860 GND.n10266 GND.n10265 0.358
R10861 GND.n10182 GND.n10181 0.358
R10862 GND.n8536 GND.n8535 0.358
R10863 GND.n8830 GND.n8829 0.358
R10864 GND.n8452 GND.n8451 0.358
R10865 GND.n10091 GND.n10090 0.358
R10866 GND.n8921 GND.n8920 0.358
R10867 GND.n9215 GND.n9212 0.358
R10868 GND.n4458 GND.n4457 0.358
R10869 GND.n4517 GND.n4516 0.358
R10870 GND.n3025 GND.n3024 0.358
R10871 GND.n3225 GND.n3224 0.358
R10872 GND.n10449 GND.n10448 0.358
R10873 GND.n15156 GND.n15155 0.358
R10874 GND.n3656 GND.n3653 0.358
R10875 GND.n3878 GND.n3877 0.358
R10876 GND.n5716 GND.n5715 0.358
R10877 GND.n12115 GND.n12096 0.329
R10878 GND.n12495 GND.n11735 0.329
R10879 GND.n12126 GND.n12124 0.329
R10880 GND.n12486 GND.n12480 0.329
R10881 GND.n13196 GND.n13195 0.329
R10882 GND.n12847 GND.n12845 0.329
R10883 GND.n7621 GND.n7619 0.329
R10884 GND.n7964 GND.n7963 0.329
R10885 GND.n15892 GND.n15890 0.329
R10886 GND.n16233 GND.n16232 0.329
R10887 GND.n10372 GND.n1172 0.329
R10888 GND.n832 GND.n830 0.329
R10889 GND.n10363 GND.n1174 0.329
R10890 GND.n9933 GND.n9932 0.329
R10891 GND.n10334 GND.n1176 0.329
R10892 GND.n9954 GND.n1528 0.329
R10893 GND.n10325 GND.n10309 0.329
R10894 GND.n8879 GND.n8872 0.329
R10895 GND.n8891 GND.n8889 0.329
R10896 GND.n9232 GND.n9231 0.329
R10897 GND.n4544 GND.n4538 0.329
R10898 GND.n5432 GND.n1915 0.329
R10899 GND.n4569 GND.n3953 0.329
R10900 GND.n5235 GND.n1917 0.329
R10901 GND.n5792 GND.n5791 0.329
R10902 GND.n5451 GND.n5449 0.329
R10903 GND.n17652 GND.n17651 0.312
R10904 GND.n14914 GND.n10573 0.28
R10905 GND.n3180 GND.n3149 0.28
R10906 GND.n5098 GND.n4923 0.28
R10907 GND.n7043 GND.n7042 0.259
R10908 GND.n8093 GND.n8092 0.259
R10909 GND.n13393 GND.n13392 0.259
R10910 GND.n12645 GND.n12644 0.259
R10911 GND.n12586 GND.n12585 0.259
R10912 GND.n13452 GND.n13451 0.259
R10913 GND.n12892 GND.n12889 0.259
R10914 GND.n11774 GND.n11771 0.259
R10915 GND.n12449 GND.n12446 0.259
R10916 GND.n12362 GND.n12361 0.259
R10917 GND.n13086 GND.n13085 0.259
R10918 GND.n12967 GND.n12966 0.259
R10919 GND.n7732 GND.n7731 0.259
R10920 GND.n7919 GND.n7916 0.259
R10921 GND.n8034 GND.n8033 0.259
R10922 GND.n7102 GND.n7101 0.259
R10923 GND.n6277 GND.n6276 0.259
R10924 GND.n11258 GND.n11257 0.259
R10925 GND.n13665 GND.n13664 0.259
R10926 GND.n14857 GND.n14856 0.259
R10927 GND.n16204 GND.n16201 0.259
R10928 GND.n876 GND.n873 0.259
R10929 GND.n934 GND.n933 0.259
R10930 GND.n1085 GND.n1084 0.259
R10931 GND.n9904 GND.n9901 0.259
R10932 GND.n1514 GND.n1511 0.259
R10933 GND.n1428 GND.n1427 0.259
R10934 GND.n1277 GND.n1276 0.259
R10935 GND.n8818 GND.n8817 0.259
R10936 GND.n10079 GND.n10078 0.259
R10937 GND.n9203 GND.n9200 0.259
R10938 GND.n5495 GND.n5492 0.259
R10939 GND.n4236 GND.n4233 0.259
R10940 GND.n4294 GND.n4293 0.259
R10941 GND.n15605 GND.n15604 0.259
R10942 GND.n4695 GND.n4694 0.259
R10943 GND.n5041 GND.n5040 0.259
R10944 GND.n4982 GND.n4981 0.259
R10945 GND.n4636 GND.n4635 0.259
R10946 GND.n3037 GND.n3036 0.259
R10947 GND.n3237 GND.n3236 0.259
R10948 GND.n14798 GND.n14797 0.259
R10949 GND.n10461 GND.n10460 0.259
R10950 GND.n15664 GND.n15663 0.259
R10951 GND.n15168 GND.n15167 0.259
R10952 GND.n3644 GND.n3641 0.259
R10953 GND.n3866 GND.n3865 0.259
R10954 GND.n5553 GND.n5552 0.259
R10955 GND.n5704 GND.n5703 0.259
R10956 GND.n11923 GND.n11921 0.241
R10957 GND.n12302 GND.n12299 0.241
R10958 GND.n13028 GND.n13026 0.241
R10959 GND.n7791 GND.n7788 0.241
R10960 GND.n16404 GND.n16319 0.229
R10961 GND.n16665 GND.n16580 0.229
R10962 GND.n16926 GND.n16841 0.229
R10963 GND.n17187 GND.n17102 0.229
R10964 GND.n17448 GND.n17363 0.229
R10965 GND.n16398 GND.n16397 0.228
R10966 GND.n16659 GND.n16658 0.228
R10967 GND.n16920 GND.n16919 0.228
R10968 GND.n17181 GND.n17180 0.228
R10969 GND.n17442 GND.n17441 0.228
R10970 GND.n16571 GND.n16570 0.228
R10971 GND.n16832 GND.n16831 0.228
R10972 GND.n17093 GND.n17092 0.228
R10973 GND.n17354 GND.n17353 0.228
R10974 GND.n17615 GND.n17614 0.228
R10975 GND.n16486 GND.n16484 0.227
R10976 GND.n16747 GND.n16745 0.227
R10977 GND.n17008 GND.n17006 0.227
R10978 GND.n17269 GND.n17267 0.227
R10979 GND.n17530 GND.n17528 0.227
R10980 GND.n15545 GND.n14028 0.222
R10981 GND.n625 GND.n540 0.215
R10982 GND.n367 GND.n282 0.215
R10983 GND.n109 GND.n24 0.215
R10984 GND.n619 GND.n618 0.214
R10985 GND.n361 GND.n360 0.214
R10986 GND.n103 GND.n102 0.214
R10987 GND.n17860 GND.n17705 0.214
R10988 GND.n789 GND.n786 0.213
R10989 GND.n531 GND.n528 0.213
R10990 GND.n273 GND.n270 0.213
R10991 GND.n705 GND.n703 0.213
R10992 GND.n447 GND.n445 0.213
R10993 GND.n189 GND.n187 0.213
R10994 GND.n9520 GND.n9519 0.212
R10995 GND.n12710 GND.n12704 0.21
R10996 GND.n13723 GND.n13722 0.21
R10997 GND.n13510 GND.n13509 0.21
R10998 GND.n13549 GND.n13546 0.21
R10999 GND.n6524 GND.n6523 0.21
R11000 GND.n8151 GND.n8150 0.21
R11001 GND.n8879 GND.n8406 0.21
R11002 GND.n7200 GND.n7199 0.21
R11003 GND.n7163 GND.n7162 0.21
R11004 GND.n8703 GND.n8702 0.21
R11005 GND.n10134 GND.n1182 0.21
R11006 GND.n3180 GND.n3179 0.21
R11007 GND.n5099 GND.n5098 0.21
R11008 GND.n3149 GND.n2673 0.21
R11009 GND.n4923 GND.n4922 0.21
R11010 GND.n15758 GND.n10573 0.21
R11011 GND.n14920 GND.n14914 0.21
R11012 GND.n5422 GND.n5421 0.19
R11013 GND.n5280 GND.n5279 0.19
R11014 GND.n1555 GND.n1554 0.19
R11015 GND.n16305 GND.n16304 0.19
R11016 GND.n16251 GND.n16250 0.19
R11017 GND.n16272 GND.n16263 0.19
R11018 GND.n9566 GND.n9565 0.19
R11019 GND.n9562 GND.n9561 0.19
R11020 GND.n5322 GND.n5321 0.19
R11021 GND.n5335 GND.n5334 0.19
R11022 GND.n5408 GND.n5394 0.19
R11023 GND.n5373 GND.n5372 0.19
R11024 GND.n5408 GND.n5407 0.19
R11025 GND.n16272 GND.n16271 0.19
R11026 GND.n16288 GND.n16287 0.19
R11027 GND.n1565 GND.n1564 0.19
R11028 GND.n9565 GND.n1539 0.19
R11029 GND.n5290 GND.n5289 0.19
R11030 GND.n5322 GND.n5260 0.19
R11031 GND.n5418 GND.n5417 0.19
R11032 GND.n3496 GND.n3489 0.185
R11033 GND.n15456 GND.n15455 0.185
R11034 GND.n5420 GND.n5419 0.18
R11035 GND.n5337 GND.n5336 0.18
R11036 GND.n9551 GND.n9550 0.18
R11037 GND.n802 GND.n801 0.18
R11038 GND.n16252 GND.n800 0.178
R11039 GND.n1556 GND.n1540 0.178
R11040 GND.n5281 GND.n5261 0.178
R11041 GND.n5374 GND.n5339 0.178
R11042 GND.n5346 GND.n5345 0.171
R11043 GND.n17663 GND.n17660 0.171
R11044 GND.n17658 GND.n17657 0.171
R11045 GND.n794 GND.n793 0.171
R11046 GND.n798 GND.n795 0.171
R11047 GND.n5342 GND.n5341 0.171
R11048 GND.n5352 GND.n5351 0.171
R11049 GND.n5356 GND.n5353 0.171
R11050 GND.n7378 GND.n7375 0.169
R11051 GND.n14671 GND.n14668 0.168
R11052 GND.n14620 GND.n14617 0.168
R11053 GND.n10626 GND.n10623 0.168
R11054 GND.n15484 GND.n15482 0.168
R11055 GND.n14348 GND.n14345 0.168
R11056 GND.n14265 GND.n14263 0.168
R11057 GND.n3570 GND.n3568 0.168
R11058 GND.n4838 GND.n4835 0.168
R11059 GND.n10758 GND.n10755 0.168
R11060 GND.n13948 GND.n13945 0.168
R11061 GND.n13820 GND.n13818 0.168
R11062 GND.n13774 GND.n13771 0.168
R11063 GND.n12761 GND.n12758 0.168
R11064 GND.n11674 GND.n11671 0.168
R11065 GND.n11570 GND.n11567 0.168
R11066 GND.n11062 GND.n11060 0.168
R11067 GND.n13275 GND.n13273 0.168
R11068 GND.n11370 GND.n11367 0.168
R11069 GND.n8210 GND.n8207 0.168
R11070 GND.n8299 GND.n8296 0.168
R11071 GND.n5984 GND.n5981 0.168
R11072 GND.n6461 GND.n6459 0.168
R11073 GND.n6896 GND.n6893 0.168
R11074 GND.n6661 GND.n6658 0.168
R11075 GND.n6758 GND.n6755 0.168
R11076 GND.n7482 GND.n7479 0.168
R11077 GND.n7536 GND.n7534 0.168
R11078 GND.n9343 GND.n9340 0.168
R11079 GND.n1748 GND.n1745 0.168
R11080 GND.n9470 GND.n9468 0.168
R11081 GND.n1850 GND.n1847 0.168
R11082 GND.n8650 GND.n8648 0.168
R11083 GND.n2541 GND.n2538 0.168
R11084 GND.n3451 GND.n3449 0.168
R11085 GND.n2447 GND.n2444 0.168
R11086 GND.n2379 GND.n2376 0.168
R11087 GND.n5150 GND.n5147 0.168
R11088 GND.n2108 GND.n2106 0.168
R11089 GND.n2188 GND.n2185 0.168
R11090 GND.n2917 GND.n2915 0.168
R11091 GND.n15825 GND.n15823 0.168
R11092 GND.n15380 GND.n15378 0.168
R11093 GND.n14971 GND.n14968 0.168
R11094 GND.n15066 GND.n15064 0.168
R11095 GND.n14016 GND.n14013 0.166
R11096 GND.n14019 GND.n14016 0.166
R11097 GND.n14022 GND.n14019 0.166
R11098 GND.n14025 GND.n14022 0.166
R11099 GND.n14028 GND.n14025 0.166
R11100 GND.n8394 GND.n8391 0.166
R11101 GND.n8397 GND.n8394 0.166
R11102 GND.n8400 GND.n8397 0.166
R11103 GND.n8403 GND.n8400 0.166
R11104 GND.n8406 GND.n8403 0.166
R11105 GND.n11921 GND.n11918 0.159
R11106 GND.n11918 GND.n11915 0.159
R11107 GND.n12305 GND.n12302 0.159
R11108 GND.n12308 GND.n12305 0.159
R11109 GND.n13026 GND.n13023 0.159
R11110 GND.n13023 GND.n13020 0.159
R11111 GND.n7794 GND.n7791 0.159
R11112 GND.n7797 GND.n7794 0.159
R11113 GND.n11968 GND.n11967 0.157
R11114 GND.n12050 GND.n12049 0.157
R11115 GND.n11794 GND.n11791 0.157
R11116 GND.n12261 GND.n12260 0.157
R11117 GND.n12154 GND.n12153 0.157
R11118 GND.n13074 GND.n13073 0.157
R11119 GND.n7749 GND.n7748 0.157
R11120 GND.n7939 GND.n7936 0.157
R11121 GND.n7307 GND.n7306 0.157
R11122 GND.n6265 GND.n6264 0.157
R11123 GND.n7273 GND.n7272 0.157
R11124 GND.n11246 GND.n11245 0.157
R11125 GND.n13653 GND.n13652 0.157
R11126 GND.n9003 GND.n9002 0.157
R11127 GND.n9704 GND.n9703 0.157
R11128 GND.n16004 GND.n16003 0.157
R11129 GND.n15913 GND.n15912 0.157
R11130 GND.n16208 GND.n16205 0.157
R11131 GND.n1073 GND.n1072 0.157
R11132 GND.n9613 GND.n9612 0.157
R11133 GND.n9908 GND.n9905 0.157
R11134 GND.n1294 GND.n1293 0.157
R11135 GND.n10241 GND.n10240 0.157
R11136 GND.n10207 GND.n10206 0.157
R11137 GND.n8511 GND.n8510 0.157
R11138 GND.n8806 GND.n8805 0.157
R11139 GND.n8477 GND.n8476 0.157
R11140 GND.n10067 GND.n10066 0.157
R11141 GND.n8912 GND.n8911 0.157
R11142 GND.n9207 GND.n9204 0.157
R11143 GND.n4433 GND.n4432 0.157
R11144 GND.n4508 GND.n4507 0.157
R11145 GND.n3049 GND.n3048 0.157
R11146 GND.n3249 GND.n3248 0.157
R11147 GND.n10473 GND.n10472 0.157
R11148 GND.n15180 GND.n15179 0.157
R11149 GND.n3648 GND.n3645 0.157
R11150 GND.n3854 GND.n3853 0.157
R11151 GND.n5692 GND.n5691 0.157
R11152 GND.n11315 GND.n11312 0.153
R11153 GND.n15282 GND.n15279 0.153
R11154 GND.n2685 GND.n2680 0.151
R11155 GND.n2690 GND.n2685 0.151
R11156 GND.n2695 GND.n2690 0.151
R11157 GND.n2700 GND.n2695 0.151
R11158 GND.n2705 GND.n2700 0.151
R11159 GND.n2708 GND.n2705 0.151
R11160 GND.n2713 GND.n2708 0.151
R11161 GND.n2718 GND.n2713 0.151
R11162 GND.n2723 GND.n2718 0.151
R11163 GND.n2730 GND.n2723 0.151
R11164 GND.n2759 GND.n2754 0.151
R11165 GND.n2764 GND.n2759 0.151
R11166 GND.n2769 GND.n2764 0.151
R11167 GND.n2774 GND.n2769 0.151
R11168 GND.n2777 GND.n2774 0.151
R11169 GND.n2782 GND.n2777 0.151
R11170 GND.n2787 GND.n2782 0.151
R11171 GND.n2792 GND.n2787 0.151
R11172 GND.n2797 GND.n2792 0.151
R11173 GND.n2804 GND.n2797 0.151
R11174 GND.n2806 GND.n2804 0.151
R11175 GND.n2809 GND.n2806 0.151
R11176 GND.n2814 GND.n2809 0.151
R11177 GND.n2817 GND.n2814 0.151
R11178 GND.n2820 GND.n2817 0.151
R11179 GND.n2823 GND.n2820 0.151
R11180 GND.n2827 GND.n2823 0.151
R11181 GND.n2830 GND.n2827 0.151
R11182 GND.n2833 GND.n2830 0.151
R11183 GND.n2836 GND.n2833 0.151
R11184 GND.n2839 GND.n2836 0.151
R11185 GND.n3971 GND.n3964 0.151
R11186 GND.n3978 GND.n3971 0.151
R11187 GND.n3985 GND.n3978 0.151
R11188 GND.n3992 GND.n3985 0.151
R11189 GND.n4006 GND.n3992 0.151
R11190 GND.n4013 GND.n4006 0.151
R11191 GND.n4020 GND.n4013 0.151
R11192 GND.n4027 GND.n4020 0.151
R11193 GND.n4034 GND.n4027 0.151
R11194 GND.n4044 GND.n4034 0.151
R11195 GND.n4081 GND.n4074 0.151
R11196 GND.n4088 GND.n4081 0.151
R11197 GND.n4095 GND.n4088 0.151
R11198 GND.n4102 GND.n4095 0.151
R11199 GND.n4116 GND.n4102 0.151
R11200 GND.n4123 GND.n4116 0.151
R11201 GND.n4130 GND.n4123 0.151
R11202 GND.n4137 GND.n4130 0.151
R11203 GND.n4144 GND.n4137 0.151
R11204 GND.n4154 GND.n4144 0.151
R11205 GND.n4156 GND.n4154 0.151
R11206 GND.n4161 GND.n4156 0.151
R11207 GND.n4165 GND.n4161 0.151
R11208 GND.n4168 GND.n4165 0.151
R11209 GND.n4171 GND.n4168 0.151
R11210 GND.n4174 GND.n4171 0.151
R11211 GND.n4177 GND.n4174 0.151
R11212 GND.n4180 GND.n4177 0.151
R11213 GND.n4183 GND.n4180 0.151
R11214 GND.n4186 GND.n4183 0.151
R11215 GND.n4189 GND.n4186 0.151
R11216 GND.n14834 GND.n14826 0.15
R11217 GND.n6255 GND.n6247 0.15
R11218 GND.n12622 GND.n12614 0.15
R11219 GND.n11236 GND.n11228 0.15
R11220 GND.n13643 GND.n13635 0.15
R11221 GND.n13429 GND.n13420 0.15
R11222 GND.n11955 GND.n11954 0.15
R11223 GND.n11915 GND.n11912 0.15
R11224 GND.n11882 GND.n11881 0.15
R11225 GND.n12267 GND.n12266 0.15
R11226 GND.n12310 GND.n12308 0.15
R11227 GND.n12340 GND.n12339 0.15
R11228 GND.n13061 GND.n13060 0.15
R11229 GND.n13020 GND.n13017 0.15
R11230 GND.n12987 GND.n12986 0.15
R11231 GND.n7755 GND.n7754 0.15
R11232 GND.n7799 GND.n7797 0.15
R11233 GND.n7829 GND.n7828 0.15
R11234 GND.n8070 GND.n8061 0.15
R11235 GND.n7079 GND.n7070 0.15
R11236 GND.n7297 GND.n7288 0.15
R11237 GND.n16013 GND.n16009 0.15
R11238 GND.n16114 GND.n16106 0.15
R11239 GND.n1060 GND.n1059 0.15
R11240 GND.n970 GND.n962 0.15
R11241 GND.n9713 GND.n9709 0.15
R11242 GND.n9814 GND.n9806 0.15
R11243 GND.n1303 GND.n1299 0.15
R11244 GND.n1405 GND.n1396 0.15
R11245 GND.n10231 GND.n10222 0.15
R11246 GND.n8796 GND.n8788 0.15
R11247 GND.n8501 GND.n8492 0.15
R11248 GND.n10057 GND.n10049 0.15
R11249 GND.n9012 GND.n9008 0.15
R11250 GND.n9113 GND.n9105 0.15
R11251 GND.n4420 GND.n4419 0.15
R11252 GND.n4330 GND.n4322 0.15
R11253 GND.n3271 GND.n3263 0.15
R11254 GND.n5018 GND.n5010 0.15
R11255 GND.n4672 GND.n4664 0.15
R11256 GND.n3071 GND.n3063 0.15
R11257 GND.n10495 GND.n10487 0.15
R11258 GND.n15641 GND.n15632 0.15
R11259 GND.n15202 GND.n15194 0.15
R11260 GND.n3841 GND.n3840 0.15
R11261 GND.n3751 GND.n3743 0.15
R11262 GND.n5679 GND.n5678 0.15
R11263 GND.n5589 GND.n5581 0.15
R11264 GND.n12836 GND.n12524 0.149
R11265 GND.n13345 GND.n13337 0.149
R11266 GND.n2736 GND.n2730 0.145
R11267 GND.n4050 GND.n4044 0.145
R11268 GND.n2742 GND.n2741 0.143
R11269 GND.n4059 GND.n4058 0.143
R11270 GND.n3352 GND.n3349 0.142
R11271 GND.n14719 GND.n14717 0.141
R11272 GND.n15296 GND.n14402 0.141
R11273 GND.n15536 GND.n15530 0.141
R11274 GND.n15726 GND.n10714 0.141
R11275 GND.n15750 GND.n10575 0.141
R11276 GND.n4761 GND.n3616 0.141
R11277 GND.n4789 GND.n4787 0.141
R11278 GND.n10877 GND.n10875 0.141
R11279 GND.n13996 GND.n13994 0.141
R11280 GND.n13869 GND.n13866 0.141
R11281 GND.n13725 GND.n13723 0.141
R11282 GND.n12712 GND.n12710 0.141
R11283 GND.n13518 GND.n11720 0.141
R11284 GND.n13542 GND.n11616 0.141
R11285 GND.n11126 GND.n11108 0.141
R11286 GND.n13330 GND.n13321 0.141
R11287 GND.n11321 GND.n11319 0.141
R11288 GND.n8161 GND.n8159 0.141
R11289 GND.n8250 GND.n8248 0.141
R11290 GND.n6117 GND.n5901 0.141
R11291 GND.n6047 GND.n6030 0.141
R11292 GND.n8382 GND.n5824 0.141
R11293 GND.n7171 GND.n6942 0.141
R11294 GND.n7195 GND.n6707 0.141
R11295 GND.n7433 GND.n7431 0.141
R11296 GND.n7583 GND.n7582 0.141
R11297 GND.n9294 GND.n1182 0.141
R11298 GND.n1699 GND.n1697 0.141
R11299 GND.n9421 GND.n9419 0.141
R11300 GND.n9259 GND.n1896 0.141
R11301 GND.n8702 GND.n8696 0.141
R11302 GND.n2492 GND.n2490 0.141
R11303 GND.n3402 GND.n3400 0.141
R11304 GND.n3366 GND.n2631 0.141
R11305 GND.n3179 GND.n3155 0.141
R11306 GND.n5101 GND.n5099 0.141
R11307 GND.n4918 GND.n1941 0.141
R11308 GND.n2669 GND.n2658 0.141
R11309 GND.n2969 GND.n2963 0.141
R11310 GND.n15872 GND.n15871 0.141
R11311 GND.n15429 GND.n15426 0.141
R11312 GND.n14922 GND.n14920 0.141
R11313 GND.n15113 GND.n15112 0.141
R11314 GND.n7618 GND.n7613 0.14
R11315 GND.n7613 GND.n7610 0.14
R11316 GND.n7610 GND.n7607 0.14
R11317 GND.n7607 GND.n7604 0.14
R11318 GND.n7604 GND.n7601 0.14
R11319 GND.n7601 GND.n7598 0.14
R11320 GND.n12123 GND.n12120 0.14
R11321 GND.n12114 GND.n12111 0.14
R11322 GND.n12111 GND.n12108 0.14
R11323 GND.n12108 GND.n12105 0.14
R11324 GND.n12105 GND.n12102 0.14
R11325 GND.n12102 GND.n12099 0.14
R11326 GND.n12099 GND.n11729 0.14
R11327 GND.n13204 GND.n13201 0.14
R11328 GND.n6143 GND.n6138 0.14
R11329 GND.n6138 GND.n6135 0.14
R11330 GND.n6135 GND.n6132 0.14
R11331 GND.n6132 GND.n6129 0.14
R11332 GND.n6129 GND.n6126 0.14
R11333 GND.n6126 GND.n6123 0.14
R11334 GND.n12494 GND.n12489 0.14
R11335 GND.n12501 GND.n12498 0.14
R11336 GND.n12504 GND.n12501 0.14
R11337 GND.n12507 GND.n12504 0.14
R11338 GND.n12510 GND.n12507 0.14
R11339 GND.n12513 GND.n12510 0.14
R11340 GND.n12516 GND.n12513 0.14
R11341 GND.n12844 GND.n12839 0.14
R11342 GND.n14417 GND.n812 0.14
R11343 GND.n9944 GND.n9941 0.14
R11344 GND.n9941 GND.n9938 0.14
R11345 GND.n829 GND.n826 0.14
R11346 GND.n826 GND.n807 0.14
R11347 GND.n9953 GND.n9948 0.14
R11348 GND.n5306 GND.n1904 0.14
R11349 GND.n4577 GND.n4574 0.14
R11350 GND.n4568 GND.n4565 0.14
R11351 GND.n4565 GND.n4562 0.14
R11352 GND.n4558 GND.n4553 0.14
R11353 GND.n4553 GND.n4550 0.14
R11354 GND.n4550 GND.n4547 0.14
R11355 GND.n4543 GND.n1910 0.14
R11356 GND.n5800 GND.n5797 0.14
R11357 GND.n5803 GND.n5800 0.14
R11358 GND.n5806 GND.n5803 0.14
R11359 GND.n5809 GND.n5806 0.14
R11360 GND.n5812 GND.n5809 0.14
R11361 GND.n5815 GND.n5812 0.14
R11362 GND.n5820 GND.n5815 0.14
R11363 GND.n8888 GND.n8885 0.14
R11364 GND.n8878 GND.n8875 0.14
R11365 GND.n10315 GND.n10312 0.14
R11366 GND.n10318 GND.n10315 0.14
R11367 GND.n10321 GND.n10318 0.14
R11368 GND.n10324 GND.n10321 0.14
R11369 GND.n10333 GND.n10330 0.14
R11370 GND.n10342 GND.n10339 0.14
R11371 GND.n10345 GND.n10342 0.14
R11372 GND.n10348 GND.n10345 0.14
R11373 GND.n10351 GND.n10348 0.14
R11374 GND.n10354 GND.n10351 0.14
R11375 GND.n10357 GND.n10354 0.14
R11376 GND.n10362 GND.n10357 0.14
R11377 GND.n10371 GND.n10366 0.14
R11378 GND.n10378 GND.n10375 0.14
R11379 GND.n10381 GND.n10378 0.14
R11380 GND.n10384 GND.n10381 0.14
R11381 GND.n10387 GND.n10384 0.14
R11382 GND.n10390 GND.n10387 0.14
R11383 GND.n10393 GND.n10390 0.14
R11384 GND.n15889 GND.n15884 0.14
R11385 GND.n5440 GND.n5437 0.14
R11386 GND.n5448 GND.n5443 0.14
R11387 GND.n5297 GND.n5294 0.14
R11388 GND.n5300 GND.n5297 0.14
R11389 GND.n5234 GND.n5229 0.14
R11390 GND.n5241 GND.n5238 0.14
R11391 GND.n5244 GND.n5241 0.14
R11392 GND.n5303 GND.n5300 0.139
R11393 GND.n13531 GND.n13528 0.132
R11394 GND.n13196 GND.n11729 0.132
R11395 GND.n12845 GND.n12516 0.132
R11396 GND.n7192 GND.n7184 0.132
R11397 GND.n16236 GND.n16233 0.132
R11398 GND.n15747 GND.n15739 0.132
R11399 GND.n15890 GND.n10393 0.132
R11400 GND.n7162 GND.n5851 0.131
R11401 GND.n7200 GND.n6527 0.131
R11402 GND.n13552 GND.n13549 0.131
R11403 GND.n13509 GND.n11724 0.131
R11404 GND.n12540 GND.n12524 0.13
R11405 GND.n13347 GND.n13345 0.13
R11406 GND.n15717 GND.n15708 0.13
R11407 GND.n15124 GND.n15122 0.13
R11408 GND.n9240 GND.n9235 0.13
R11409 GND.n5307 GND.n5303 0.13
R11410 GND.n2981 GND.n2979 0.13
R11411 GND.n10325 GND.n10324 0.128
R11412 GND.n14678 GND.n14676 0.127
R11413 GND.n14685 GND.n14683 0.127
R11414 GND.n14692 GND.n14690 0.127
R11415 GND.n14699 GND.n14697 0.127
R11416 GND.n14706 GND.n14704 0.127
R11417 GND.n14713 GND.n14711 0.127
R11418 GND.n14613 GND.n14610 0.127
R11419 GND.n14606 GND.n14603 0.127
R11420 GND.n14599 GND.n14596 0.127
R11421 GND.n14384 GND.n14382 0.127
R11422 GND.n14391 GND.n14389 0.127
R11423 GND.n14398 GND.n14396 0.127
R11424 GND.n10584 GND.n10581 0.127
R11425 GND.n10591 GND.n10588 0.127
R11426 GND.n10598 GND.n10595 0.127
R11427 GND.n10605 GND.n10602 0.127
R11428 GND.n10612 GND.n10609 0.127
R11429 GND.n10619 GND.n10616 0.127
R11430 GND.n15526 GND.n15524 0.127
R11431 GND.n15519 GND.n15517 0.127
R11432 GND.n15512 GND.n15510 0.127
R11433 GND.n15505 GND.n15503 0.127
R11434 GND.n15498 GND.n15496 0.127
R11435 GND.n15491 GND.n15489 0.127
R11436 GND.n14341 GND.n14338 0.127
R11437 GND.n14334 GND.n14331 0.127
R11438 GND.n14327 GND.n14324 0.127
R11439 GND.n10703 GND.n10701 0.127
R11440 GND.n10710 GND.n10708 0.127
R11441 GND.n14258 GND.n14255 0.127
R11442 GND.n14251 GND.n14248 0.127
R11443 GND.n14244 GND.n14241 0.127
R11444 GND.n14237 GND.n14234 0.127
R11445 GND.n14230 GND.n14227 0.127
R11446 GND.n14223 GND.n14220 0.127
R11447 GND.n14914 GND.n14913 0.127
R11448 GND.n14739 GND.n14737 0.127
R11449 GND.n3612 GND.n3610 0.127
R11450 GND.n3605 GND.n3603 0.127
R11451 GND.n3598 GND.n3596 0.127
R11452 GND.n3591 GND.n3589 0.127
R11453 GND.n3584 GND.n3582 0.127
R11454 GND.n3577 GND.n3575 0.127
R11455 GND.n4796 GND.n4793 0.127
R11456 GND.n4803 GND.n4800 0.127
R11457 GND.n4810 GND.n4807 0.127
R11458 GND.n4817 GND.n4814 0.127
R11459 GND.n4824 GND.n4821 0.127
R11460 GND.n4831 GND.n4828 0.127
R11461 GND.n6524 GND.n6331 0.127
R11462 GND.n8388 GND.n5822 0.127
R11463 GND.n12704 GND.n12701 0.127
R11464 GND.n10751 GND.n10748 0.127
R11465 GND.n10744 GND.n10741 0.127
R11466 GND.n10857 GND.n10855 0.127
R11467 GND.n10864 GND.n10862 0.127
R11468 GND.n10871 GND.n10869 0.127
R11469 GND.n13955 GND.n13953 0.127
R11470 GND.n13962 GND.n13960 0.127
R11471 GND.n13969 GND.n13967 0.127
R11472 GND.n13976 GND.n13974 0.127
R11473 GND.n13983 GND.n13981 0.127
R11474 GND.n13990 GND.n13988 0.127
R11475 GND.n13862 GND.n13860 0.127
R11476 GND.n13855 GND.n13853 0.127
R11477 GND.n13848 GND.n13846 0.127
R11478 GND.n13841 GND.n13839 0.127
R11479 GND.n13834 GND.n13832 0.127
R11480 GND.n13827 GND.n13825 0.127
R11481 GND.n13732 GND.n13729 0.127
R11482 GND.n13739 GND.n13736 0.127
R11483 GND.n13746 GND.n13743 0.127
R11484 GND.n13753 GND.n13750 0.127
R11485 GND.n13760 GND.n13757 0.127
R11486 GND.n13767 GND.n13764 0.127
R11487 GND.n13549 GND.n11006 0.127
R11488 GND.n13722 GND.n13719 0.127
R11489 GND.n14010 GND.n10717 0.127
R11490 GND.n12719 GND.n12716 0.127
R11491 GND.n12726 GND.n12723 0.127
R11492 GND.n12733 GND.n12730 0.127
R11493 GND.n12740 GND.n12737 0.127
R11494 GND.n12747 GND.n12744 0.127
R11495 GND.n12754 GND.n12751 0.127
R11496 GND.n11681 GND.n11679 0.127
R11497 GND.n11688 GND.n11686 0.127
R11498 GND.n11695 GND.n11693 0.127
R11499 GND.n11702 GND.n11700 0.127
R11500 GND.n11709 GND.n11707 0.127
R11501 GND.n11716 GND.n11714 0.127
R11502 GND.n11577 GND.n11575 0.127
R11503 GND.n11584 GND.n11582 0.127
R11504 GND.n11591 GND.n11589 0.127
R11505 GND.n11598 GND.n11596 0.127
R11506 GND.n11605 GND.n11603 0.127
R11507 GND.n11612 GND.n11610 0.127
R11508 GND.n11104 GND.n11102 0.127
R11509 GND.n11097 GND.n11095 0.127
R11510 GND.n11090 GND.n11088 0.127
R11511 GND.n11083 GND.n11081 0.127
R11512 GND.n11076 GND.n11074 0.127
R11513 GND.n11069 GND.n11067 0.127
R11514 GND.n13317 GND.n13315 0.127
R11515 GND.n13310 GND.n13308 0.127
R11516 GND.n13303 GND.n13301 0.127
R11517 GND.n13296 GND.n13294 0.127
R11518 GND.n13289 GND.n13287 0.127
R11519 GND.n13282 GND.n13280 0.127
R11520 GND.n11328 GND.n11325 0.127
R11521 GND.n11335 GND.n11332 0.127
R11522 GND.n11342 GND.n11339 0.127
R11523 GND.n11349 GND.n11346 0.127
R11524 GND.n11356 GND.n11353 0.127
R11525 GND.n11363 GND.n11360 0.127
R11526 GND.n13509 GND.n13508 0.127
R11527 GND.n8168 GND.n8165 0.127
R11528 GND.n8175 GND.n8172 0.127
R11529 GND.n8182 GND.n8179 0.127
R11530 GND.n8189 GND.n8186 0.127
R11531 GND.n8196 GND.n8193 0.127
R11532 GND.n8203 GND.n8200 0.127
R11533 GND.n8257 GND.n8254 0.127
R11534 GND.n8264 GND.n8261 0.127
R11535 GND.n8271 GND.n8268 0.127
R11536 GND.n8278 GND.n8275 0.127
R11537 GND.n8285 GND.n8282 0.127
R11538 GND.n8292 GND.n8289 0.127
R11539 GND.n5862 GND.n5860 0.127
R11540 GND.n5869 GND.n5867 0.127
R11541 GND.n5876 GND.n5874 0.127
R11542 GND.n5883 GND.n5881 0.127
R11543 GND.n5890 GND.n5888 0.127
R11544 GND.n5897 GND.n5895 0.127
R11545 GND.n5991 GND.n5989 0.127
R11546 GND.n5998 GND.n5996 0.127
R11547 GND.n6005 GND.n6003 0.127
R11548 GND.n6012 GND.n6010 0.127
R11549 GND.n6019 GND.n6017 0.127
R11550 GND.n6026 GND.n6024 0.127
R11551 GND.n6454 GND.n6451 0.127
R11552 GND.n6447 GND.n6444 0.127
R11553 GND.n6440 GND.n6437 0.127
R11554 GND.n6433 GND.n6430 0.127
R11555 GND.n6426 GND.n6423 0.127
R11556 GND.n6419 GND.n6416 0.127
R11557 GND.n8150 GND.n8149 0.127
R11558 GND.n7975 GND.n7973 0.127
R11559 GND.n7587 GND.n6149 0.127
R11560 GND.n7162 GND.n7159 0.127
R11561 GND.n6903 GND.n6901 0.127
R11562 GND.n6910 GND.n6908 0.127
R11563 GND.n6917 GND.n6915 0.127
R11564 GND.n6924 GND.n6922 0.127
R11565 GND.n6931 GND.n6929 0.127
R11566 GND.n6938 GND.n6936 0.127
R11567 GND.n6668 GND.n6666 0.127
R11568 GND.n6675 GND.n6673 0.127
R11569 GND.n6682 GND.n6680 0.127
R11570 GND.n6689 GND.n6687 0.127
R11571 GND.n6696 GND.n6694 0.127
R11572 GND.n6703 GND.n6701 0.127
R11573 GND.n6716 GND.n6713 0.127
R11574 GND.n6723 GND.n6720 0.127
R11575 GND.n6730 GND.n6727 0.127
R11576 GND.n6737 GND.n6734 0.127
R11577 GND.n6744 GND.n6741 0.127
R11578 GND.n6751 GND.n6748 0.127
R11579 GND.n7440 GND.n7437 0.127
R11580 GND.n7447 GND.n7444 0.127
R11581 GND.n7454 GND.n7451 0.127
R11582 GND.n7461 GND.n7458 0.127
R11583 GND.n7468 GND.n7465 0.127
R11584 GND.n7475 GND.n7472 0.127
R11585 GND.n7578 GND.n7576 0.127
R11586 GND.n7571 GND.n7569 0.127
R11587 GND.n7564 GND.n7562 0.127
R11588 GND.n7557 GND.n7555 0.127
R11589 GND.n7550 GND.n7548 0.127
R11590 GND.n7543 GND.n7541 0.127
R11591 GND.n7202 GND.n7200 0.127
R11592 GND.n8703 GND.n8579 0.127
R11593 GND.n9241 GND.n1899 0.127
R11594 GND.n9301 GND.n9298 0.127
R11595 GND.n9308 GND.n9305 0.127
R11596 GND.n9315 GND.n9312 0.127
R11597 GND.n9322 GND.n9319 0.127
R11598 GND.n9329 GND.n9326 0.127
R11599 GND.n9336 GND.n9333 0.127
R11600 GND.n1706 GND.n1703 0.127
R11601 GND.n1713 GND.n1710 0.127
R11602 GND.n1720 GND.n1717 0.127
R11603 GND.n1727 GND.n1724 0.127
R11604 GND.n1734 GND.n1731 0.127
R11605 GND.n1741 GND.n1738 0.127
R11606 GND.n9463 GND.n9460 0.127
R11607 GND.n9456 GND.n9453 0.127
R11608 GND.n9449 GND.n9446 0.127
R11609 GND.n9442 GND.n9439 0.127
R11610 GND.n9435 GND.n9432 0.127
R11611 GND.n9428 GND.n9425 0.127
R11612 GND.n1857 GND.n1855 0.127
R11613 GND.n1864 GND.n1862 0.127
R11614 GND.n1871 GND.n1869 0.127
R11615 GND.n1878 GND.n1876 0.127
R11616 GND.n1885 GND.n1883 0.127
R11617 GND.n1892 GND.n1890 0.127
R11618 GND.n8692 GND.n8690 0.127
R11619 GND.n8685 GND.n8683 0.127
R11620 GND.n8678 GND.n8676 0.127
R11621 GND.n8671 GND.n8669 0.127
R11622 GND.n8664 GND.n8662 0.127
R11623 GND.n8657 GND.n8655 0.127
R11624 GND.n10134 GND.n10133 0.127
R11625 GND.n9965 GND.n9963 0.127
R11626 GND.n2499 GND.n2496 0.127
R11627 GND.n2506 GND.n2503 0.127
R11628 GND.n2513 GND.n2510 0.127
R11629 GND.n2520 GND.n2517 0.127
R11630 GND.n2527 GND.n2524 0.127
R11631 GND.n2534 GND.n2531 0.127
R11632 GND.n3182 GND.n3180 0.127
R11633 GND.n3444 GND.n3441 0.127
R11634 GND.n3437 GND.n3434 0.127
R11635 GND.n3430 GND.n3427 0.127
R11636 GND.n3423 GND.n3420 0.127
R11637 GND.n3416 GND.n3413 0.127
R11638 GND.n3409 GND.n3406 0.127
R11639 GND.n2440 GND.n2437 0.127
R11640 GND.n2433 GND.n2430 0.127
R11641 GND.n2426 GND.n2423 0.127
R11642 GND.n2613 GND.n2611 0.127
R11643 GND.n2620 GND.n2618 0.127
R11644 GND.n2627 GND.n2625 0.127
R11645 GND.n2344 GND.n2341 0.127
R11646 GND.n2351 GND.n2348 0.127
R11647 GND.n2358 GND.n2355 0.127
R11648 GND.n2365 GND.n2362 0.127
R11649 GND.n2372 GND.n2369 0.127
R11650 GND.n5098 GND.n5097 0.127
R11651 GND.n5226 GND.n1919 0.127
R11652 GND.n5108 GND.n5105 0.127
R11653 GND.n5115 GND.n5112 0.127
R11654 GND.n5122 GND.n5119 0.127
R11655 GND.n5129 GND.n5126 0.127
R11656 GND.n5136 GND.n5133 0.127
R11657 GND.n5143 GND.n5140 0.127
R11658 GND.n2101 GND.n2098 0.127
R11659 GND.n2094 GND.n2091 0.127
R11660 GND.n2087 GND.n2084 0.127
R11661 GND.n2080 GND.n2077 0.127
R11662 GND.n2073 GND.n2070 0.127
R11663 GND.n2066 GND.n2063 0.127
R11664 GND.n2181 GND.n2178 0.127
R11665 GND.n2174 GND.n2171 0.127
R11666 GND.n2167 GND.n2164 0.127
R11667 GND.n2640 GND.n2638 0.127
R11668 GND.n2647 GND.n2645 0.127
R11669 GND.n2654 GND.n2652 0.127
R11670 GND.n2959 GND.n2957 0.127
R11671 GND.n2952 GND.n2950 0.127
R11672 GND.n2945 GND.n2943 0.127
R11673 GND.n2938 GND.n2936 0.127
R11674 GND.n2931 GND.n2929 0.127
R11675 GND.n2924 GND.n2922 0.127
R11676 GND.n4752 GND.n4751 0.127
R11677 GND.n4923 GND.n1934 0.127
R11678 GND.n3149 GND.n3148 0.127
R11679 GND.n15881 GND.n10395 0.127
R11680 GND.n10573 GND.n10572 0.127
R11681 GND.n15547 GND.n15545 0.127
R11682 GND.n15867 GND.n15865 0.127
R11683 GND.n15860 GND.n15858 0.127
R11684 GND.n15853 GND.n15851 0.127
R11685 GND.n15846 GND.n15844 0.127
R11686 GND.n15839 GND.n15837 0.127
R11687 GND.n15832 GND.n15830 0.127
R11688 GND.n15422 GND.n15420 0.127
R11689 GND.n15415 GND.n15413 0.127
R11690 GND.n15408 GND.n15406 0.127
R11691 GND.n15401 GND.n15399 0.127
R11692 GND.n15394 GND.n15392 0.127
R11693 GND.n15387 GND.n15385 0.127
R11694 GND.n14929 GND.n14926 0.127
R11695 GND.n14936 GND.n14933 0.127
R11696 GND.n14943 GND.n14940 0.127
R11697 GND.n14950 GND.n14947 0.127
R11698 GND.n14957 GND.n14954 0.127
R11699 GND.n14964 GND.n14961 0.127
R11700 GND.n15108 GND.n15106 0.127
R11701 GND.n15101 GND.n15099 0.127
R11702 GND.n15094 GND.n15092 0.127
R11703 GND.n15087 GND.n15085 0.127
R11704 GND.n15080 GND.n15078 0.127
R11705 GND.n15073 GND.n15071 0.127
R11706 GND.n2754 GND.n2751 0.126
R11707 GND.n4074 GND.n4070 0.126
R11708 GND.n16237 GND.n807 0.126
R11709 GND.n2741 GND.n2738 0.125
R11710 GND.n4058 GND.n4052 0.125
R11711 GND.n4547 GND.n4544 0.125
R11712 GND.n5432 GND.n5431 0.125
R11713 GND.n9545 GND.n9544 0.125
R11714 GND.n5362 GND.n5343 0.125
R11715 GND.n9586 GND.n9577 0.119
R11716 GND.n16247 GND.n16246 0.119
R11717 GND.n5427 GND.n5424 0.119
R11718 GND.n14909 GND.n14901 0.114
R11719 GND.n14897 GND.n14888 0.114
R11720 GND.n14884 GND.n14876 0.114
R11721 GND.n14872 GND.n14863 0.114
R11722 GND.n14859 GND.n14851 0.114
R11723 GND.n14815 GND.n14813 0.114
R11724 GND.n14802 GND.n14800 0.114
R11725 GND.n14790 GND.n14788 0.114
R11726 GND.n14777 GND.n14775 0.114
R11727 GND.n14765 GND.n14763 0.114
R11728 GND.n14752 GND.n14750 0.114
R11729 GND.n6327 GND.n6319 0.114
R11730 GND.n6315 GND.n6307 0.114
R11731 GND.n6303 GND.n6295 0.114
R11732 GND.n6291 GND.n6283 0.114
R11733 GND.n6279 GND.n6271 0.114
R11734 GND.n6267 GND.n6259 0.114
R11735 GND.n6225 GND.n6223 0.114
R11736 GND.n6213 GND.n6211 0.114
R11737 GND.n6201 GND.n6199 0.114
R11738 GND.n6189 GND.n6187 0.114
R11739 GND.n6176 GND.n6174 0.114
R11740 GND.n12697 GND.n12689 0.114
R11741 GND.n12685 GND.n12676 0.114
R11742 GND.n12672 GND.n12664 0.114
R11743 GND.n12660 GND.n12651 0.114
R11744 GND.n12647 GND.n12639 0.114
R11745 GND.n12603 GND.n12601 0.114
R11746 GND.n12590 GND.n12588 0.114
R11747 GND.n12578 GND.n12576 0.114
R11748 GND.n12565 GND.n12563 0.114
R11749 GND.n12553 GND.n12551 0.114
R11750 GND.n11308 GND.n11300 0.114
R11751 GND.n11296 GND.n11288 0.114
R11752 GND.n11284 GND.n11276 0.114
R11753 GND.n11272 GND.n11264 0.114
R11754 GND.n11260 GND.n11252 0.114
R11755 GND.n11218 GND.n11216 0.114
R11756 GND.n11206 GND.n11204 0.114
R11757 GND.n11194 GND.n11192 0.114
R11758 GND.n11182 GND.n11180 0.114
R11759 GND.n11170 GND.n11168 0.114
R11760 GND.n11158 GND.n11156 0.114
R11761 GND.n13715 GND.n13707 0.114
R11762 GND.n13703 GND.n13695 0.114
R11763 GND.n13691 GND.n13683 0.114
R11764 GND.n13679 GND.n13671 0.114
R11765 GND.n13667 GND.n13659 0.114
R11766 GND.n13625 GND.n13623 0.114
R11767 GND.n13613 GND.n13611 0.114
R11768 GND.n13601 GND.n13599 0.114
R11769 GND.n13589 GND.n13587 0.114
R11770 GND.n13577 GND.n13575 0.114
R11771 GND.n13565 GND.n13563 0.114
R11772 GND.n13360 GND.n13358 0.114
R11773 GND.n13372 GND.n13370 0.114
R11774 GND.n13385 GND.n13383 0.114
R11775 GND.n13397 GND.n13395 0.114
R11776 GND.n13442 GND.n13433 0.114
R11777 GND.n13454 GND.n13446 0.114
R11778 GND.n13467 GND.n13458 0.114
R11779 GND.n13479 GND.n13471 0.114
R11780 GND.n13492 GND.n13483 0.114
R11781 GND.n13504 GND.n13496 0.114
R11782 GND.n12092 GND.n12024 0.114
R11783 GND.n12020 GND.n12012 0.114
R11784 GND.n12008 GND.n11999 0.114
R11785 GND.n11995 GND.n11987 0.114
R11786 GND.n11983 GND.n11974 0.114
R11787 GND.n11952 GND.n11950 0.114
R11788 GND.n11948 GND.n11946 0.114
R11789 GND.n11943 GND.n11941 0.114
R11790 GND.n11938 GND.n11936 0.114
R11791 GND.n11933 GND.n11931 0.114
R11792 GND.n11928 GND.n11926 0.114
R11793 GND.n11908 GND.n11907 0.114
R11794 GND.n11903 GND.n11902 0.114
R11795 GND.n11898 GND.n11897 0.114
R11796 GND.n11894 GND.n11893 0.114
R11797 GND.n11890 GND.n11889 0.114
R11798 GND.n11886 GND.n11885 0.114
R11799 GND.n11867 GND.n11865 0.114
R11800 GND.n11855 GND.n11853 0.114
R11801 GND.n11843 GND.n11841 0.114
R11802 GND.n11830 GND.n11828 0.114
R11803 GND.n11818 GND.n11816 0.114
R11804 GND.n12198 GND.n12196 0.114
R11805 GND.n12210 GND.n12208 0.114
R11806 GND.n12223 GND.n12221 0.114
R11807 GND.n12235 GND.n12233 0.114
R11808 GND.n12248 GND.n12246 0.114
R11809 GND.n12271 GND.n12270 0.114
R11810 GND.n12275 GND.n12274 0.114
R11811 GND.n12280 GND.n12279 0.114
R11812 GND.n12285 GND.n12284 0.114
R11813 GND.n12290 GND.n12289 0.114
R11814 GND.n12295 GND.n12294 0.114
R11815 GND.n12315 GND.n12313 0.114
R11816 GND.n12320 GND.n12318 0.114
R11817 GND.n12325 GND.n12323 0.114
R11818 GND.n12329 GND.n12327 0.114
R11819 GND.n12333 GND.n12331 0.114
R11820 GND.n12337 GND.n12335 0.114
R11821 GND.n12364 GND.n12356 0.114
R11822 GND.n12377 GND.n12368 0.114
R11823 GND.n12389 GND.n12381 0.114
R11824 GND.n12402 GND.n12393 0.114
R11825 GND.n12476 GND.n12406 0.114
R11826 GND.n13191 GND.n13128 0.114
R11827 GND.n13124 GND.n13116 0.114
R11828 GND.n13112 GND.n13104 0.114
R11829 GND.n13100 GND.n13092 0.114
R11830 GND.n13088 GND.n13080 0.114
R11831 GND.n13058 GND.n13056 0.114
R11832 GND.n13053 GND.n13051 0.114
R11833 GND.n13048 GND.n13046 0.114
R11834 GND.n13043 GND.n13041 0.114
R11835 GND.n13038 GND.n13036 0.114
R11836 GND.n13033 GND.n13031 0.114
R11837 GND.n13013 GND.n13012 0.114
R11838 GND.n13008 GND.n13007 0.114
R11839 GND.n13003 GND.n13002 0.114
R11840 GND.n12999 GND.n12998 0.114
R11841 GND.n12995 GND.n12994 0.114
R11842 GND.n12991 GND.n12990 0.114
R11843 GND.n12971 GND.n12969 0.114
R11844 GND.n12959 GND.n12957 0.114
R11845 GND.n12946 GND.n12944 0.114
R11846 GND.n12934 GND.n12932 0.114
R11847 GND.n12921 GND.n12919 0.114
R11848 GND.n7688 GND.n7686 0.114
R11849 GND.n7700 GND.n7698 0.114
R11850 GND.n7712 GND.n7710 0.114
R11851 GND.n7724 GND.n7722 0.114
R11852 GND.n7736 GND.n7734 0.114
R11853 GND.n7759 GND.n7758 0.114
R11854 GND.n7764 GND.n7763 0.114
R11855 GND.n7769 GND.n7768 0.114
R11856 GND.n7774 GND.n7773 0.114
R11857 GND.n7779 GND.n7778 0.114
R11858 GND.n7784 GND.n7783 0.114
R11859 GND.n7804 GND.n7802 0.114
R11860 GND.n7809 GND.n7807 0.114
R11861 GND.n7814 GND.n7812 0.114
R11862 GND.n7818 GND.n7816 0.114
R11863 GND.n7822 GND.n7820 0.114
R11864 GND.n7826 GND.n7824 0.114
R11865 GND.n7852 GND.n7844 0.114
R11866 GND.n7864 GND.n7856 0.114
R11867 GND.n7877 GND.n7868 0.114
R11868 GND.n7889 GND.n7881 0.114
R11869 GND.n7959 GND.n7893 0.114
R11870 GND.n8145 GND.n8137 0.114
R11871 GND.n8133 GND.n8124 0.114
R11872 GND.n8120 GND.n8112 0.114
R11873 GND.n8108 GND.n8099 0.114
R11874 GND.n8095 GND.n8087 0.114
R11875 GND.n8083 GND.n8074 0.114
R11876 GND.n8038 GND.n8036 0.114
R11877 GND.n8026 GND.n8024 0.114
R11878 GND.n8013 GND.n8011 0.114
R11879 GND.n8001 GND.n7999 0.114
R11880 GND.n7988 GND.n7986 0.114
R11881 GND.n6997 GND.n6995 0.114
R11882 GND.n7010 GND.n7008 0.114
R11883 GND.n7022 GND.n7020 0.114
R11884 GND.n7035 GND.n7033 0.114
R11885 GND.n7047 GND.n7045 0.114
R11886 GND.n7092 GND.n7083 0.114
R11887 GND.n7104 GND.n7096 0.114
R11888 GND.n7117 GND.n7108 0.114
R11889 GND.n7129 GND.n7121 0.114
R11890 GND.n7142 GND.n7133 0.114
R11891 GND.n7155 GND.n7146 0.114
R11892 GND.n7371 GND.n7363 0.114
R11893 GND.n7359 GND.n7351 0.114
R11894 GND.n7347 GND.n7338 0.114
R11895 GND.n7334 GND.n7326 0.114
R11896 GND.n7322 GND.n7313 0.114
R11897 GND.n7277 GND.n7275 0.114
R11898 GND.n7265 GND.n7263 0.114
R11899 GND.n7252 GND.n7250 0.114
R11900 GND.n7240 GND.n7238 0.114
R11901 GND.n7227 GND.n7225 0.114
R11902 GND.n7215 GND.n7213 0.114
R11903 GND.n15941 GND.n15939 0.114
R11904 GND.n15953 GND.n15951 0.114
R11905 GND.n15966 GND.n15964 0.114
R11906 GND.n15978 GND.n15976 0.114
R11907 GND.n15991 GND.n15989 0.114
R11908 GND.n16021 GND.n16017 0.114
R11909 GND.n16029 GND.n16025 0.114
R11910 GND.n16037 GND.n16033 0.114
R11911 GND.n16045 GND.n16041 0.114
R11912 GND.n16053 GND.n16049 0.114
R11913 GND.n16061 GND.n16057 0.114
R11914 GND.n16072 GND.n16070 0.114
R11915 GND.n16077 GND.n16075 0.114
R11916 GND.n16082 GND.n16080 0.114
R11917 GND.n16086 GND.n16084 0.114
R11918 GND.n16089 GND.n16088 0.114
R11919 GND.n16126 GND.n16118 0.114
R11920 GND.n16138 GND.n16130 0.114
R11921 GND.n16150 GND.n16142 0.114
R11922 GND.n16162 GND.n16154 0.114
R11923 GND.n16175 GND.n16166 0.114
R11924 GND.n16228 GND.n16179 0.114
R11925 GND.n1168 GND.n1127 0.114
R11926 GND.n1123 GND.n1115 0.114
R11927 GND.n1111 GND.n1103 0.114
R11928 GND.n1099 GND.n1091 0.114
R11929 GND.n1087 GND.n1079 0.114
R11930 GND.n1053 GND.n1051 0.114
R11931 GND.n1045 GND.n1043 0.114
R11932 GND.n1037 GND.n1035 0.114
R11933 GND.n1029 GND.n1027 0.114
R11934 GND.n1021 GND.n1019 0.114
R11935 GND.n1013 GND.n1011 0.114
R11936 GND.n999 GND.n998 0.114
R11937 GND.n994 GND.n993 0.114
R11938 GND.n989 GND.n988 0.114
R11939 GND.n985 GND.n984 0.114
R11940 GND.n981 GND.n980 0.114
R11941 GND.n951 GND.n949 0.114
R11942 GND.n938 GND.n936 0.114
R11943 GND.n926 GND.n924 0.114
R11944 GND.n913 GND.n911 0.114
R11945 GND.n901 GND.n899 0.114
R11946 GND.n888 GND.n886 0.114
R11947 GND.n9641 GND.n9639 0.114
R11948 GND.n9653 GND.n9651 0.114
R11949 GND.n9666 GND.n9664 0.114
R11950 GND.n9678 GND.n9676 0.114
R11951 GND.n9691 GND.n9689 0.114
R11952 GND.n9721 GND.n9717 0.114
R11953 GND.n9729 GND.n9725 0.114
R11954 GND.n9737 GND.n9733 0.114
R11955 GND.n9745 GND.n9741 0.114
R11956 GND.n9753 GND.n9749 0.114
R11957 GND.n9761 GND.n9757 0.114
R11958 GND.n9772 GND.n9770 0.114
R11959 GND.n9777 GND.n9775 0.114
R11960 GND.n9782 GND.n9780 0.114
R11961 GND.n9786 GND.n9784 0.114
R11962 GND.n9789 GND.n9788 0.114
R11963 GND.n9826 GND.n9818 0.114
R11964 GND.n9838 GND.n9830 0.114
R11965 GND.n9850 GND.n9842 0.114
R11966 GND.n9862 GND.n9854 0.114
R11967 GND.n9875 GND.n9866 0.114
R11968 GND.n9928 GND.n9879 0.114
R11969 GND.n1233 GND.n1231 0.114
R11970 GND.n1245 GND.n1243 0.114
R11971 GND.n1257 GND.n1255 0.114
R11972 GND.n1269 GND.n1267 0.114
R11973 GND.n1281 GND.n1279 0.114
R11974 GND.n1311 GND.n1307 0.114
R11975 GND.n1319 GND.n1315 0.114
R11976 GND.n1327 GND.n1323 0.114
R11977 GND.n1335 GND.n1331 0.114
R11978 GND.n1343 GND.n1339 0.114
R11979 GND.n1351 GND.n1347 0.114
R11980 GND.n1362 GND.n1360 0.114
R11981 GND.n1367 GND.n1365 0.114
R11982 GND.n1372 GND.n1370 0.114
R11983 GND.n1376 GND.n1374 0.114
R11984 GND.n1379 GND.n1378 0.114
R11985 GND.n1418 GND.n1409 0.114
R11986 GND.n1430 GND.n1422 0.114
R11987 GND.n1443 GND.n1434 0.114
R11988 GND.n1455 GND.n1447 0.114
R11989 GND.n1468 GND.n1459 0.114
R11990 GND.n1524 GND.n1472 0.114
R11991 GND.n10305 GND.n10297 0.114
R11992 GND.n10293 GND.n10285 0.114
R11993 GND.n10281 GND.n10272 0.114
R11994 GND.n10268 GND.n10260 0.114
R11995 GND.n10256 GND.n10247 0.114
R11996 GND.n10211 GND.n10209 0.114
R11997 GND.n10199 GND.n10197 0.114
R11998 GND.n10186 GND.n10184 0.114
R11999 GND.n10174 GND.n10172 0.114
R12000 GND.n10161 GND.n10159 0.114
R12001 GND.n10149 GND.n10147 0.114
R12002 GND.n8868 GND.n8860 0.114
R12003 GND.n8856 GND.n8848 0.114
R12004 GND.n8844 GND.n8836 0.114
R12005 GND.n8832 GND.n8824 0.114
R12006 GND.n8820 GND.n8812 0.114
R12007 GND.n8778 GND.n8776 0.114
R12008 GND.n8766 GND.n8764 0.114
R12009 GND.n8754 GND.n8752 0.114
R12010 GND.n8742 GND.n8740 0.114
R12011 GND.n8730 GND.n8728 0.114
R12012 GND.n8718 GND.n8716 0.114
R12013 GND.n8575 GND.n8567 0.114
R12014 GND.n8563 GND.n8555 0.114
R12015 GND.n8551 GND.n8542 0.114
R12016 GND.n8538 GND.n8530 0.114
R12017 GND.n8526 GND.n8517 0.114
R12018 GND.n8481 GND.n8479 0.114
R12019 GND.n8469 GND.n8467 0.114
R12020 GND.n8456 GND.n8454 0.114
R12021 GND.n8444 GND.n8442 0.114
R12022 GND.n8431 GND.n8429 0.114
R12023 GND.n8419 GND.n8417 0.114
R12024 GND.n10129 GND.n10121 0.114
R12025 GND.n10117 GND.n10109 0.114
R12026 GND.n10105 GND.n10097 0.114
R12027 GND.n10093 GND.n10085 0.114
R12028 GND.n10081 GND.n10073 0.114
R12029 GND.n10039 GND.n10037 0.114
R12030 GND.n10027 GND.n10025 0.114
R12031 GND.n10015 GND.n10013 0.114
R12032 GND.n10003 GND.n10001 0.114
R12033 GND.n9991 GND.n9989 0.114
R12034 GND.n9978 GND.n9976 0.114
R12035 GND.n8940 GND.n8938 0.114
R12036 GND.n8952 GND.n8950 0.114
R12037 GND.n8965 GND.n8963 0.114
R12038 GND.n8977 GND.n8975 0.114
R12039 GND.n8990 GND.n8988 0.114
R12040 GND.n9020 GND.n9016 0.114
R12041 GND.n9028 GND.n9024 0.114
R12042 GND.n9036 GND.n9032 0.114
R12043 GND.n9044 GND.n9040 0.114
R12044 GND.n9052 GND.n9048 0.114
R12045 GND.n9060 GND.n9056 0.114
R12046 GND.n9071 GND.n9069 0.114
R12047 GND.n9076 GND.n9074 0.114
R12048 GND.n9081 GND.n9079 0.114
R12049 GND.n9085 GND.n9083 0.114
R12050 GND.n9088 GND.n9087 0.114
R12051 GND.n9125 GND.n9117 0.114
R12052 GND.n9137 GND.n9129 0.114
R12053 GND.n9149 GND.n9141 0.114
R12054 GND.n9161 GND.n9153 0.114
R12055 GND.n9174 GND.n9165 0.114
R12056 GND.n9227 GND.n9178 0.114
R12057 GND.n4534 GND.n4489 0.114
R12058 GND.n4485 GND.n4477 0.114
R12059 GND.n4473 GND.n4464 0.114
R12060 GND.n4460 GND.n4452 0.114
R12061 GND.n4448 GND.n4439 0.114
R12062 GND.n4413 GND.n4411 0.114
R12063 GND.n4405 GND.n4403 0.114
R12064 GND.n4397 GND.n4395 0.114
R12065 GND.n4389 GND.n4387 0.114
R12066 GND.n4381 GND.n4379 0.114
R12067 GND.n4373 GND.n4371 0.114
R12068 GND.n4359 GND.n4358 0.114
R12069 GND.n4354 GND.n4353 0.114
R12070 GND.n4349 GND.n4348 0.114
R12071 GND.n4345 GND.n4344 0.114
R12072 GND.n4341 GND.n4340 0.114
R12073 GND.n4311 GND.n4309 0.114
R12074 GND.n4298 GND.n4296 0.114
R12075 GND.n4286 GND.n4284 0.114
R12076 GND.n4273 GND.n4271 0.114
R12077 GND.n4261 GND.n4259 0.114
R12078 GND.n4248 GND.n4246 0.114
R12079 GND.n3193 GND.n3191 0.114
R12080 GND.n3205 GND.n3203 0.114
R12081 GND.n3217 GND.n3215 0.114
R12082 GND.n3229 GND.n3227 0.114
R12083 GND.n3241 GND.n3239 0.114
R12084 GND.n3283 GND.n3275 0.114
R12085 GND.n3295 GND.n3287 0.114
R12086 GND.n3307 GND.n3299 0.114
R12087 GND.n3319 GND.n3311 0.114
R12088 GND.n3332 GND.n3323 0.114
R12089 GND.n3345 GND.n3336 0.114
R12090 GND.n5093 GND.n5085 0.114
R12091 GND.n5081 GND.n5072 0.114
R12092 GND.n5068 GND.n5060 0.114
R12093 GND.n5056 GND.n5047 0.114
R12094 GND.n5043 GND.n5035 0.114
R12095 GND.n4999 GND.n4997 0.114
R12096 GND.n4986 GND.n4984 0.114
R12097 GND.n4974 GND.n4972 0.114
R12098 GND.n4961 GND.n4959 0.114
R12099 GND.n4949 GND.n4947 0.114
R12100 GND.n4936 GND.n4934 0.114
R12101 GND.n4747 GND.n4739 0.114
R12102 GND.n4735 GND.n4726 0.114
R12103 GND.n4722 GND.n4714 0.114
R12104 GND.n4710 GND.n4701 0.114
R12105 GND.n4697 GND.n4689 0.114
R12106 GND.n4653 GND.n4651 0.114
R12107 GND.n4640 GND.n4638 0.114
R12108 GND.n4628 GND.n4626 0.114
R12109 GND.n4615 GND.n4613 0.114
R12110 GND.n4603 GND.n4601 0.114
R12111 GND.n4590 GND.n4588 0.114
R12112 GND.n2993 GND.n2991 0.114
R12113 GND.n3005 GND.n3003 0.114
R12114 GND.n3017 GND.n3015 0.114
R12115 GND.n3029 GND.n3027 0.114
R12116 GND.n3041 GND.n3039 0.114
R12117 GND.n3083 GND.n3075 0.114
R12118 GND.n3095 GND.n3087 0.114
R12119 GND.n3107 GND.n3099 0.114
R12120 GND.n3119 GND.n3111 0.114
R12121 GND.n3132 GND.n3123 0.114
R12122 GND.n3144 GND.n3136 0.114
R12123 GND.n10417 GND.n10415 0.114
R12124 GND.n10429 GND.n10427 0.114
R12125 GND.n10441 GND.n10439 0.114
R12126 GND.n10453 GND.n10451 0.114
R12127 GND.n10465 GND.n10463 0.114
R12128 GND.n10507 GND.n10499 0.114
R12129 GND.n10519 GND.n10511 0.114
R12130 GND.n10531 GND.n10523 0.114
R12131 GND.n10543 GND.n10535 0.114
R12132 GND.n10555 GND.n10547 0.114
R12133 GND.n10568 GND.n10559 0.114
R12134 GND.n15559 GND.n15557 0.114
R12135 GND.n15572 GND.n15570 0.114
R12136 GND.n15584 GND.n15582 0.114
R12137 GND.n15597 GND.n15595 0.114
R12138 GND.n15609 GND.n15607 0.114
R12139 GND.n15654 GND.n15645 0.114
R12140 GND.n15666 GND.n15658 0.114
R12141 GND.n15679 GND.n15670 0.114
R12142 GND.n15691 GND.n15683 0.114
R12143 GND.n15704 GND.n15695 0.114
R12144 GND.n15136 GND.n15134 0.114
R12145 GND.n15148 GND.n15146 0.114
R12146 GND.n15160 GND.n15158 0.114
R12147 GND.n15172 GND.n15170 0.114
R12148 GND.n15214 GND.n15206 0.114
R12149 GND.n15226 GND.n15218 0.114
R12150 GND.n15238 GND.n15230 0.114
R12151 GND.n15251 GND.n15242 0.114
R12152 GND.n15263 GND.n15255 0.114
R12153 GND.n15275 GND.n15267 0.114
R12154 GND.n3949 GND.n3908 0.114
R12155 GND.n3904 GND.n3896 0.114
R12156 GND.n3892 GND.n3884 0.114
R12157 GND.n3880 GND.n3872 0.114
R12158 GND.n3868 GND.n3860 0.114
R12159 GND.n3834 GND.n3832 0.114
R12160 GND.n3826 GND.n3824 0.114
R12161 GND.n3818 GND.n3816 0.114
R12162 GND.n3810 GND.n3808 0.114
R12163 GND.n3802 GND.n3800 0.114
R12164 GND.n3794 GND.n3792 0.114
R12165 GND.n3780 GND.n3779 0.114
R12166 GND.n3775 GND.n3774 0.114
R12167 GND.n3770 GND.n3769 0.114
R12168 GND.n3766 GND.n3765 0.114
R12169 GND.n3762 GND.n3761 0.114
R12170 GND.n3733 GND.n3731 0.114
R12171 GND.n3721 GND.n3719 0.114
R12172 GND.n3709 GND.n3707 0.114
R12173 GND.n3697 GND.n3695 0.114
R12174 GND.n3685 GND.n3683 0.114
R12175 GND.n3672 GND.n3670 0.114
R12176 GND.n5787 GND.n5746 0.114
R12177 GND.n5742 GND.n5734 0.114
R12178 GND.n5730 GND.n5722 0.114
R12179 GND.n5718 GND.n5710 0.114
R12180 GND.n5706 GND.n5698 0.114
R12181 GND.n5672 GND.n5670 0.114
R12182 GND.n5664 GND.n5662 0.114
R12183 GND.n5656 GND.n5654 0.114
R12184 GND.n5648 GND.n5646 0.114
R12185 GND.n5640 GND.n5638 0.114
R12186 GND.n5632 GND.n5630 0.114
R12187 GND.n5618 GND.n5617 0.114
R12188 GND.n5613 GND.n5612 0.114
R12189 GND.n5608 GND.n5607 0.114
R12190 GND.n5604 GND.n5603 0.114
R12191 GND.n5600 GND.n5599 0.114
R12192 GND.n5570 GND.n5568 0.114
R12193 GND.n5557 GND.n5555 0.114
R12194 GND.n5545 GND.n5543 0.114
R12195 GND.n5532 GND.n5530 0.114
R12196 GND.n5520 GND.n5518 0.114
R12197 GND.n5507 GND.n5505 0.114
R12198 GND.n7595 GND.n7592 0.113
R12199 GND.n7972 GND.n7967 0.113
R12200 GND.n9962 GND.n9957 0.113
R12201 GND.n13517 GND.n13515 0.11
R12202 GND.n13545 GND.n13544 0.11
R12203 GND.n8158 GND.n8156 0.11
R12204 GND.n7198 GND.n7197 0.11
R12205 GND.n7170 GND.n7168 0.11
R12206 GND.n3178 GND.n3177 0.11
R12207 GND.n2672 GND.n2671 0.11
R12208 GND.n4921 GND.n4920 0.11
R12209 GND.n15757 GND.n15752 0.11
R12210 GND.n15725 GND.n15723 0.11
R12211 GND.n15446 GND.n15444 0.11
R12212 GND.n7423 GND.n7422 0.11
R12213 GND.n8374 GND.n8373 0.11
R12214 GND.n9256 GND.n9255 0.11
R12215 GND.n8391 GND.n8388 0.11
R12216 GND.n7619 GND.n7595 0.109
R12217 GND.n7967 GND.n7964 0.109
R12218 GND.n9957 GND.n9954 0.109
R12219 GND.n10334 GND.n10333 0.109
R12220 GND.n4569 GND.n4568 0.106
R12221 GND.n5792 GND.n1910 0.106
R12222 GND.n5449 GND.n5440 0.106
R12223 GND.n5238 GND.n5235 0.106
R12224 GND.n14490 GND.n14489 0.103
R12225 GND.n15448 GND.n15447 0.103
R12226 GND.n15739 GND.n10694 0.103
R12227 GND.n15718 GND.n10715 0.103
R12228 GND.n14119 GND.n14118 0.103
R12229 GND.n4922 GND.n1935 0.103
R12230 GND.n4907 GND.n4904 0.103
R12231 GND.n10783 GND.n10782 0.103
R12232 GND.n13883 GND.n13882 0.103
R12233 GND.n10905 GND.n10904 0.103
R12234 GND.n14001 GND.n10718 0.103
R12235 GND.n12829 GND.n12828 0.103
R12236 GND.n13531 GND.n11653 0.103
R12237 GND.n13510 GND.n11721 0.103
R12238 GND.n13546 GND.n11434 0.103
R12239 GND.n6108 GND.n6106 0.103
R12240 GND.n8369 GND.n8367 0.103
R12241 GND.n8151 GND.n5848 0.103
R12242 GND.n5913 GND.n5912 0.103
R12243 GND.n6523 GND.n6517 0.103
R12244 GND.n7384 GND.n7379 0.103
R12245 GND.n7184 GND.n6826 0.103
R12246 GND.n7199 GND.n6576 0.103
R12247 GND.n7163 GND.n6985 0.103
R12248 GND.n9409 GND.n9408 0.103
R12249 GND.n9278 GND.n1815 0.103
R12250 GND.n1684 GND.n1681 0.103
R12251 GND.n1582 GND.n1581 0.103
R12252 GND.n9245 GND.n1897 0.103
R12253 GND.n5308 GND.n5307 0.103
R12254 GND.n3382 GND.n2608 0.103
R12255 GND.n2477 GND.n2474 0.103
R12256 GND.n3175 GND.n3164 0.103
R12257 GND.n5217 GND.n5216 0.103
R12258 GND.n1960 GND.n1959 0.103
R12259 GND.n15759 GND.n15758 0.103
R12260 GND.n15313 GND.n15312 0.103
R12261 GND.n14728 GND.n14464 0.103
R12262 GND.n15286 GND.n14403 0.103
R12263 GND.n8879 GND.n8878 0.102
R12264 GND.n17684 GND.n17683 0.101
R12265 GND.n4562 GND.n4559 0.1
R12266 GND.n12115 GND.n12114 0.098
R12267 GND.n12498 GND.n12495 0.098
R12268 GND.n830 GND.n829 0.098
R12269 GND.n10375 GND.n10372 0.098
R12270 GND.n14013 GND.n14010 0.097
R12271 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SUBSTRATE GND.n14838
+ 0.096
R12272 GND.n2979 GND.n2839 0.096
R12273 GND.n4559 GND.n4189 0.096
R12274 GND.n6237 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE
+ 0.096
R12275 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE GND.n12626
+ 0.096
R12276 GND.n13410 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE
+ 0.096
R12277 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE GND.n11957
+ 0.096
R12278 GND.n11879 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.096
R12279 GND.n7752 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE
+ 0.096
R12280 GND.n7831 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE
+ 0.096
R12281 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE GND.n7301
+ 0.096
R12282 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE GND.n1062
+ 0.096
R12283 GND.n973 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE
+ 0.096
R12284 GND.n1297 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE
+ 0.096
R12285 GND.n1386 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.096
R12286 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SUBSTRATE GND.n8800
+ 0.096
R12287 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE GND.n8505
+ 0.096
R12288 GND.n3253 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SUBSTRATE
+ 0.096
R12289 GND.n3053 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SUBSTRATE
+ 0.096
R12290 GND.n10477 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SUBSTRATE
+ 0.096
R12291 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SUBSTRATE GND.n3843
+ 0.096
R12292 GND.n3754 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE
+ 0.096
R12293 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE GND.n5681
+ 0.096
R12294 GND.n5592 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE
+ 0.096
R12295 GND.n5362 GND.n5357 0.093
R12296 GND.n5431 GND.n5428 0.089
R12297 GND.n9235 GND.n9232 0.083
R12298 GND.n8889 GND.n8888 0.083
R12299 GND.n12839 GND.n12836 0.08
R12300 GND.n13337 GND.n13204 0.08
R12301 GND.n14737 GND.n14417 0.08
R12302 GND.n15884 GND.n15881 0.08
R12303 GND.n12124 GND.n12123 0.079
R12304 GND.n12489 GND.n12486 0.079
R12305 GND.n9933 GND.n9589 0.079
R12306 GND.n10366 GND.n10363 0.079
R12307 GND.n10632 GND.n10631 0.078
R12308 GND.n15477 GND.n15474 0.078
R12309 GND.n13941 GND.n13938 0.078
R12310 GND.n13813 GND.n13810 0.078
R12311 GND.n13780 GND.n13779 0.078
R12312 GND.n11563 GND.n11560 0.078
R12313 GND.n11055 GND.n11052 0.078
R12314 GND.n11376 GND.n11375 0.078
R12315 GND.n8216 GND.n8215 0.078
R12316 GND.n6764 GND.n6763 0.078
R12317 GND.n7529 GND.n7526 0.078
R12318 GND.n9349 GND.n9348 0.078
R12319 GND.n1754 GND.n1753 0.078
R12320 GND.n8643 GND.n8640 0.078
R12321 GND.n2547 GND.n2546 0.078
R12322 GND.n5156 GND.n5155 0.078
R12323 GND.n4844 GND.n4843 0.078
R12324 GND.n3563 GND.n3560 0.078
R12325 GND.n15373 GND.n15370 0.078
R12326 GND.n14977 GND.n14976 0.078
R12327 GND.n15059 GND.n15056 0.078
R12328 GND.n10764 GND.n10763 0.078
R12329 GND.n12767 GND.n12766 0.078
R12330 GND.n11667 GND.n11664 0.078
R12331 GND.n13268 GND.n13265 0.078
R12332 GND.n8305 GND.n8304 0.078
R12333 GND.n6359 GND.n6353 0.078
R12334 GND.n5977 GND.n5974 0.078
R12335 GND.n6467 GND.n6466 0.078
R12336 GND.n6889 GND.n6886 0.078
R12337 GND.n6654 GND.n6651 0.078
R12338 GND.n7488 GND.n7487 0.078
R12339 GND.n2385 GND.n2384 0.078
R12340 GND.n15818 GND.n15815 0.078
R12341 GND.n9945 GND.n9944 0.077
R12342 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE GND.n13531 0.075
R12343 GND.n5912 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE 0.075
R12344 GND.n7184 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE 0.075
R12345 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/GATE GND.n4907 0.075
R12346 GND.n15739 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/GATE 0.075
R12347 GND.n10669 GND.n10667 0.073
R12348 GND.n14057 GND.n14056 0.073
R12349 GND.n3529 GND.n3528 0.073
R12350 GND.n4880 GND.n4878 0.073
R12351 GND.n10810 GND.n10809 0.073
R12352 GND.n13909 GND.n13908 0.073
R12353 GND.n10929 GND.n10928 0.073
R12354 GND.n10978 GND.n10977 0.073
R12355 GND.n12803 GND.n12801 0.073
R12356 GND.n11471 GND.n11470 0.073
R12357 GND.n11531 GND.n11530 0.073
R12358 GND.n11628 GND.n11626 0.073
R12359 GND.n13233 GND.n13232 0.073
R12360 GND.n11410 GND.n11408 0.073
R12361 GND.n6081 GND.n6079 0.073
R12362 GND.n8342 GND.n8340 0.073
R12363 GND.n6392 GND.n6390 0.073
R12364 GND.n5940 GND.n5939 0.073
R12365 GND.n6495 GND.n6493 0.073
R12366 GND.n6853 GND.n6852 0.073
R12367 GND.n6618 GND.n6617 0.073
R12368 GND.n6801 GND.n6799 0.073
R12369 GND.n6551 GND.n6549 0.073
R12370 GND.n6960 GND.n6958 0.073
R12371 GND.n9384 GND.n9382 0.073
R12372 GND.n1791 GND.n1789 0.073
R12373 GND.n8613 GND.n8612 0.073
R12374 GND.n2583 GND.n2581 0.073
R12375 GND.n2321 GND.n2319 0.073
R12376 GND.n5191 GND.n5189 0.073
R12377 GND.n2875 GND.n2874 0.073
R12378 GND.n15783 GND.n15782 0.073
R12379 GND.n15337 GND.n15336 0.073
R12380 GND.n14440 GND.n14438 0.073
R12381 GND.n15029 GND.n15028 0.073
R12382 GND.n10686 GND.n10685 0.073
R12383 GND.n14043 GND.n14040 0.073
R12384 GND.n3514 GND.n3511 0.073
R12385 GND.n4897 GND.n4896 0.073
R12386 GND.n10794 GND.n10791 0.073
R12387 GND.n13894 GND.n13891 0.073
R12388 GND.n10915 GND.n10912 0.073
R12389 GND.n10964 GND.n10961 0.073
R12390 GND.n12820 GND.n12819 0.073
R12391 GND.n11455 GND.n11452 0.073
R12392 GND.n11516 GND.n11513 0.073
R12393 GND.n11645 GND.n11644 0.073
R12394 GND.n13219 GND.n13216 0.073
R12395 GND.n11427 GND.n11426 0.073
R12396 GND.n6098 GND.n6097 0.073
R12397 GND.n8359 GND.n8358 0.073
R12398 GND.n5841 GND.n5840 0.073
R12399 GND.n5924 GND.n5921 0.073
R12400 GND.n6510 GND.n6509 0.073
R12401 GND.n6837 GND.n6834 0.073
R12402 GND.n6602 GND.n6599 0.073
R12403 GND.n6818 GND.n6817 0.073
R12404 GND.n6568 GND.n6567 0.073
R12405 GND.n6977 GND.n6976 0.073
R12406 GND.n9401 GND.n9400 0.073
R12407 GND.n1808 GND.n1807 0.073
R12408 GND.n8598 GND.n8595 0.073
R12409 GND.n2600 GND.n2599 0.073
R12410 GND.n2309 GND.n2306 0.073
R12411 GND.n5208 GND.n5207 0.073
R12412 GND.n2860 GND.n2857 0.073
R12413 GND.n15769 GND.n15766 0.073
R12414 GND.n15323 GND.n15320 0.073
R12415 GND.n14457 GND.n14456 0.073
R12416 GND.n15015 GND.n15012 0.073
R12417 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE GND.n13869 0.073
R12418 GND.n1697 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE 0.073
R12419 GND.n2490 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/GATE 0.073
R12420 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/GATE GND.n15429 0.073
R12421 GND.n13899 GND.n13898 0.072
R12422 GND.n10969 GND.n10968 0.072
R12423 GND.n11521 GND.n11520 0.072
R12424 GND.n11420 GND.n11418 0.072
R12425 GND.n8603 GND.n8602 0.072
R12426 GND.n5201 GND.n5199 0.072
R12427 GND.n2593 GND.n2591 0.072
R12428 GND.n2329 GND.n2313 0.072
R12429 GND.n2865 GND.n2864 0.072
R12430 GND.n14450 GND.n14448 0.072
R12431 GND.n2296 GND.n2295 0.072
R12432 GND.n10679 GND.n10677 0.072
R12433 GND.n14048 GND.n14047 0.072
R12434 GND.n3519 GND.n3518 0.072
R12435 GND.n4890 GND.n4888 0.072
R12436 GND.n10800 GND.n10799 0.072
R12437 GND.n10920 GND.n10919 0.072
R12438 GND.n12813 GND.n12811 0.072
R12439 GND.n11461 GND.n11460 0.072
R12440 GND.n11638 GND.n11636 0.072
R12441 GND.n13224 GND.n13223 0.072
R12442 GND.n6091 GND.n6089 0.072
R12443 GND.n8352 GND.n8350 0.072
R12444 GND.n6401 GND.n6400 0.072
R12445 GND.n5930 GND.n5929 0.072
R12446 GND.n6504 GND.n6502 0.072
R12447 GND.n6843 GND.n6842 0.072
R12448 GND.n6608 GND.n6607 0.072
R12449 GND.n6811 GND.n6809 0.072
R12450 GND.n6561 GND.n6559 0.072
R12451 GND.n6970 GND.n6968 0.072
R12452 GND.n9394 GND.n9392 0.072
R12453 GND.n1801 GND.n1799 0.072
R12454 GND.n15774 GND.n15773 0.072
R12455 GND.n15328 GND.n15327 0.072
R12456 GND.n15020 GND.n15019 0.072
R12457 GND.n6383 GND.n6366 0.071
R12458 GND.n5968 GND.n5962 0.071
R12459 GND.n6473 GND.n6472 0.071
R12460 GND.n6880 GND.n6875 0.071
R12461 GND.n6645 GND.n6640 0.071
R12462 GND.n16454 GND.n16452 0.071
R12463 GND.n16715 GND.n16713 0.071
R12464 GND.n16976 GND.n16974 0.071
R12465 GND.n17237 GND.n17235 0.071
R12466 GND.n17498 GND.n17496 0.071
R12467 GND.n10659 GND.n10657 0.068
R12468 GND.n14067 GND.n14066 0.068
R12469 GND.n3539 GND.n3538 0.068
R12470 GND.n4870 GND.n4868 0.068
R12471 GND.n10820 GND.n10819 0.068
R12472 GND.n13919 GND.n13918 0.068
R12473 GND.n10939 GND.n10938 0.068
R12474 GND.n10988 GND.n10987 0.068
R12475 GND.n12793 GND.n12791 0.068
R12476 GND.n11481 GND.n11480 0.068
R12477 GND.n11541 GND.n11540 0.068
R12478 GND.n13243 GND.n13242 0.068
R12479 GND.n11400 GND.n11398 0.068
R12480 GND.n6071 GND.n6069 0.068
R12481 GND.n8332 GND.n8330 0.068
R12482 GND.n6371 GND.n6370 0.068
R12483 GND.n5950 GND.n5949 0.068
R12484 GND.n6486 GND.n6484 0.068
R12485 GND.n6863 GND.n6862 0.068
R12486 GND.n6628 GND.n6627 0.068
R12487 GND.n6791 GND.n6789 0.068
R12488 GND.n6541 GND.n6539 0.068
R12489 GND.n6950 GND.n6948 0.068
R12490 GND.n9374 GND.n9372 0.068
R12491 GND.n1781 GND.n1779 0.068
R12492 GND.n8623 GND.n8622 0.068
R12493 GND.n2573 GND.n2571 0.068
R12494 GND.n2281 GND.n2280 0.068
R12495 GND.n5181 GND.n5179 0.068
R12496 GND.n2885 GND.n2884 0.068
R12497 GND.n15793 GND.n15792 0.068
R12498 GND.n15347 GND.n15346 0.068
R12499 GND.n14430 GND.n14428 0.068
R12500 GND.n15039 GND.n15038 0.068
R12501 GND.n16467 GND.n16465 0.068
R12502 GND.n16542 GND.n16541 0.068
R12503 GND.n16367 GND.n16366 0.068
R12504 GND.n16728 GND.n16726 0.068
R12505 GND.n16803 GND.n16802 0.068
R12506 GND.n16628 GND.n16627 0.068
R12507 GND.n16989 GND.n16987 0.068
R12508 GND.n17064 GND.n17063 0.068
R12509 GND.n16889 GND.n16888 0.068
R12510 GND.n17250 GND.n17248 0.068
R12511 GND.n17325 GND.n17324 0.068
R12512 GND.n17150 GND.n17149 0.068
R12513 GND.n17511 GND.n17509 0.068
R12514 GND.n17586 GND.n17585 0.068
R12515 GND.n17411 GND.n17410 0.068
R12516 GND.n655 GND.n654 0.068
R12517 GND.n758 GND.n757 0.068
R12518 GND.n590 GND.n589 0.068
R12519 GND.n397 GND.n396 0.068
R12520 GND.n500 GND.n499 0.068
R12521 GND.n332 GND.n331 0.068
R12522 GND.n139 GND.n138 0.068
R12523 GND.n242 GND.n241 0.068
R12524 GND.n74 GND.n73 0.068
R12525 GND.n17754 GND.n17753 0.068
R12526 GND.n17831 GND.n17830 0.068
R12527 GND.n17910 GND.n17909 0.068
R12528 GND.n17616 GND.n17615 0.068
R12529 GND.n17449 GND.n17448 0.068
R12530 GND.n17355 GND.n17354 0.068
R12531 GND.n17188 GND.n17187 0.068
R12532 GND.n17094 GND.n17093 0.068
R12533 GND.n16927 GND.n16926 0.068
R12534 GND.n16833 GND.n16832 0.068
R12535 GND.n16666 GND.n16665 0.068
R12536 GND.n16572 GND.n16571 0.068
R12537 GND.n16405 GND.n16404 0.068
R12538 GND.n10 GND.n9 0.068
R12539 GND.n17701 GND.n17700 0.068
R12540 GND.n274 GND.n273 0.068
R12541 GND.n110 GND.n109 0.068
R12542 GND.n532 GND.n531 0.068
R12543 GND.n368 GND.n367 0.068
R12544 GND.n790 GND.n789 0.068
R12545 GND.n626 GND.n625 0.068
R12546 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE GND.n11240
+ 0.068
R12547 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE GND.n13647
+ 0.068
R12548 GND.n12264 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE
+ 0.068
R12549 GND.n12342 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE
+ 0.068
R12550 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE GND.n13063
+ 0.068
R12551 GND.n12984 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.068
R12552 GND.n8051 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE
+ 0.068
R12553 GND.n7060 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE
+ 0.068
R12554 GND.n16007 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE
+ 0.068
R12555 GND.n16096 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE
+ 0.068
R12556 GND.n9707 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE
+ 0.068
R12557 GND.n9796 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.068
R12558 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SUBSTRATE GND.n10235
+ 0.068
R12559 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE GND.n10061
+ 0.068
R12560 GND.n9006 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE
+ 0.068
R12561 GND.n9095 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE
+ 0.068
R12562 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SUBSTRATE GND.n4422
+ 0.068
R12563 GND.n4333 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE
+ 0.068
R12564 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SUBSTRATE GND.n5022
+ 0.068
R12565 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SUBSTRATE GND.n4676
+ 0.068
R12566 GND.n15622 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SUBSTRATE
+ 0.068
R12567 GND.n15184 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SUBSTRATE
+ 0.068
R12568 GND.n17670 GND.n17669 0.065
R12569 GND.n644 GND.n643 0.065
R12570 GND.n746 GND.n745 0.065
R12571 GND.n578 GND.n577 0.065
R12572 GND.n386 GND.n385 0.065
R12573 GND.n488 GND.n487 0.065
R12574 GND.n320 GND.n319 0.065
R12575 GND.n128 GND.n127 0.065
R12576 GND.n230 GND.n229 0.065
R12577 GND.n62 GND.n61 0.065
R12578 GND.n17743 GND.n17742 0.065
R12579 GND.n17819 GND.n17818 0.065
R12580 GND.n17898 GND.n17897 0.065
R12581 GND.n16479 GND.n16477 0.064
R12582 GND.n16514 GND.n16512 0.064
R12583 GND.n16356 GND.n16355 0.064
R12584 GND.n16740 GND.n16738 0.064
R12585 GND.n16775 GND.n16773 0.064
R12586 GND.n16617 GND.n16616 0.064
R12587 GND.n17001 GND.n16999 0.064
R12588 GND.n17036 GND.n17034 0.064
R12589 GND.n16878 GND.n16877 0.064
R12590 GND.n17262 GND.n17260 0.064
R12591 GND.n17297 GND.n17295 0.064
R12592 GND.n17139 GND.n17138 0.064
R12593 GND.n17523 GND.n17521 0.064
R12594 GND.n17558 GND.n17556 0.064
R12595 GND.n17400 GND.n17399 0.064
R12596 GND.n14499 GND.n14498 0.06
R12597 GND.n14524 GND.n14523 0.06
R12598 GND.n14515 GND.n14513 0.06
R12599 GND.n14636 GND.n14476 0.06
R12600 GND.n14548 GND.n14547 0.06
R12601 GND.n14559 GND.n14558 0.06
R12602 GND.n14570 GND.n14569 0.06
R12603 GND.n14128 GND.n14127 0.06
R12604 GND.n14137 GND.n14136 0.06
R12605 GND.n14148 GND.n14147 0.06
R12606 GND.n14292 GND.n14158 0.06
R12607 GND.n14170 GND.n14169 0.06
R12608 GND.n14190 GND.n14189 0.06
R12609 GND.n14201 GND.n14200 0.06
R12610 GND.n14291 GND.n14211 0.06
R12611 GND.n12124 GND.n11744 0.06
R12612 GND.n12486 GND.n12485 0.06
R12613 GND.n9938 GND.n9933 0.06
R12614 GND.n1674 GND.n1673 0.06
R12615 GND.n1665 GND.n1664 0.06
R12616 GND.n1656 GND.n1654 0.06
R12617 GND.n9496 GND.n1636 0.06
R12618 GND.n1591 GND.n1590 0.06
R12619 GND.n1612 GND.n1611 0.06
R12620 GND.n1623 GND.n1622 0.06
R12621 GND.n1634 GND.n1633 0.06
R12622 GND.n2467 GND.n2466 0.06
R12623 GND.n2245 GND.n2244 0.06
R12624 GND.n2256 GND.n2255 0.06
R12625 GND.n3477 GND.n2266 0.06
R12626 GND.n2216 GND.n2215 0.06
R12627 GND.n2227 GND.n2226 0.06
R12628 GND.n2238 GND.n2237 0.06
R12629 GND.n2012 GND.n2011 0.06
R12630 GND.n2032 GND.n2031 0.06
R12631 GND.n2043 GND.n2042 0.06
R12632 GND.n2134 GND.n2053 0.06
R12633 GND.n1969 GND.n1968 0.06
R12634 GND.n1979 GND.n1978 0.06
R12635 GND.n1990 GND.n1989 0.06
R12636 GND.n2135 GND.n2000 0.06
R12637 GND.n10363 GND.n10362 0.06
R12638 GND.n2910 GND.n2907 0.06
R12639 GND.n714 GND.n712 0.06
R12640 GND.n566 GND.n565 0.06
R12641 GND.n688 GND.n686 0.06
R12642 GND.n456 GND.n454 0.06
R12643 GND.n308 GND.n307 0.06
R12644 GND.n430 GND.n428 0.06
R12645 GND.n198 GND.n196 0.06
R12646 GND.n50 GND.n49 0.06
R12647 GND.n172 GND.n170 0.06
R12648 GND.n17708 GND.n17706 0.06
R12649 GND.n17886 GND.n17885 0.06
R12650 GND.n17787 GND.n17785 0.06
R12651 GND.n16488 GND.n16487 0.059
R12652 GND.n16749 GND.n16748 0.059
R12653 GND.n17010 GND.n17009 0.059
R12654 GND.n17271 GND.n17270 0.059
R12655 GND.n17532 GND.n17531 0.059
R12656 GND.n707 GND.n706 0.059
R12657 GND.n449 GND.n448 0.059
R12658 GND.n191 GND.n190 0.059
R12659 GND.n4 GND.n3 0.059
R12660 GND.n10840 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN 0.059
R12661 GND.n11501 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN 0.059
R12662 GND.n8228 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN 0.059
R12663 GND.n6583 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN 0.059
R12664 GND.n13877 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE 0.058
R12665 GND.n9948 GND.n9945 0.058
R12666 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE GND.n1694 0.058
R12667 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/GATE GND.n2487 0.058
R12668 GND.n15437 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/GATE 0.058
R12669 GND.n12835 GND.n12832 0.057
R12670 GND.n14009 GND.n14004 0.057
R12671 GND.n13336 GND.n13333 0.057
R12672 GND.n11318 GND.n11315 0.057
R12673 GND.n3355 GND.n3352 0.057
R12674 GND.n5225 GND.n5220 0.057
R12675 GND.n2978 GND.n2972 0.057
R12676 GND.n4760 GND.n4757 0.057
R12677 GND.n15880 GND.n15875 0.057
R12678 GND.n15544 GND.n15539 0.057
R12679 GND.n14736 GND.n14731 0.057
R12680 GND.n15285 GND.n15282 0.057
R12681 GND.n16436 GND.n16435 0.057
R12682 GND.n16522 GND.n16521 0.057
R12683 GND.n16345 GND.n16344 0.057
R12684 GND.n16697 GND.n16696 0.057
R12685 GND.n16783 GND.n16782 0.057
R12686 GND.n16606 GND.n16605 0.057
R12687 GND.n16958 GND.n16957 0.057
R12688 GND.n17044 GND.n17043 0.057
R12689 GND.n16867 GND.n16866 0.057
R12690 GND.n17219 GND.n17218 0.057
R12691 GND.n17305 GND.n17304 0.057
R12692 GND.n17128 GND.n17127 0.057
R12693 GND.n17480 GND.n17479 0.057
R12694 GND.n17566 GND.n17565 0.057
R12695 GND.n17389 GND.n17388 0.057
R12696 GND.n10803 GND.n10800 0.057
R12697 GND.n10923 GND.n10920 0.057
R12698 GND.n12811 GND.n12810 0.057
R12699 GND.n11464 GND.n11461 0.057
R12700 GND.n11636 GND.n11635 0.057
R12701 GND.n13227 GND.n13224 0.057
R12702 GND.n6089 GND.n6088 0.057
R12703 GND.n8350 GND.n8349 0.057
R12704 GND.n5933 GND.n5930 0.057
R12705 GND.n6401 GND.n6398 0.057
R12706 GND.n6502 GND.n6501 0.057
R12707 GND.n6846 GND.n6843 0.057
R12708 GND.n6611 GND.n6608 0.057
R12709 GND.n6809 GND.n6808 0.057
R12710 GND.n6559 GND.n6558 0.057
R12711 GND.n6968 GND.n6967 0.057
R12712 GND.n1799 GND.n1798 0.057
R12713 GND.n9392 GND.n9391 0.057
R12714 GND.n4888 GND.n4887 0.057
R12715 GND.n3522 GND.n3519 0.057
R12716 GND.n14051 GND.n14048 0.057
R12717 GND.n10677 GND.n10676 0.057
R12718 GND.n15777 GND.n15774 0.057
R12719 GND.n15331 GND.n15328 0.057
R12720 GND.n15023 GND.n15020 0.057
R12721 GND.n13902 GND.n13899 0.057
R12722 GND.n10972 GND.n10969 0.057
R12723 GND.n11524 GND.n11521 0.057
R12724 GND.n11418 GND.n11417 0.057
R12725 GND.n8606 GND.n8603 0.057
R12726 GND.n2591 GND.n2590 0.057
R12727 GND.n2329 GND.n2328 0.057
R12728 GND.n5199 GND.n5198 0.057
R12729 GND.n2868 GND.n2865 0.057
R12730 GND.n14448 GND.n14447 0.057
R12731 GND.n13539 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE 0.056
R12732 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE GND.n5909 0.056
R12733 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE GND.n7181 0.056
R12734 GND.n9232 GND.n1904 0.056
R12735 GND.n4915 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/GATE 0.056
R12736 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/GATE GND.n15736 0.056
R12737 GND.n8889 GND.n5820 0.056
R12738 GND.n10832 GND.n10831 0.055
R12739 GND.n11493 GND.n11492 0.055
R12740 GND.n16392 GND.n16391 0.055
R12741 GND.n16566 GND.n16565 0.055
R12742 GND.n16653 GND.n16652 0.055
R12743 GND.n16827 GND.n16826 0.055
R12744 GND.n16914 GND.n16913 0.055
R12745 GND.n17088 GND.n17087 0.055
R12746 GND.n17175 GND.n17174 0.055
R12747 GND.n17349 GND.n17348 0.055
R12748 GND.n17436 GND.n17435 0.055
R12749 GND.n17610 GND.n17609 0.055
R12750 GND.n613 GND.n612 0.055
R12751 GND.n679 GND.n678 0.055
R12752 GND.n782 GND.n781 0.055
R12753 GND.n355 GND.n354 0.055
R12754 GND.n421 GND.n420 0.055
R12755 GND.n524 GND.n523 0.055
R12756 GND.n97 GND.n96 0.055
R12757 GND.n163 GND.n162 0.055
R12758 GND.n266 GND.n265 0.055
R12759 GND.n17933 GND.n17932 0.055
R12760 GND.n17778 GND.n17777 0.055
R12761 GND.n17855 GND.n17854 0.055
R12762 GND.n10688 GND.n10686 0.054
R12763 GND.n14040 GND.n14039 0.054
R12764 GND.n3511 GND.n3510 0.054
R12765 GND.n4899 GND.n4897 0.054
R12766 GND.n10791 GND.n10790 0.054
R12767 GND.n13891 GND.n13890 0.054
R12768 GND.n10912 GND.n10911 0.054
R12769 GND.n10961 GND.n10960 0.054
R12770 GND.n12822 GND.n12820 0.054
R12771 GND.n11452 GND.n11451 0.054
R12772 GND.n11513 GND.n11512 0.054
R12773 GND.n11647 GND.n11645 0.054
R12774 GND.n13216 GND.n13215 0.054
R12775 GND.n11429 GND.n11427 0.054
R12776 GND.n6100 GND.n6098 0.054
R12777 GND.n8361 GND.n8359 0.054
R12778 GND.n5843 GND.n5841 0.054
R12779 GND.n5921 GND.n5920 0.054
R12780 GND.n6512 GND.n6510 0.054
R12781 GND.n6834 GND.n6833 0.054
R12782 GND.n6599 GND.n6598 0.054
R12783 GND.n6820 GND.n6818 0.054
R12784 GND.n6570 GND.n6568 0.054
R12785 GND.n6979 GND.n6977 0.054
R12786 GND.n9403 GND.n9401 0.054
R12787 GND.n1810 GND.n1808 0.054
R12788 GND.n8595 GND.n8594 0.054
R12789 GND.n2602 GND.n2600 0.054
R12790 GND.n2306 GND.n2305 0.054
R12791 GND.n5210 GND.n5208 0.054
R12792 GND.n2857 GND.n2856 0.054
R12793 GND.n15766 GND.n15765 0.054
R12794 GND.n15320 GND.n15319 0.054
R12795 GND.n14459 GND.n14457 0.054
R12796 GND.n15012 GND.n15011 0.054
R12797 GND.n13799 GND.n10949 0.054
R12798 GND.n12781 GND.n12779 0.054
R12799 GND.n11041 GND.n11028 0.054
R12800 GND.n13254 GND.n13253 0.054
R12801 GND.n8227 GND.n5831 0.054
R12802 GND.n8320 GND.n8318 0.054
R12803 GND.n6779 GND.n6777 0.054
R12804 GND.n7500 GND.n6163 0.054
R12805 GND.n7520 GND.n7519 0.054
R12806 GND.n9362 GND.n9360 0.054
R12807 GND.n1769 GND.n1767 0.054
R12808 GND.n5169 GND.n5167 0.054
R12809 GND.n2561 GND.n2559 0.054
R12810 GND.n4858 GND.n4856 0.054
R12811 GND.n3550 GND.n3549 0.054
R12812 GND.n15464 GND.n14077 0.054
R12813 GND.n10647 GND.n10645 0.054
R12814 GND.n15804 GND.n15803 0.054
R12815 GND.n15358 GND.n15357 0.054
R12816 GND.n15050 GND.n15049 0.054
R12817 GND.n13931 GND.n13930 0.054
R12818 GND.n13932 GND.n13931 0.054
R12819 GND.n13790 GND.n13789 0.054
R12820 GND.n13790 GND.n10998 0.054
R12821 GND.n11553 GND.n11552 0.054
R12822 GND.n11554 GND.n11553 0.054
R12823 GND.n11386 GND.n11385 0.054
R12824 GND.n11388 GND.n11386 0.054
R12825 GND.n8635 GND.n8634 0.054
R12826 GND.n8634 GND.n8633 0.054
R12827 GND.n2902 GND.n2896 0.054
R12828 GND.n2896 GND.n2895 0.054
R12829 GND.n14988 GND.n14987 0.054
R12830 GND.n14988 GND.n14413 0.054
R12831 GND.n10645 GND.n10644 0.054
R12832 GND.n15469 GND.n15464 0.054
R12833 GND.n3555 GND.n3550 0.054
R12834 GND.n4856 GND.n4855 0.054
R12835 GND.n13805 GND.n13799 0.054
R12836 GND.n12779 GND.n12778 0.054
R12837 GND.n11047 GND.n11041 0.054
R12838 GND.n13260 GND.n13254 0.054
R12839 GND.n8227 GND.n8226 0.054
R12840 GND.n8318 GND.n8317 0.054
R12841 GND.n6777 GND.n6776 0.054
R12842 GND.n7500 GND.n7499 0.054
R12843 GND.n7521 GND.n7520 0.054
R12844 GND.n9360 GND.n9359 0.054
R12845 GND.n1767 GND.n1766 0.054
R12846 GND.n2559 GND.n2558 0.054
R12847 GND.n5167 GND.n5166 0.054
R12848 GND.n15810 GND.n15804 0.054
R12849 GND.n15365 GND.n15358 0.054
R12850 GND.n15051 GND.n15050 0.054
R12851 GND.n5229 GND.n5226 0.054
R12852 GND.n4752 GND.n4577 0.054
R12853 GND.n10832 GND.n10769 0.054
R12854 GND.n16566 GND.n16553 0.054
R12855 GND.n16392 GND.n16379 0.054
R12856 GND.n16827 GND.n16814 0.054
R12857 GND.n16653 GND.n16640 0.054
R12858 GND.n17088 GND.n17075 0.054
R12859 GND.n16914 GND.n16901 0.054
R12860 GND.n17349 GND.n17336 0.054
R12861 GND.n17175 GND.n17162 0.054
R12862 GND.n17610 GND.n17597 0.054
R12863 GND.n17436 GND.n17423 0.054
R12864 GND.n679 GND.n666 0.054
R12865 GND.n782 GND.n769 0.054
R12866 GND.n613 GND.n600 0.054
R12867 GND.n421 GND.n408 0.054
R12868 GND.n524 GND.n511 0.054
R12869 GND.n355 GND.n342 0.054
R12870 GND.n163 GND.n150 0.054
R12871 GND.n266 GND.n253 0.054
R12872 GND.n97 GND.n84 0.054
R12873 GND.n17778 GND.n17765 0.054
R12874 GND.n17855 GND.n17842 0.054
R12875 GND.n17933 GND.n17920 0.054
R12876 GND.n14649 GND.n14648 0.053
R12877 GND.n14654 GND.n14649 0.053
R12878 GND.n14589 GND.n14583 0.053
R12879 GND.n14314 GND.n14308 0.053
R12880 GND.n14281 GND.n14279 0.053
R12881 GND.n14279 GND.n14278 0.053
R12882 GND.n9486 GND.n9484 0.053
R12883 GND.n9484 GND.n9483 0.053
R12884 GND.n1828 GND.n1827 0.053
R12885 GND.n1833 GND.n1828 0.053
R12886 GND.n3467 GND.n3465 0.053
R12887 GND.n3465 GND.n3464 0.053
R12888 GND.n2416 GND.n2409 0.053
R12889 GND.n2124 GND.n2122 0.053
R12890 GND.n2122 GND.n2121 0.053
R12891 GND.n2157 GND.n2151 0.053
R12892 GND.n7068 GND.n7067 0.053
R12893 GND.n8068 GND.n8067 0.053
R12894 GND.n13418 GND.n13417 0.053
R12895 GND.n12620 GND.n12619 0.053
R12896 GND.n12612 GND.n12611 0.053
R12897 GND.n13427 GND.n13426 0.053
R12898 GND.n12910 GND.n12906 0.053
R12899 GND.n11782 GND.n11779 0.053
R12900 GND.n12467 GND.n12463 0.053
R12901 GND.n12471 GND.n12470 0.053
R12902 GND.n13137 GND.n13134 0.053
R12903 GND.n12914 GND.n12913 0.053
R12904 GND.n7632 GND.n7629 0.053
R12905 GND.n7927 GND.n7924 0.053
R12906 GND.n8059 GND.n8058 0.053
R12907 GND.n7077 GND.n7076 0.053
R12908 GND.n6253 GND.n6252 0.053
R12909 GND.n11234 GND.n11233 0.053
R12910 GND.n13641 GND.n13640 0.053
R12911 GND.n14832 GND.n14831 0.053
R12912 GND.n16104 GND.n16103 0.053
R12913 GND.n968 GND.n967 0.053
R12914 GND.n960 GND.n959 0.053
R12915 GND.n1136 GND.n1133 0.053
R12916 GND.n9804 GND.n9803 0.053
R12917 GND.n1394 GND.n1393 0.053
R12918 GND.n1403 GND.n1402 0.053
R12919 GND.n1199 GND.n1196 0.053
R12920 GND.n8794 GND.n8793 0.053
R12921 GND.n10055 GND.n10054 0.053
R12922 GND.n9103 GND.n9102 0.053
R12923 GND.n5587 GND.n5586 0.053
R12924 GND.n4328 GND.n4327 0.053
R12925 GND.n4320 GND.n4319 0.053
R12926 GND.n15630 GND.n15629 0.053
R12927 GND.n4670 GND.n4669 0.053
R12928 GND.n5016 GND.n5015 0.053
R12929 GND.n5008 GND.n5007 0.053
R12930 GND.n4662 GND.n4661 0.053
R12931 GND.n3061 GND.n3060 0.053
R12932 GND.n3261 GND.n3260 0.053
R12933 GND.n14824 GND.n14823 0.053
R12934 GND.n10485 GND.n10484 0.053
R12935 GND.n15639 GND.n15638 0.053
R12936 GND.n15192 GND.n15191 0.053
R12937 GND.n3749 GND.n3748 0.053
R12938 GND.n3917 GND.n3914 0.053
R12939 GND.n5579 GND.n5578 0.053
R12940 GND.n5755 GND.n5752 0.053
R12941 GND.n7973 GND.n6120 0.053
R12942 GND.n7587 GND.n7586 0.053
R12943 GND.n9963 GND.n1185 0.053
R12944 GND.n2907 GND.n2906 0.053
R12945 GND.n16558 GND.n16556 0.053
R12946 GND.n16819 GND.n16817 0.053
R12947 GND.n17080 GND.n17078 0.053
R12948 GND.n17341 GND.n17339 0.053
R12949 GND.n17602 GND.n17600 0.053
R12950 GND.n774 GND.n772 0.053
R12951 GND.n516 GND.n514 0.053
R12952 GND.n258 GND.n256 0.053
R12953 GND.n17847 GND.n17845 0.053
R12954 GND.n12710 GND.n12709 0.051
R12955 GND.n13723 GND.n11004 0.051
R12956 GND.n13515 GND.n13510 0.051
R12957 GND.n13546 GND.n13545 0.051
R12958 GND.n6523 GND.n6522 0.051
R12959 GND.n8156 GND.n8151 0.051
R12960 GND.n7199 GND.n7198 0.051
R12961 GND.n7168 GND.n7163 0.051
R12962 GND.n8702 GND.n8701 0.051
R12963 GND.n1182 GND.n1181 0.051
R12964 GND.n3179 GND.n3178 0.051
R12965 GND.n5099 GND.n1932 0.051
R12966 GND.n2673 GND.n2672 0.051
R12967 GND.n4922 GND.n4921 0.051
R12968 GND.n15758 GND.n15757 0.051
R12969 GND.n15723 GND.n15718 0.051
R12970 GND.n14920 GND.n14919 0.051
R12971 GND.n14664 GND.n14661 0.05
R12972 GND.n14626 GND.n14625 0.05
R12973 GND.n14354 GND.n14353 0.05
R12974 GND.n14271 GND.n14270 0.05
R12975 GND.n9476 GND.n9475 0.05
R12976 GND.n1843 GND.n1840 0.05
R12977 GND.n3457 GND.n3456 0.05
R12978 GND.n2453 GND.n2452 0.05
R12979 GND.n2114 GND.n2113 0.05
R12980 GND.n2194 GND.n2193 0.05
R12981 GND.n557 GND.n556 0.05
R12982 GND.n299 GND.n298 0.05
R12983 GND.n41 GND.n40 0.05
R12984 GND.n17877 GND.n17876 0.05
R12985 GND.n16440 GND.n16437 0.049
R12986 GND.n16526 GND.n16523 0.049
R12987 GND.n16349 GND.n16346 0.049
R12988 GND.n16701 GND.n16698 0.049
R12989 GND.n16787 GND.n16784 0.049
R12990 GND.n16610 GND.n16607 0.049
R12991 GND.n16962 GND.n16959 0.049
R12992 GND.n17048 GND.n17045 0.049
R12993 GND.n16871 GND.n16868 0.049
R12994 GND.n17223 GND.n17220 0.049
R12995 GND.n17309 GND.n17306 0.049
R12996 GND.n17132 GND.n17129 0.049
R12997 GND.n17484 GND.n17481 0.049
R12998 GND.n17570 GND.n17567 0.049
R12999 GND.n17393 GND.n17390 0.049
R13000 GND.n699 GND.n697 0.049
R13001 GND.n726 GND.n724 0.049
R13002 GND.n441 GND.n439 0.049
R13003 GND.n468 GND.n466 0.049
R13004 GND.n183 GND.n181 0.049
R13005 GND.n210 GND.n208 0.049
R13006 GND.n17798 GND.n17796 0.049
R13007 GND.n17720 GND.n17718 0.049
R13008 GND.n6043 GND.n6040 0.049
R13009 GND.n7411 GND.n7403 0.049
R13010 GND.n9275 GND.n9272 0.049
R13011 GND.n10657 GND.n10656 0.048
R13012 GND.n14070 GND.n14067 0.048
R13013 GND.n3542 GND.n3539 0.048
R13014 GND.n4868 GND.n4867 0.048
R13015 GND.n10823 GND.n10820 0.048
R13016 GND.n13922 GND.n13919 0.048
R13017 GND.n10942 GND.n10939 0.048
R13018 GND.n10991 GND.n10988 0.048
R13019 GND.n12791 GND.n12790 0.048
R13020 GND.n11484 GND.n11481 0.048
R13021 GND.n11544 GND.n11541 0.048
R13022 GND.n11021 GND.n11018 0.048
R13023 GND.n13246 GND.n13243 0.048
R13024 GND.n11398 GND.n11397 0.048
R13025 GND.n6069 GND.n6068 0.048
R13026 GND.n8330 GND.n8329 0.048
R13027 GND.n6374 GND.n6371 0.048
R13028 GND.n5953 GND.n5950 0.048
R13029 GND.n6484 GND.n6483 0.048
R13030 GND.n6866 GND.n6863 0.048
R13031 GND.n6631 GND.n6628 0.048
R13032 GND.n6789 GND.n6788 0.048
R13033 GND.n6539 GND.n6538 0.048
R13034 GND.n6948 GND.n6947 0.048
R13035 GND.n9372 GND.n9371 0.048
R13036 GND.n1779 GND.n1778 0.048
R13037 GND.n8626 GND.n8623 0.048
R13038 GND.n2571 GND.n2570 0.048
R13039 GND.n2284 GND.n2281 0.048
R13040 GND.n5179 GND.n5178 0.048
R13041 GND.n2888 GND.n2885 0.048
R13042 GND.n15796 GND.n15793 0.048
R13043 GND.n15350 GND.n15347 0.048
R13044 GND.n14428 GND.n14427 0.048
R13045 GND.n15042 GND.n15039 0.048
R13046 GND.n16424 GND.n16423 0.048
R13047 GND.n16505 GND.n16503 0.048
R13048 GND.n16685 GND.n16684 0.048
R13049 GND.n16766 GND.n16764 0.048
R13050 GND.n16946 GND.n16945 0.048
R13051 GND.n17027 GND.n17025 0.048
R13052 GND.n17207 GND.n17206 0.048
R13053 GND.n17288 GND.n17286 0.048
R13054 GND.n17468 GND.n17467 0.048
R13055 GND.n17549 GND.n17547 0.048
R13056 GND.n16334 GND.n16333 0.048
R13057 GND.n16595 GND.n16594 0.048
R13058 GND.n16856 GND.n16855 0.048
R13059 GND.n17117 GND.n17116 0.048
R13060 GND.n17378 GND.n17377 0.048
R13061 GND.n636 GND.n633 0.048
R13062 GND.n738 GND.n735 0.048
R13063 GND.n570 GND.n567 0.048
R13064 GND.n378 GND.n375 0.048
R13065 GND.n480 GND.n477 0.048
R13066 GND.n312 GND.n309 0.048
R13067 GND.n120 GND.n117 0.048
R13068 GND.n222 GND.n219 0.048
R13069 GND.n54 GND.n51 0.048
R13070 GND.n17735 GND.n17732 0.048
R13071 GND.n17811 GND.n17808 0.048
R13072 GND.n17890 GND.n17887 0.048
R13073 GND.n5428 GND.n5244 0.047
R13074 GND.n17653 GND.n17652 0.047
R13075 GND.n11248 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE
+ 0.045
R13076 GND.n13655 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE
+ 0.045
R13077 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE GND.n12263
+ 0.045
R13078 GND.n12352 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE
+ 0.045
R13079 GND.n13076 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE
+ 0.045
R13080 GND.n12974 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.045
R13081 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE GND.n8049
+ 0.045
R13082 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE GND.n7058
+ 0.045
R13083 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE GND.n16006
+ 0.045
R13084 GND.n16091 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE
+ 0.045
R13085 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE GND.n9706
+ 0.045
R13086 GND.n9791 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.045
R13087 GND.n10243 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SUBSTRATE
+ 0.045
R13088 GND.n10069 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE
+ 0.045
R13089 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE GND.n9005
+ 0.045
R13090 GND.n9090 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE
+ 0.045
R13091 GND.n4435 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SUBSTRATE
+ 0.045
R13092 GND.n4338 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE
+ 0.045
R13093 GND.n5031 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SUBSTRATE
+ 0.045
R13094 GND.n4685 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SUBSTRATE
+ 0.045
R13095 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SUBSTRATE GND.n15620
+ 0.045
R13096 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SUBSTRATE GND.n15182
+ 0.045
R13097 GND.n16476 GND.n16475 0.045
R13098 GND.n16535 GND.n16532 0.045
R13099 GND.n16360 GND.n16357 0.045
R13100 GND.n16737 GND.n16736 0.045
R13101 GND.n16796 GND.n16793 0.045
R13102 GND.n16621 GND.n16618 0.045
R13103 GND.n16998 GND.n16997 0.045
R13104 GND.n17057 GND.n17054 0.045
R13105 GND.n16882 GND.n16879 0.045
R13106 GND.n17259 GND.n17258 0.045
R13107 GND.n17318 GND.n17315 0.045
R13108 GND.n17143 GND.n17140 0.045
R13109 GND.n17520 GND.n17519 0.045
R13110 GND.n17579 GND.n17576 0.045
R13111 GND.n17404 GND.n17401 0.045
R13112 GND.n8387 GND.n8382 0.044
R13113 GND.n7431 GND.n7378 0.044
R13114 GND.n9245 GND.n9244 0.044
R13115 GND.n14502 GND.n14499 0.043
R13116 GND.n14660 GND.n14659 0.043
R13117 GND.n14541 GND.n14538 0.043
R13118 GND.n14628 GND.n14627 0.043
R13119 GND.n14131 GND.n14128 0.043
R13120 GND.n14357 GND.n14355 0.043
R13121 GND.n14173 GND.n14170 0.043
R13122 GND.n14274 GND.n14272 0.043
R13123 GND.n1673 GND.n1672 0.043
R13124 GND.n9479 GND.n9477 0.043
R13125 GND.n1594 GND.n1591 0.043
R13126 GND.n1839 GND.n1838 0.043
R13127 GND.n2466 GND.n2465 0.043
R13128 GND.n3460 GND.n3458 0.043
R13129 GND.n2209 GND.n2206 0.043
R13130 GND.n2456 GND.n2454 0.043
R13131 GND.n2015 GND.n2012 0.043
R13132 GND.n2117 GND.n2115 0.043
R13133 GND.n1972 GND.n1969 0.043
R13134 GND.n2197 GND.n2195 0.043
R13135 GND.n648 GND.n645 0.043
R13136 GND.n750 GND.n747 0.043
R13137 GND.n582 GND.n579 0.043
R13138 GND.n390 GND.n387 0.043
R13139 GND.n492 GND.n489 0.043
R13140 GND.n324 GND.n321 0.043
R13141 GND.n132 GND.n129 0.043
R13142 GND.n234 GND.n231 0.043
R13143 GND.n66 GND.n63 0.043
R13144 GND.n17747 GND.n17744 0.043
R13145 GND.n17823 GND.n17820 0.043
R13146 GND.n17902 GND.n17899 0.043
R13147 GND.n9244 GND.n9241 0.042
R13148 GND.n12120 GND.n12115 0.041
R13149 GND.n12495 GND.n12494 0.041
R13150 GND.n8388 GND.n8387 0.041
R13151 GND.n8375 GND.n8369 0.041
R13152 GND.n6111 GND.n6108 0.041
R13153 GND.n7424 GND.n7418 0.041
R13154 GND.n7384 GND.n7382 0.041
R13155 GND.n830 GND.n823 0.041
R13156 GND.n9259 GND.n9257 0.041
R13157 GND.n9419 GND.n9417 0.041
R13158 GND.n10372 GND.n10371 0.041
R13159 GND.n16338 GND.n16335 0.04
R13160 GND.n16599 GND.n16596 0.04
R13161 GND.n16860 GND.n16857 0.04
R13162 GND.n17121 GND.n17118 0.04
R13163 GND.n17382 GND.n17379 0.04
R13164 GND.n14640 GND.n14637 0.04
R13165 GND.n14574 GND.n14571 0.04
R13166 GND.n14296 GND.n14293 0.04
R13167 GND.n14290 GND.n14289 0.04
R13168 GND.n8150 GND.n5851 0.04
R13169 GND.n6527 GND.n6524 0.04
R13170 GND.n13722 GND.n13552 0.04
R13171 GND.n12704 GND.n11724 0.04
R13172 GND.n9495 GND.n9494 0.04
R13173 GND.n1819 GND.n1816 0.04
R13174 GND.n3476 GND.n3475 0.04
R13175 GND.n2397 GND.n2394 0.04
R13176 GND.n2133 GND.n2132 0.04
R13177 GND.n2139 GND.n2136 0.04
R13178 GND.n16464 GND.n16463 0.04
R13179 GND.n16546 GND.n16543 0.04
R13180 GND.n16371 GND.n16368 0.04
R13181 GND.n16725 GND.n16724 0.04
R13182 GND.n16807 GND.n16804 0.04
R13183 GND.n16632 GND.n16629 0.04
R13184 GND.n16986 GND.n16985 0.04
R13185 GND.n17068 GND.n17065 0.04
R13186 GND.n16893 GND.n16890 0.04
R13187 GND.n17247 GND.n17246 0.04
R13188 GND.n17329 GND.n17326 0.04
R13189 GND.n17154 GND.n17151 0.04
R13190 GND.n17508 GND.n17507 0.04
R13191 GND.n17590 GND.n17587 0.04
R13192 GND.n17415 GND.n17412 0.04
R13193 GND.n17624 GND.n17623 0.04
R13194 GND.n17631 GND.n17630 0.04
R13195 GND.n17638 GND.n17637 0.04
R13196 GND.n17645 GND.n17644 0.04
R13197 GND.n659 GND.n656 0.04
R13198 GND.n762 GND.n759 0.04
R13199 GND.n594 GND.n591 0.04
R13200 GND.n401 GND.n398 0.04
R13201 GND.n504 GND.n501 0.04
R13202 GND.n336 GND.n333 0.04
R13203 GND.n143 GND.n140 0.04
R13204 GND.n246 GND.n243 0.04
R13205 GND.n78 GND.n75 0.04
R13206 GND.n17758 GND.n17755 0.04
R13207 GND.n17835 GND.n17832 0.04
R13208 GND.n17914 GND.n17911 0.04
R13209 GND.n17691 GND.n17690 0.04
R13210 GND.n17677 GND.n17676 0.04
R13211 GND.n10667 GND.n10666 0.039
R13212 GND.n14060 GND.n14057 0.039
R13213 GND.n3532 GND.n3529 0.039
R13214 GND.n4878 GND.n4877 0.039
R13215 GND.n10813 GND.n10810 0.039
R13216 GND.n13912 GND.n13909 0.039
R13217 GND.n10932 GND.n10929 0.039
R13218 GND.n10981 GND.n10978 0.039
R13219 GND.n12801 GND.n12800 0.039
R13220 GND.n11474 GND.n11471 0.039
R13221 GND.n11534 GND.n11531 0.039
R13222 GND.n11626 GND.n11625 0.039
R13223 GND.n13236 GND.n13233 0.039
R13224 GND.n11408 GND.n11407 0.039
R13225 GND.n6079 GND.n6078 0.039
R13226 GND.n8340 GND.n8339 0.039
R13227 GND.n6390 GND.n6389 0.039
R13228 GND.n5943 GND.n5940 0.039
R13229 GND.n6493 GND.n6492 0.039
R13230 GND.n6856 GND.n6853 0.039
R13231 GND.n6621 GND.n6618 0.039
R13232 GND.n6799 GND.n6798 0.039
R13233 GND.n6549 GND.n6548 0.039
R13234 GND.n6958 GND.n6957 0.039
R13235 GND.n9382 GND.n9381 0.039
R13236 GND.n1789 GND.n1788 0.039
R13237 GND.n8616 GND.n8613 0.039
R13238 GND.n2581 GND.n2580 0.039
R13239 GND.n2319 GND.n2318 0.039
R13240 GND.n5189 GND.n5188 0.039
R13241 GND.n2878 GND.n2875 0.039
R13242 GND.n15786 GND.n15783 0.039
R13243 GND.n15340 GND.n15337 0.039
R13244 GND.n14438 GND.n14437 0.039
R13245 GND.n15032 GND.n15029 0.039
R13246 GND.n4559 GND.n4558 0.039
R13247 GND.n14492 GND.n14490 0.038
R13248 GND.n14666 GND.n14664 0.038
R13249 GND.n14676 GND.n14673 0.038
R13250 GND.n15450 GND.n15448 0.038
R13251 GND.n14625 GND.n14622 0.038
R13252 GND.n14615 GND.n14613 0.038
R13253 GND.n10621 GND.n10619 0.038
R13254 GND.n10631 GND.n10628 0.038
R13255 GND.n10694 GND.n10693 0.038
R13256 GND.n15489 GND.n15486 0.038
R13257 GND.n15479 GND.n15477 0.038
R13258 GND.n14035 GND.n10715 0.038
R13259 GND.n14121 GND.n14119 0.038
R13260 GND.n14353 GND.n14350 0.038
R13261 GND.n14343 GND.n14341 0.038
R13262 GND.n14163 GND.n14161 0.038
R13263 GND.n14270 GND.n14267 0.038
R13264 GND.n14260 GND.n14258 0.038
R13265 GND.n3575 GND.n3572 0.038
R13266 GND.n3565 GND.n3563 0.038
R13267 GND.n3506 GND.n1935 0.038
R13268 GND.n4833 GND.n4831 0.038
R13269 GND.n4843 GND.n4840 0.038
R13270 GND.n4904 GND.n4903 0.038
R13271 GND.n10785 GND.n10783 0.038
R13272 GND.n10763 GND.n10760 0.038
R13273 GND.n10753 GND.n10751 0.038
R13274 GND.n13885 GND.n13883 0.038
R13275 GND.n13943 GND.n13941 0.038
R13276 GND.n13953 GND.n13950 0.038
R13277 GND.n13825 GND.n13822 0.038
R13278 GND.n13815 GND.n13813 0.038
R13279 GND.n10907 GND.n10905 0.038
R13280 GND.n13769 GND.n13767 0.038
R13281 GND.n13779 GND.n13776 0.038
R13282 GND.n10956 GND.n10718 0.038
R13283 GND.n12756 GND.n12754 0.038
R13284 GND.n12766 GND.n12763 0.038
R13285 GND.n12828 GND.n12827 0.038
R13286 GND.n11446 GND.n11444 0.038
R13287 GND.n11669 GND.n11667 0.038
R13288 GND.n11679 GND.n11676 0.038
R13289 GND.n11507 GND.n11505 0.038
R13290 GND.n11565 GND.n11563 0.038
R13291 GND.n11575 GND.n11572 0.038
R13292 GND.n11067 GND.n11064 0.038
R13293 GND.n11057 GND.n11055 0.038
R13294 GND.n11653 GND.n11652 0.038
R13295 GND.n13280 GND.n13277 0.038
R13296 GND.n13270 GND.n13268 0.038
R13297 GND.n13211 GND.n11721 0.038
R13298 GND.n11365 GND.n11363 0.038
R13299 GND.n11375 GND.n11372 0.038
R13300 GND.n11434 GND.n11433 0.038
R13301 GND.n8205 GND.n8203 0.038
R13302 GND.n8215 GND.n8212 0.038
R13303 GND.n6106 GND.n6105 0.038
R13304 GND.n8294 GND.n8292 0.038
R13305 GND.n8304 GND.n8301 0.038
R13306 GND.n8367 GND.n8366 0.038
R13307 GND.n5848 GND.n5847 0.038
R13308 GND.n6353 GND.n6350 0.038
R13309 GND.n5860 GND.n5857 0.038
R13310 GND.n5915 GND.n5913 0.038
R13311 GND.n5979 GND.n5977 0.038
R13312 GND.n5989 GND.n5986 0.038
R13313 GND.n6517 GND.n6516 0.038
R13314 GND.n6466 GND.n6463 0.038
R13315 GND.n6456 GND.n6454 0.038
R13316 GND.n6891 GND.n6889 0.038
R13317 GND.n6901 GND.n6898 0.038
R13318 GND.n6593 GND.n6591 0.038
R13319 GND.n6656 GND.n6654 0.038
R13320 GND.n6666 GND.n6663 0.038
R13321 GND.n6753 GND.n6751 0.038
R13322 GND.n6763 GND.n6760 0.038
R13323 GND.n6826 GND.n6825 0.038
R13324 GND.n7477 GND.n7475 0.038
R13325 GND.n7487 GND.n7484 0.038
R13326 GND.n6576 GND.n6575 0.038
R13327 GND.n7541 GND.n7538 0.038
R13328 GND.n7531 GND.n7529 0.038
R13329 GND.n6985 GND.n6984 0.038
R13330 GND.n9338 GND.n9336 0.038
R13331 GND.n9348 GND.n9345 0.038
R13332 GND.n9408 GND.n9407 0.038
R13333 GND.n1743 GND.n1741 0.038
R13334 GND.n1753 GND.n1750 0.038
R13335 GND.n1815 GND.n1814 0.038
R13336 GND.n1681 GND.n1680 0.038
R13337 GND.n9475 GND.n9472 0.038
R13338 GND.n9465 GND.n9463 0.038
R13339 GND.n1584 GND.n1582 0.038
R13340 GND.n1845 GND.n1843 0.038
R13341 GND.n1855 GND.n1852 0.038
R13342 GND.n8655 GND.n8652 0.038
R13343 GND.n8645 GND.n8643 0.038
R13344 GND.n8590 GND.n1897 0.038
R13345 GND.n2536 GND.n2534 0.038
R13346 GND.n2546 GND.n2543 0.038
R13347 GND.n2608 GND.n2607 0.038
R13348 GND.n2474 GND.n2473 0.038
R13349 GND.n3456 GND.n3453 0.038
R13350 GND.n3446 GND.n3444 0.038
R13351 GND.n3164 GND.n3163 0.038
R13352 GND.n2452 GND.n2449 0.038
R13353 GND.n2442 GND.n2440 0.038
R13354 GND.n2374 GND.n2372 0.038
R13355 GND.n2384 GND.n2381 0.038
R13356 GND.n2301 GND.n2299 0.038
R13357 GND.n5145 GND.n5143 0.038
R13358 GND.n5155 GND.n5152 0.038
R13359 GND.n5216 GND.n5215 0.038
R13360 GND.n2005 GND.n2003 0.038
R13361 GND.n2113 GND.n2110 0.038
R13362 GND.n2103 GND.n2101 0.038
R13363 GND.n1962 GND.n1960 0.038
R13364 GND.n2193 GND.n2190 0.038
R13365 GND.n2183 GND.n2181 0.038
R13366 GND.n2922 GND.n2919 0.038
R13367 GND.n2912 GND.n2910 0.038
R13368 GND.n2852 GND.n2850 0.038
R13369 GND.n15830 GND.n15827 0.038
R13370 GND.n15820 GND.n15818 0.038
R13371 GND.n15761 GND.n15759 0.038
R13372 GND.n15385 GND.n15382 0.038
R13373 GND.n15375 GND.n15373 0.038
R13374 GND.n15315 GND.n15313 0.038
R13375 GND.n14966 GND.n14964 0.038
R13376 GND.n14976 GND.n14973 0.038
R13377 GND.n14464 GND.n14463 0.038
R13378 GND.n15071 GND.n15068 0.038
R13379 GND.n15061 GND.n15059 0.038
R13380 GND.n15007 GND.n14403 0.038
R13381 GND.n561 GND.n558 0.037
R13382 GND.n303 GND.n300 0.037
R13383 GND.n45 GND.n42 0.037
R13384 GND.n17881 GND.n17878 0.037
R13385 GND.n13791 GND 0.037
R13386 GND.n11008 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SOURCE 0.037
R13387 GND.n6360 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SOURCE 0.037
R13388 GND.n7511 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SOURCE 0.037
R13389 GND.n9511 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE 0.037
R13390 GND.n1925 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SOURCE
+ 0.037
R13391 GND.n3490 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SOURCE
+ 0.037
R13392 GND.n15461 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SOURCE
+ 0.037
R13393 GND.n14999 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SOURCE
+ 0.037
R13394 GND.n8885 GND.n8879 0.037
R13395 GND.n16321 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE
+ 0.037
R13396 GND.n16582 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE
+ 0.037
R13397 GND.n16843 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SOURCE
+ 0.037
R13398 GND.n17104 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SOURCE
+ 0.037
R13399 GND.n17365 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SOURCE
+ 0.037
R13400 GND.n542 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SOURCE 0.037
R13401 GND.n284 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE 0.037
R13402 GND.n26 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SOURCE 0.037
R13403 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SOURCE GND.n17936
+ 0.037
R13404 GND.n5962 GND.n5961 0.036
R13405 GND.n6383 GND.n6382 0.036
R13406 GND.n6475 GND.n6473 0.036
R13407 GND.n6875 GND.n6874 0.036
R13408 GND.n6640 GND.n6639 0.036
R13409 GND.n16452 GND.n16451 0.036
R13410 GND.n16713 GND.n16712 0.036
R13411 GND.n16974 GND.n16973 0.036
R13412 GND.n17235 GND.n17234 0.036
R13413 GND.n17496 GND.n17495 0.036
R13414 GND.n10765 GND.n10764 0.036
R13415 GND.n12769 GND.n12767 0.036
R13416 GND.n11664 GND.n11663 0.036
R13417 GND.n13265 GND.n13264 0.036
R13418 GND.n8307 GND.n8305 0.036
R13419 GND.n6359 GND.n6358 0.036
R13420 GND.n5974 GND.n5973 0.036
R13421 GND.n6468 GND.n6467 0.036
R13422 GND.n6886 GND.n6885 0.036
R13423 GND.n6651 GND.n6650 0.036
R13424 GND.n7490 GND.n7488 0.036
R13425 GND.n2385 GND.n2334 0.036
R13426 GND.n15815 GND.n15814 0.036
R13427 GND.n16384 GND.n16382 0.036
R13428 GND.n16645 GND.n16643 0.036
R13429 GND.n16906 GND.n16904 0.036
R13430 GND.n17167 GND.n17165 0.036
R13431 GND.n17428 GND.n17426 0.036
R13432 GND.n605 GND.n603 0.036
R13433 GND.n671 GND.n669 0.036
R13434 GND.n347 GND.n345 0.036
R13435 GND.n413 GND.n411 0.036
R13436 GND.n89 GND.n87 0.036
R13437 GND.n155 GND.n153 0.036
R13438 GND.n17925 GND.n17923 0.036
R13439 GND.n17770 GND.n17768 0.036
R13440 GND.n2296 GND.n2290 0.036
R13441 GND.n14523 GND.n14522 0.036
R13442 GND.n14549 GND.n14548 0.036
R13443 GND.n14138 GND.n14137 0.036
R13444 GND.n14191 GND.n14190 0.036
R13445 GND.n10904 GND.n10890 0.036
R13446 GND.n11126 GND.n11123 0.036
R13447 GND.n1664 GND.n1663 0.036
R13448 GND.n1613 GND.n1612 0.036
R13449 GND.n2246 GND.n2245 0.036
R13450 GND.n2217 GND.n2216 0.036
R13451 GND.n2033 GND.n2032 0.036
R13452 GND.n1980 GND.n1979 0.036
R13453 GND.n14100 GND.n14097 0.036
R13454 GND.n15312 GND.n14379 0.036
R13455 GND.n10634 GND.n10632 0.036
R13456 GND.n15474 GND.n15473 0.036
R13457 GND.n3560 GND.n3559 0.036
R13458 GND.n4846 GND.n4844 0.036
R13459 GND.n13938 GND.n13937 0.036
R13460 GND.n13810 GND.n13809 0.036
R13461 GND.n13781 GND.n13780 0.036
R13462 GND.n11560 GND.n11559 0.036
R13463 GND.n11052 GND.n11051 0.036
R13464 GND.n11377 GND.n11376 0.036
R13465 GND.n8218 GND.n8216 0.036
R13466 GND.n6766 GND.n6764 0.036
R13467 GND.n7526 GND.n7525 0.036
R13468 GND.n9351 GND.n9349 0.036
R13469 GND.n1756 GND.n1754 0.036
R13470 GND.n8640 GND.n8639 0.036
R13471 GND.n2549 GND.n2547 0.036
R13472 GND.n5158 GND.n5156 0.036
R13473 GND.n15370 GND.n15369 0.036
R13474 GND.n14978 GND.n14977 0.036
R13475 GND.n15056 GND.n15055 0.036
R13476 GND.n15456 GND.n14360 0.035
R13477 GND.n9519 GND.n9504 0.035
R13478 GND.n2460 GND.n2459 0.035
R13479 GND.n3496 GND.n2200 0.035
R13480 GND.n14994 GND.n14409 0.035
R13481 GND.n14000 GND.n13999 0.035
R13482 GND.n11145 GND.n11144 0.035
R13483 GND.n15294 GND.n15291 0.035
R13484 GND.n14838 GND.n14836 0.034
R13485 GND.n14817 GND.n14815 0.034
R13486 GND.n6259 GND.n6257 0.034
R13487 GND.n6239 GND.n6237 0.034
R13488 GND.n12626 GND.n12624 0.034
R13489 GND.n12605 GND.n12603 0.034
R13490 GND.n10838 GND.n10837 0.034
R13491 GND.n12536 GND.n12535 0.034
R13492 GND.n13796 GND.n13795 0.034
R13493 GND.n11240 GND.n11238 0.034
R13494 GND.n11220 GND.n11218 0.034
R13495 GND.n13647 GND.n13645 0.034
R13496 GND.n13627 GND.n13625 0.034
R13497 GND.n11499 GND.n11498 0.034
R13498 GND.n11034 GND.n11033 0.034
R13499 GND.n11038 GND.n11037 0.034
R13500 GND.n13412 GND.n13410 0.034
R13501 GND.n13433 GND.n13431 0.034
R13502 GND.n11957 GND.n11956 0.034
R13503 GND.n11953 GND.n11952 0.034
R13504 GND.n11885 GND.n11883 0.034
R13505 GND.n11880 GND.n11879 0.034
R13506 GND.n12265 GND.n12264 0.034
R13507 GND.n12270 GND.n12268 0.034
R13508 GND.n12338 GND.n12337 0.034
R13509 GND.n12342 GND.n12341 0.034
R13510 GND.n13063 GND.n13062 0.034
R13511 GND.n13059 GND.n13058 0.034
R13512 GND.n12990 GND.n12988 0.034
R13513 GND.n12985 GND.n12984 0.034
R13514 GND.n7753 GND.n7752 0.034
R13515 GND.n7758 GND.n7756 0.034
R13516 GND.n7827 GND.n7826 0.034
R13517 GND.n7831 GND.n7830 0.034
R13518 GND.n8233 GND.n8232 0.034
R13519 GND.n6410 GND.n6409 0.034
R13520 GND.n6405 GND.n6404 0.034
R13521 GND.n8074 GND.n8072 0.034
R13522 GND.n8053 GND.n8051 0.034
R13523 GND.n7062 GND.n7060 0.034
R13524 GND.n7083 GND.n7081 0.034
R13525 GND.n6588 GND.n6587 0.034
R13526 GND.n7504 GND.n7503 0.034
R13527 GND.n7509 GND.n7508 0.034
R13528 GND.n7301 GND.n7299 0.034
R13529 GND.n7279 GND.n7277 0.034
R13530 GND.n16008 GND.n16007 0.034
R13531 GND.n16017 GND.n16015 0.034
R13532 GND.n16098 GND.n16096 0.034
R13533 GND.n16118 GND.n16116 0.034
R13534 GND.n1062 GND.n1061 0.034
R13535 GND.n1055 GND.n1053 0.034
R13536 GND.n973 GND.n972 0.034
R13537 GND.n953 GND.n951 0.034
R13538 GND.n9708 GND.n9707 0.034
R13539 GND.n9717 GND.n9715 0.034
R13540 GND.n9798 GND.n9796 0.034
R13541 GND.n9818 GND.n9816 0.034
R13542 GND.n1298 GND.n1297 0.034
R13543 GND.n1307 GND.n1305 0.034
R13544 GND.n1388 GND.n1386 0.034
R13545 GND.n1409 GND.n1407 0.034
R13546 GND.n10235 GND.n10233 0.034
R13547 GND.n10213 GND.n10211 0.034
R13548 GND.n8800 GND.n8798 0.034
R13549 GND.n8780 GND.n8778 0.034
R13550 GND.n8505 GND.n8503 0.034
R13551 GND.n8483 GND.n8481 0.034
R13552 GND.n9510 GND.n9509 0.034
R13553 GND.n9516 GND.n9515 0.034
R13554 GND.n10061 GND.n10059 0.034
R13555 GND.n10041 GND.n10039 0.034
R13556 GND.n9007 GND.n9006 0.034
R13557 GND.n9016 GND.n9014 0.034
R13558 GND.n9097 GND.n9095 0.034
R13559 GND.n9117 GND.n9115 0.034
R13560 GND.n4422 GND.n4421 0.034
R13561 GND.n4415 GND.n4413 0.034
R13562 GND.n4333 GND.n4332 0.034
R13563 GND.n4313 GND.n4311 0.034
R13564 GND.n3255 GND.n3253 0.034
R13565 GND.n3275 GND.n3273 0.034
R13566 GND.n5022 GND.n5020 0.034
R13567 GND.n5001 GND.n4999 0.034
R13568 GND.n2389 GND.n2388 0.034
R13569 GND.n2393 GND.n2392 0.034
R13570 GND.n2844 GND.n2843 0.034
R13571 GND.n3495 GND.n3494 0.034
R13572 GND.n4676 GND.n4674 0.034
R13573 GND.n4655 GND.n4653 0.034
R13574 GND.n3055 GND.n3053 0.034
R13575 GND.n3075 GND.n3073 0.034
R13576 GND.n10479 GND.n10477 0.034
R13577 GND.n10499 GND.n10497 0.034
R13578 GND.n15624 GND.n15622 0.034
R13579 GND.n15645 GND.n15643 0.034
R13580 GND.n14366 GND.n14365 0.034
R13581 GND.n15459 GND.n15458 0.034
R13582 GND.n14992 GND.n14991 0.034
R13583 GND.n14997 GND.n14996 0.034
R13584 GND.n15186 GND.n15184 0.034
R13585 GND.n15206 GND.n15204 0.034
R13586 GND.n3843 GND.n3842 0.034
R13587 GND.n3836 GND.n3834 0.034
R13588 GND.n3754 GND.n3753 0.034
R13589 GND.n3735 GND.n3733 0.034
R13590 GND.n4574 GND.n4569 0.034
R13591 GND.n5797 GND.n5792 0.034
R13592 GND.n5681 GND.n5680 0.034
R13593 GND.n5674 GND.n5672 0.034
R13594 GND.n5592 GND.n5591 0.034
R13595 GND.n5572 GND.n5570 0.034
R13596 GND.n5449 GND.n5448 0.034
R13597 GND.n5235 GND.n5234 0.034
R13598 GND.n14683 GND.n14680 0.033
R13599 GND.n14608 GND.n14606 0.033
R13600 GND.n10614 GND.n10612 0.033
R13601 GND.n15496 GND.n15493 0.033
R13602 GND.n14336 GND.n14334 0.033
R13603 GND.n14253 GND.n14251 0.033
R13604 GND.n3582 GND.n3579 0.033
R13605 GND.n4826 GND.n4824 0.033
R13606 GND.n10746 GND.n10744 0.033
R13607 GND.n13960 GND.n13957 0.033
R13608 GND.n13832 GND.n13829 0.033
R13609 GND.n13762 GND.n13760 0.033
R13610 GND.n12749 GND.n12747 0.033
R13611 GND.n11686 GND.n11683 0.033
R13612 GND.n11582 GND.n11579 0.033
R13613 GND.n11074 GND.n11071 0.033
R13614 GND.n13287 GND.n13284 0.033
R13615 GND.n11358 GND.n11356 0.033
R13616 GND.n8198 GND.n8196 0.033
R13617 GND.n8287 GND.n8285 0.033
R13618 GND.n5867 GND.n5864 0.033
R13619 GND.n5996 GND.n5993 0.033
R13620 GND.n6449 GND.n6447 0.033
R13621 GND.n6120 GND.n6117 0.033
R13622 GND.n6908 GND.n6905 0.033
R13623 GND.n6673 GND.n6670 0.033
R13624 GND.n6746 GND.n6744 0.033
R13625 GND.n7470 GND.n7468 0.033
R13626 GND.n7586 GND.n7583 0.033
R13627 GND.n7548 GND.n7545 0.033
R13628 GND.n9331 GND.n9329 0.033
R13629 GND.n1736 GND.n1734 0.033
R13630 GND.n9458 GND.n9456 0.033
R13631 GND.n1862 GND.n1859 0.033
R13632 GND.n8662 GND.n8659 0.033
R13633 GND.n9409 GND.n1185 0.033
R13634 GND.n2529 GND.n2527 0.033
R13635 GND.n3439 GND.n3437 0.033
R13636 GND.n2435 GND.n2433 0.033
R13637 GND.n2367 GND.n2365 0.033
R13638 GND.n5138 GND.n5136 0.033
R13639 GND.n2096 GND.n2094 0.033
R13640 GND.n2176 GND.n2174 0.033
R13641 GND.n2929 GND.n2926 0.033
R13642 GND.n15837 GND.n15834 0.033
R13643 GND.n15392 GND.n15389 0.033
R13644 GND.n14959 GND.n14957 0.033
R13645 GND.n15078 GND.n15075 0.033
R13646 GND.n3382 GND.n3379 0.032
R13647 GND.n4787 GND.n3500 0.032
R13648 GND.n16429 GND.n16426 0.032
R13649 GND.n16501 GND.n16500 0.032
R13650 GND.n16690 GND.n16687 0.032
R13651 GND.n16762 GND.n16761 0.032
R13652 GND.n16951 GND.n16948 0.032
R13653 GND.n17023 GND.n17022 0.032
R13654 GND.n17212 GND.n17209 0.032
R13655 GND.n17284 GND.n17283 0.032
R13656 GND.n17473 GND.n17470 0.032
R13657 GND.n17545 GND.n17544 0.032
R13658 GND.n14497 GND.n14495 0.031
R13659 GND.n14508 GND.n14507 0.031
R13660 GND.n14644 GND.n14642 0.031
R13661 GND.n14715 GND.n14713 0.031
R13662 GND.n14567 GND.n14565 0.031
R13663 GND.n14400 GND.n14398 0.031
R13664 GND.n10581 GND.n10579 0.031
R13665 GND.n10653 GND.n10651 0.031
R13666 GND.n10663 GND.n10661 0.031
R13667 GND.n15528 GND.n15526 0.031
R13668 GND.n14074 GND.n14072 0.031
R13669 GND.n14064 GND.n14062 0.031
R13670 GND.n14156 GND.n14154 0.031
R13671 GND.n10712 GND.n10710 0.031
R13672 GND.n14209 GND.n14207 0.031
R13673 GND.n14286 GND.n14285 0.031
R13674 GND.n14220 GND.n14218 0.031
R13675 GND.n3614 GND.n3612 0.031
R13676 GND.n3546 GND.n3544 0.031
R13677 GND.n3536 GND.n3534 0.031
R13678 GND.n4793 GND.n4791 0.031
R13679 GND.n4864 GND.n4862 0.031
R13680 GND.n4874 GND.n4872 0.031
R13681 GND.n10817 GND.n10815 0.031
R13682 GND.n10827 GND.n10825 0.031
R13683 GND.n10873 GND.n10871 0.031
R13684 GND.n13916 GND.n13914 0.031
R13685 GND.n13926 GND.n13924 0.031
R13686 GND.n13992 GND.n13990 0.031
R13687 GND.n13864 GND.n13862 0.031
R13688 GND.n10946 GND.n10944 0.031
R13689 GND.n10936 GND.n10934 0.031
R13690 GND.n13729 GND.n13727 0.031
R13691 GND.n10995 GND.n10993 0.031
R13692 GND.n10985 GND.n10983 0.031
R13693 GND.n12716 GND.n12714 0.031
R13694 GND.n12787 GND.n12785 0.031
R13695 GND.n12797 GND.n12795 0.031
R13696 GND.n11478 GND.n11476 0.031
R13697 GND.n11488 GND.n11486 0.031
R13698 GND.n11718 GND.n11716 0.031
R13699 GND.n11538 GND.n11536 0.031
R13700 GND.n11548 GND.n11546 0.031
R13701 GND.n11614 GND.n11612 0.031
R13702 GND.n11106 GND.n11104 0.031
R13703 GND.n11025 GND.n11023 0.031
R13704 GND.n11622 GND.n11620 0.031
R13705 GND.n13319 GND.n13317 0.031
R13706 GND.n13250 GND.n13248 0.031
R13707 GND.n13240 GND.n13238 0.031
R13708 GND.n11325 GND.n11323 0.031
R13709 GND.n11394 GND.n11392 0.031
R13710 GND.n11404 GND.n11402 0.031
R13711 GND.n8165 GND.n8163 0.031
R13712 GND.n6065 GND.n6063 0.031
R13713 GND.n6075 GND.n6073 0.031
R13714 GND.n8254 GND.n8252 0.031
R13715 GND.n8326 GND.n8324 0.031
R13716 GND.n8336 GND.n8334 0.031
R13717 GND.n6378 GND.n6376 0.031
R13718 GND.n5899 GND.n5897 0.031
R13719 GND.n5947 GND.n5945 0.031
R13720 GND.n5957 GND.n5955 0.031
R13721 GND.n6028 GND.n6026 0.031
R13722 GND.n6489 GND.n6488 0.031
R13723 GND.n6480 GND.n6479 0.031
R13724 GND.n6416 GND.n6414 0.031
R13725 GND.n6860 GND.n6858 0.031
R13726 GND.n6870 GND.n6868 0.031
R13727 GND.n6940 GND.n6938 0.031
R13728 GND.n6625 GND.n6623 0.031
R13729 GND.n6635 GND.n6633 0.031
R13730 GND.n6705 GND.n6703 0.031
R13731 GND.n6713 GND.n6711 0.031
R13732 GND.n6785 GND.n6783 0.031
R13733 GND.n6795 GND.n6793 0.031
R13734 GND.n7437 GND.n7435 0.031
R13735 GND.n6535 GND.n6533 0.031
R13736 GND.n6545 GND.n6543 0.031
R13737 GND.n7580 GND.n7578 0.031
R13738 GND.n6954 GND.n6952 0.031
R13739 GND.n9298 GND.n9296 0.031
R13740 GND.n9368 GND.n9366 0.031
R13741 GND.n9378 GND.n9376 0.031
R13742 GND.n1703 GND.n1701 0.031
R13743 GND.n1775 GND.n1773 0.031
R13744 GND.n1785 GND.n1783 0.031
R13745 GND.n1649 GND.n1648 0.031
R13746 GND.n9491 GND.n9490 0.031
R13747 GND.n9425 GND.n9423 0.031
R13748 GND.n1631 GND.n1629 0.031
R13749 GND.n1823 GND.n1821 0.031
R13750 GND.n1894 GND.n1892 0.031
R13751 GND.n8694 GND.n8692 0.031
R13752 GND.n8630 GND.n8628 0.031
R13753 GND.n8620 GND.n8618 0.031
R13754 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE GND.n9278 0.031
R13755 GND.n2496 GND.n2494 0.031
R13756 GND.n2567 GND.n2565 0.031
R13757 GND.n2577 GND.n2575 0.031
R13758 GND.n2264 GND.n2262 0.031
R13759 GND.n3472 GND.n3471 0.031
R13760 GND.n3406 GND.n3404 0.031
R13761 GND.n2235 GND.n2233 0.031
R13762 GND.n2629 GND.n2627 0.031
R13763 GND.n3153 GND.n3151 0.031
R13764 GND.n2287 GND.n2285 0.031
R13765 GND.n5105 GND.n5103 0.031
R13766 GND.n5175 GND.n5173 0.031
R13767 GND.n5185 GND.n5183 0.031
R13768 GND.n2051 GND.n2049 0.031
R13769 GND.n2129 GND.n2128 0.031
R13770 GND.n2063 GND.n2061 0.031
R13771 GND.n1998 GND.n1996 0.031
R13772 GND.n2656 GND.n2654 0.031
R13773 GND.n2961 GND.n2959 0.031
R13774 GND.n2892 GND.n2890 0.031
R13775 GND.n2882 GND.n2880 0.031
R13776 GND.n15869 GND.n15867 0.031
R13777 GND.n15800 GND.n15798 0.031
R13778 GND.n15790 GND.n15788 0.031
R13779 GND.n15424 GND.n15422 0.031
R13780 GND.n15354 GND.n15352 0.031
R13781 GND.n15344 GND.n15342 0.031
R13782 GND.n14926 GND.n14924 0.031
R13783 GND.n14424 GND.n14422 0.031
R13784 GND.n14434 GND.n14432 0.031
R13785 GND.n15110 GND.n15108 0.031
R13786 GND.n15046 GND.n15044 0.031
R13787 GND.n15036 GND.n15034 0.031
R13788 GND.n16460 GND.n16458 0.031
R13789 GND.n16550 GND.n16548 0.031
R13790 GND.n16375 GND.n16373 0.031
R13791 GND.n16721 GND.n16719 0.031
R13792 GND.n16811 GND.n16809 0.031
R13793 GND.n16636 GND.n16634 0.031
R13794 GND.n16982 GND.n16980 0.031
R13795 GND.n17072 GND.n17070 0.031
R13796 GND.n16897 GND.n16895 0.031
R13797 GND.n17243 GND.n17241 0.031
R13798 GND.n17333 GND.n17331 0.031
R13799 GND.n17158 GND.n17156 0.031
R13800 GND.n17504 GND.n17502 0.031
R13801 GND.n17594 GND.n17592 0.031
R13802 GND.n17419 GND.n17417 0.031
R13803 GND.n663 GND.n661 0.031
R13804 GND.n766 GND.n764 0.031
R13805 GND.n597 GND.n595 0.031
R13806 GND.n405 GND.n403 0.031
R13807 GND.n508 GND.n506 0.031
R13808 GND.n339 GND.n337 0.031
R13809 GND.n147 GND.n145 0.031
R13810 GND.n250 GND.n248 0.031
R13811 GND.n81 GND.n79 0.031
R13812 GND.n17762 GND.n17760 0.031
R13813 GND.n17839 GND.n17837 0.031
R13814 GND.n17917 GND.n17915 0.031
R13815 GND.n14851 GND.n14849 0.03
R13816 GND.n14804 GND.n14802 0.03
R13817 GND.n3999 GND.n3998 0.03
R13818 GND.n4000 GND.n3999 0.03
R13819 GND.n4109 GND.n4108 0.03
R13820 GND.n4110 GND.n4109 0.03
R13821 GND.n4112 GND.n4111 0.03
R13822 GND.n4111 GND.n4110 0.03
R13823 GND.n4002 GND.n4001 0.03
R13824 GND.n4001 GND.n4000 0.03
R13825 GND.n6271 GND.n6269 0.03
R13826 GND.n6227 GND.n6225 0.03
R13827 GND.n12639 GND.n12637 0.03
R13828 GND.n12592 GND.n12590 0.03
R13829 GND.n11252 GND.n11250 0.03
R13830 GND.n11208 GND.n11206 0.03
R13831 GND.n13659 GND.n13657 0.03
R13832 GND.n13615 GND.n13613 0.03
R13833 GND.n13399 GND.n13397 0.03
R13834 GND.n13446 GND.n13444 0.03
R13835 GND.n11974 GND.n11972 0.03
R13836 GND.n11949 GND.n11948 0.03
R13837 GND.n11889 GND.n11887 0.03
R13838 GND.n11869 GND.n11867 0.03
R13839 GND.n12250 GND.n12248 0.03
R13840 GND.n12274 GND.n12272 0.03
R13841 GND.n12334 GND.n12333 0.03
R13842 GND.n12356 GND.n12354 0.03
R13843 GND.n7619 GND.n7618 0.03
R13844 GND.n13080 GND.n13078 0.03
R13845 GND.n13055 GND.n13053 0.03
R13846 GND.n12994 GND.n12992 0.03
R13847 GND.n12973 GND.n12971 0.03
R13848 GND.n7964 GND.n6143 0.03
R13849 GND.n7738 GND.n7736 0.03
R13850 GND.n7763 GND.n7761 0.03
R13851 GND.n7823 GND.n7822 0.03
R13852 GND.n7844 GND.n7842 0.03
R13853 GND.n8087 GND.n8085 0.03
R13854 GND.n8040 GND.n8038 0.03
R13855 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE GND.n6047 0.03
R13856 GND.n7049 GND.n7047 0.03
R13857 GND.n7096 GND.n7094 0.03
R13858 GND.n7400 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE 0.03
R13859 GND.n7313 GND.n7311 0.03
R13860 GND.n7267 GND.n7265 0.03
R13861 GND.n15993 GND.n15991 0.03
R13862 GND.n16025 GND.n16023 0.03
R13863 GND.n16090 GND.n16089 0.03
R13864 GND.n16130 GND.n16128 0.03
R13865 GND.n1079 GND.n1077 0.03
R13866 GND.n1047 GND.n1045 0.03
R13867 GND.n980 GND.n979 0.03
R13868 GND.n940 GND.n938 0.03
R13869 GND.n9693 GND.n9691 0.03
R13870 GND.n9725 GND.n9723 0.03
R13871 GND.n9790 GND.n9789 0.03
R13872 GND.n9830 GND.n9828 0.03
R13873 GND.n1283 GND.n1281 0.03
R13874 GND.n1315 GND.n1313 0.03
R13875 GND.n1380 GND.n1379 0.03
R13876 GND.n1422 GND.n1420 0.03
R13877 GND.n9954 GND.n9953 0.03
R13878 GND.n10247 GND.n10245 0.03
R13879 GND.n10201 GND.n10199 0.03
R13880 GND.n8812 GND.n8810 0.03
R13881 GND.n8768 GND.n8766 0.03
R13882 GND.n8517 GND.n8515 0.03
R13883 GND.n8471 GND.n8469 0.03
R13884 GND.n10073 GND.n10071 0.03
R13885 GND.n10029 GND.n10027 0.03
R13886 GND.n8992 GND.n8990 0.03
R13887 GND.n9024 GND.n9022 0.03
R13888 GND.n9089 GND.n9088 0.03
R13889 GND.n9129 GND.n9127 0.03
R13890 GND.n4439 GND.n4437 0.03
R13891 GND.n4407 GND.n4405 0.03
R13892 GND.n4340 GND.n4339 0.03
R13893 GND.n4300 GND.n4298 0.03
R13894 GND.n3243 GND.n3241 0.03
R13895 GND.n3287 GND.n3285 0.03
R13896 GND.n5035 GND.n5033 0.03
R13897 GND.n4988 GND.n4986 0.03
R13898 GND.n4689 GND.n4687 0.03
R13899 GND.n4642 GND.n4640 0.03
R13900 GND.n3043 GND.n3041 0.03
R13901 GND.n3087 GND.n3085 0.03
R13902 GND.n10467 GND.n10465 0.03
R13903 GND.n10511 GND.n10509 0.03
R13904 GND.n15611 GND.n15609 0.03
R13905 GND.n15658 GND.n15656 0.03
R13906 GND.n15174 GND.n15172 0.03
R13907 GND.n15218 GND.n15216 0.03
R13908 GND.n3860 GND.n3858 0.03
R13909 GND.n3828 GND.n3826 0.03
R13910 GND.n3761 GND.n3760 0.03
R13911 GND.n3723 GND.n3721 0.03
R13912 GND.n10339 GND.n10334 0.03
R13913 GND.n5698 GND.n5696 0.03
R13914 GND.n5666 GND.n5664 0.03
R13915 GND.n5599 GND.n5598 0.03
R13916 GND.n5559 GND.n5557 0.03
R13917 GND.n15453 GND.n14371 0.03
R13918 GND.n14126 GND.n14124 0.03
R13919 GND.n14168 GND.n14166 0.03
R13920 GND.n1677 GND.n1676 0.03
R13921 GND.n1589 GND.n1587 0.03
R13922 GND.n2470 GND.n2469 0.03
R13923 GND.n2204 GND.n2203 0.03
R13924 GND.n2010 GND.n2008 0.03
R13925 GND.n1967 GND.n1965 0.03
R13926 GND.n3398 GND.n1924 0.03
R13927 GND.n4769 GND.n4766 0.03
R13928 GND.n695 GND.n694 0.029
R13929 GND.n722 GND.n721 0.029
R13930 GND.n437 GND.n436 0.029
R13931 GND.n464 GND.n463 0.029
R13932 GND.n179 GND.n178 0.029
R13933 GND.n206 GND.n205 0.029
R13934 GND.n17794 GND.n17793 0.029
R13935 GND.n17716 GND.n17715 0.029
R13936 GND.n17654 GND.n17653 0.029
R13937 GND.n14690 GND.n14687 0.028
R13938 GND.n14601 GND.n14599 0.028
R13939 GND.n10607 GND.n10605 0.028
R13940 GND.n15503 GND.n15500 0.028
R13941 GND.n14329 GND.n14327 0.028
R13942 GND.n14246 GND.n14244 0.028
R13943 GND.n14911 GND.n14909 0.028
R13944 GND.n14750 GND.n14741 0.028
R13945 GND.n3589 GND.n3586 0.028
R13946 GND.n4819 GND.n4817 0.028
R13947 GND.n6329 GND.n6327 0.028
R13948 GND.n6174 GND.n6165 0.028
R13949 GND.n12699 GND.n12697 0.028
R13950 GND.n10739 GND.n10737 0.028
R13951 GND.n13967 GND.n13964 0.028
R13952 GND.n13839 GND.n13836 0.028
R13953 GND.n13755 GND.n13753 0.028
R13954 GND.n11310 GND.n11308 0.028
R13955 GND.n11156 GND.n11147 0.028
R13956 GND.n13717 GND.n13715 0.028
R13957 GND.n13563 GND.n13554 0.028
R13958 GND.n12742 GND.n12740 0.028
R13959 GND.n11693 GND.n11690 0.028
R13960 GND.n11589 GND.n11586 0.028
R13961 GND.n11081 GND.n11078 0.028
R13962 GND.n13294 GND.n13291 0.028
R13963 GND.n11351 GND.n11349 0.028
R13964 GND.n13506 GND.n13504 0.028
R13965 GND.n12094 GND.n12092 0.028
R13966 GND.n11926 GND.n11925 0.028
R13967 GND.n11910 GND.n11908 0.028
R13968 GND.n11816 GND.n11750 0.028
R13969 GND.n12196 GND.n12128 0.028
R13970 GND.n12297 GND.n12295 0.028
R13971 GND.n12313 GND.n12312 0.028
R13972 GND.n12478 GND.n12476 0.028
R13973 GND.n13193 GND.n13191 0.028
R13974 GND.n13031 GND.n13030 0.028
R13975 GND.n13015 GND.n13013 0.028
R13976 GND.n12919 GND.n12849 0.028
R13977 GND.n7686 GND.n7623 0.028
R13978 GND.n7786 GND.n7784 0.028
R13979 GND.n7802 GND.n7801 0.028
R13980 GND.n7961 GND.n7959 0.028
R13981 GND.n8191 GND.n8189 0.028
R13982 GND.n8280 GND.n8278 0.028
R13983 GND.n5874 GND.n5871 0.028
R13984 GND.n6003 GND.n6000 0.028
R13985 GND.n6442 GND.n6440 0.028
R13986 GND.n8147 GND.n8145 0.028
R13987 GND.n7986 GND.n7977 0.028
R13988 GND.n6995 GND.n6987 0.028
R13989 GND.n7157 GND.n7155 0.028
R13990 GND.n6915 GND.n6912 0.028
R13991 GND.n6680 GND.n6677 0.028
R13992 GND.n6739 GND.n6737 0.028
R13993 GND.n7463 GND.n7461 0.028
R13994 GND.n7555 GND.n7552 0.028
R13995 GND.n7373 GND.n7371 0.028
R13996 GND.n7213 GND.n7204 0.028
R13997 GND.n15939 GND.n15894 0.028
R13998 GND.n16063 GND.n16061 0.028
R13999 GND.n16070 GND.n16069 0.028
R14000 GND.n16230 GND.n16228 0.028
R14001 GND.n1170 GND.n1168 0.028
R14002 GND.n1011 GND.n1007 0.028
R14003 GND.n1001 GND.n999 0.028
R14004 GND.n886 GND.n834 0.028
R14005 GND.n9639 GND.n9594 0.028
R14006 GND.n9763 GND.n9761 0.028
R14007 GND.n9770 GND.n9769 0.028
R14008 GND.n9930 GND.n9928 0.028
R14009 GND.n1231 GND.n1190 0.028
R14010 GND.n1353 GND.n1351 0.028
R14011 GND.n1360 GND.n1359 0.028
R14012 GND.n1526 GND.n1524 0.028
R14013 GND.n10307 GND.n10305 0.028
R14014 GND.n10147 GND.n10138 0.028
R14015 GND.n8870 GND.n8868 0.028
R14016 GND.n8716 GND.n8707 0.028
R14017 GND.n8577 GND.n8575 0.028
R14018 GND.n8417 GND.n8408 0.028
R14019 GND.n9324 GND.n9322 0.028
R14020 GND.n1729 GND.n1727 0.028
R14021 GND.n9451 GND.n9449 0.028
R14022 GND.n1869 GND.n1866 0.028
R14023 GND.n8669 GND.n8666 0.028
R14024 GND.n10131 GND.n10129 0.028
R14025 GND.n9976 GND.n9967 0.028
R14026 GND.n8938 GND.n8893 0.028
R14027 GND.n9062 GND.n9060 0.028
R14028 GND.n9069 GND.n9068 0.028
R14029 GND.n9229 GND.n9227 0.028
R14030 GND.n4536 GND.n4534 0.028
R14031 GND.n4371 GND.n4367 0.028
R14032 GND.n4361 GND.n4359 0.028
R14033 GND.n4246 GND.n4194 0.028
R14034 GND.n2522 GND.n2520 0.028
R14035 GND.n3191 GND.n3184 0.028
R14036 GND.n3347 GND.n3345 0.028
R14037 GND.n3432 GND.n3430 0.028
R14038 GND.n2428 GND.n2426 0.028
R14039 GND.n2360 GND.n2358 0.028
R14040 GND.n5095 GND.n5093 0.028
R14041 GND.n4934 GND.n4925 0.028
R14042 GND.n5131 GND.n5129 0.028
R14043 GND.n2089 GND.n2087 0.028
R14044 GND.n2169 GND.n2167 0.028
R14045 GND.n2936 GND.n2933 0.028
R14046 GND.n4749 GND.n4747 0.028
R14047 GND.n4588 GND.n4579 0.028
R14048 GND.n2991 GND.n2983 0.028
R14049 GND.n3146 GND.n3144 0.028
R14050 GND.n10415 GND.n10407 0.028
R14051 GND.n10570 GND.n10568 0.028
R14052 GND.n15557 GND.n15549 0.028
R14053 GND.n15844 GND.n15841 0.028
R14054 GND.n15399 GND.n15396 0.028
R14055 GND.n14952 GND.n14950 0.028
R14056 GND.n15085 GND.n15082 0.028
R14057 GND.n15277 GND.n15275 0.028
R14058 GND.n3951 GND.n3949 0.028
R14059 GND.n3792 GND.n3788 0.028
R14060 GND.n3782 GND.n3780 0.028
R14061 GND.n3670 GND.n3621 0.028
R14062 GND.n5789 GND.n5787 0.028
R14063 GND.n5630 GND.n5626 0.028
R14064 GND.n5620 GND.n5618 0.028
R14065 GND.n5505 GND.n5453 0.028
R14066 GND.n10689 GND.n10688 0.028
R14067 GND.n14039 GND.n14037 0.028
R14068 GND.n3510 GND.n3508 0.028
R14069 GND.n4900 GND.n4899 0.028
R14070 GND.n10911 GND.n10909 0.028
R14071 GND.n10960 GND.n10958 0.028
R14072 GND.n12823 GND.n12822 0.028
R14073 GND.n11648 GND.n11647 0.028
R14074 GND.n13215 GND.n13213 0.028
R14075 GND.n11430 GND.n11429 0.028
R14076 GND.n6101 GND.n6100 0.028
R14077 GND.n5844 GND.n5843 0.028
R14078 GND.n5920 GND.n5918 0.028
R14079 GND.n6513 GND.n6512 0.028
R14080 GND.n6833 GND.n6831 0.028
R14081 GND.n6598 GND.n6596 0.028
R14082 GND.n6821 GND.n6820 0.028
R14083 GND.n6980 GND.n6979 0.028
R14084 GND.n9404 GND.n9403 0.028
R14085 GND.n1811 GND.n1810 0.028
R14086 GND.n2603 GND.n2602 0.028
R14087 GND.n2305 GND.n2303 0.028
R14088 GND.n5211 GND.n5210 0.028
R14089 GND.n15765 GND.n15763 0.028
R14090 GND.n15319 GND.n15317 0.028
R14091 GND.n14460 GND.n14459 0.028
R14092 GND.n15011 GND.n15009 0.028
R14093 GND.n16470 GND.n16469 0.028
R14094 GND.n16539 GND.n16537 0.028
R14095 GND.n16364 GND.n16362 0.028
R14096 GND.n16731 GND.n16730 0.028
R14097 GND.n16800 GND.n16798 0.028
R14098 GND.n16625 GND.n16623 0.028
R14099 GND.n16992 GND.n16991 0.028
R14100 GND.n17061 GND.n17059 0.028
R14101 GND.n16886 GND.n16884 0.028
R14102 GND.n17253 GND.n17252 0.028
R14103 GND.n17322 GND.n17320 0.028
R14104 GND.n17147 GND.n17145 0.028
R14105 GND.n17514 GND.n17513 0.028
R14106 GND.n17583 GND.n17581 0.028
R14107 GND.n17408 GND.n17406 0.028
R14108 GND.n1541 GND.n802 0.027
R14109 GND.n9543 GND.n9534 0.026
R14110 GND.n14527 GND.n14526 0.026
R14111 GND.n14518 GND.n14517 0.026
R14112 GND.n14513 GND.n14512 0.026
R14113 GND.n14512 GND.n14511 0.026
R14114 GND.n14708 GND.n14706 0.026
R14115 GND.n14546 GND.n14544 0.026
R14116 GND.n14556 GND.n14554 0.026
R14117 GND.n14560 GND.n14559 0.026
R14118 GND.n14563 GND.n14560 0.026
R14119 GND.n14393 GND.n14391 0.026
R14120 GND.n10588 GND.n10586 0.026
R14121 GND.n10673 GND.n10671 0.026
R14122 GND.n10681 GND.n10679 0.026
R14123 GND.n15521 GND.n15519 0.026
R14124 GND.n14054 GND.n14052 0.026
R14125 GND.n14047 GND.n14045 0.026
R14126 GND.n14135 GND.n14133 0.026
R14127 GND.n14145 GND.n14143 0.026
R14128 GND.n14149 GND.n14148 0.026
R14129 GND.n14152 GND.n14149 0.026
R14130 GND.n10705 GND.n10703 0.026
R14131 GND.n14188 GND.n14186 0.026
R14132 GND.n14198 GND.n14196 0.026
R14133 GND.n14202 GND.n14201 0.026
R14134 GND.n14205 GND.n14202 0.026
R14135 GND.n14227 GND.n14225 0.026
R14136 GND.n3607 GND.n3605 0.026
R14137 GND.n3526 GND.n3524 0.026
R14138 GND.n3518 GND.n3516 0.026
R14139 GND.n4800 GND.n4798 0.026
R14140 GND.n4884 GND.n4882 0.026
R14141 GND.n4892 GND.n4890 0.026
R14142 GND.n2738 GND.n2737 0.026
R14143 GND.n4052 GND.n4051 0.026
R14144 GND.n10799 GND.n10797 0.026
R14145 GND.n10807 GND.n10805 0.026
R14146 GND.n10866 GND.n10864 0.026
R14147 GND.n13898 GND.n13896 0.026
R14148 GND.n13906 GND.n13904 0.026
R14149 GND.n13985 GND.n13983 0.026
R14150 GND.n13857 GND.n13855 0.026
R14151 GND.n10926 GND.n10924 0.026
R14152 GND.n10919 GND.n10917 0.026
R14153 GND.n13736 GND.n13734 0.026
R14154 GND.n10975 GND.n10973 0.026
R14155 GND.n10968 GND.n10966 0.026
R14156 GND.n14010 GND.n14009 0.026
R14157 GND.n12723 GND.n12721 0.026
R14158 GND.n12807 GND.n12805 0.026
R14159 GND.n12815 GND.n12813 0.026
R14160 GND.n10782 GND.n10781 0.026
R14161 GND.n13882 GND.n13879 0.026
R14162 GND.n11460 GND.n11458 0.026
R14163 GND.n11468 GND.n11466 0.026
R14164 GND.n11711 GND.n11709 0.026
R14165 GND.n11520 GND.n11518 0.026
R14166 GND.n11528 GND.n11526 0.026
R14167 GND.n11607 GND.n11605 0.026
R14168 GND.n11099 GND.n11097 0.026
R14169 GND.n11632 GND.n11630 0.026
R14170 GND.n11640 GND.n11638 0.026
R14171 GND.n13312 GND.n13310 0.026
R14172 GND.n13230 GND.n13228 0.026
R14173 GND.n13223 GND.n13221 0.026
R14174 GND.n11332 GND.n11330 0.026
R14175 GND.n11414 GND.n11412 0.026
R14176 GND.n11422 GND.n11420 0.026
R14177 GND.n13520 GND.n13518 0.026
R14178 GND.n13542 GND.n13541 0.026
R14179 GND.n8172 GND.n8170 0.026
R14180 GND.n6085 GND.n6083 0.026
R14181 GND.n6093 GND.n6091 0.026
R14182 GND.n8261 GND.n8259 0.026
R14183 GND.n8346 GND.n8344 0.026
R14184 GND.n8354 GND.n8352 0.026
R14185 GND.n6395 GND.n6394 0.026
R14186 GND.n5892 GND.n5890 0.026
R14187 GND.n5929 GND.n5927 0.026
R14188 GND.n5937 GND.n5935 0.026
R14189 GND.n6021 GND.n6019 0.026
R14190 GND.n6505 GND.n6504 0.026
R14191 GND.n6498 GND.n6497 0.026
R14192 GND.n6423 GND.n6421 0.026
R14193 GND.n8248 GND.n8247 0.026
R14194 GND.n8159 GND.n5833 0.026
R14195 GND.n6842 GND.n6840 0.026
R14196 GND.n6850 GND.n6848 0.026
R14197 GND.n6933 GND.n6931 0.026
R14198 GND.n6607 GND.n6605 0.026
R14199 GND.n6615 GND.n6613 0.026
R14200 GND.n6698 GND.n6696 0.026
R14201 GND.n6720 GND.n6718 0.026
R14202 GND.n6805 GND.n6803 0.026
R14203 GND.n6813 GND.n6811 0.026
R14204 GND.n7444 GND.n7442 0.026
R14205 GND.n6555 GND.n6553 0.026
R14206 GND.n6563 GND.n6561 0.026
R14207 GND.n7573 GND.n7571 0.026
R14208 GND.n6964 GND.n6962 0.026
R14209 GND.n6972 GND.n6970 0.026
R14210 GND.n7195 GND.n7194 0.026
R14211 GND.n7173 GND.n7171 0.026
R14212 GND.n9305 GND.n9303 0.026
R14213 GND.n9388 GND.n9386 0.026
R14214 GND.n9396 GND.n9394 0.026
R14215 GND.n1710 GND.n1708 0.026
R14216 GND.n1795 GND.n1793 0.026
R14217 GND.n1803 GND.n1801 0.026
R14218 GND.n1668 GND.n1667 0.026
R14219 GND.n1659 GND.n1658 0.026
R14220 GND.n1654 GND.n1653 0.026
R14221 GND.n1653 GND.n1652 0.026
R14222 GND.n9432 GND.n9430 0.026
R14223 GND.n1610 GND.n1608 0.026
R14224 GND.n1620 GND.n1618 0.026
R14225 GND.n1624 GND.n1623 0.026
R14226 GND.n1627 GND.n1624 0.026
R14227 GND.n1887 GND.n1885 0.026
R14228 GND.n8687 GND.n8685 0.026
R14229 GND.n8610 GND.n8608 0.026
R14230 GND.n8602 GND.n8600 0.026
R14231 GND.n1581 GND.n1580 0.026
R14232 GND.n1686 GND.n1684 0.026
R14233 GND.n2503 GND.n2501 0.026
R14234 GND.n2587 GND.n2585 0.026
R14235 GND.n2595 GND.n2593 0.026
R14236 GND.n2243 GND.n2241 0.026
R14237 GND.n2253 GND.n2251 0.026
R14238 GND.n2257 GND.n2256 0.026
R14239 GND.n2260 GND.n2257 0.026
R14240 GND.n3413 GND.n3411 0.026
R14241 GND.n2214 GND.n2212 0.026
R14242 GND.n2224 GND.n2222 0.026
R14243 GND.n2228 GND.n2227 0.026
R14244 GND.n2231 GND.n2228 0.026
R14245 GND.n2622 GND.n2620 0.026
R14246 GND.n2341 GND.n2339 0.026
R14247 GND.n2325 GND.n2323 0.026
R14248 GND.n2313 GND.n2311 0.026
R14249 GND.n3175 GND.n3174 0.026
R14250 GND.n2479 GND.n2477 0.026
R14251 GND.n5112 GND.n5110 0.026
R14252 GND.n5195 GND.n5193 0.026
R14253 GND.n5203 GND.n5201 0.026
R14254 GND.n2030 GND.n2028 0.026
R14255 GND.n2040 GND.n2038 0.026
R14256 GND.n2044 GND.n2043 0.026
R14257 GND.n2047 GND.n2044 0.026
R14258 GND.n2070 GND.n2068 0.026
R14259 GND.n1977 GND.n1975 0.026
R14260 GND.n1987 GND.n1985 0.026
R14261 GND.n1991 GND.n1990 0.026
R14262 GND.n1994 GND.n1991 0.026
R14263 GND.n2649 GND.n2647 0.026
R14264 GND.n2954 GND.n2952 0.026
R14265 GND.n2872 GND.n2870 0.026
R14266 GND.n2864 GND.n2862 0.026
R14267 GND.n2669 GND.n2668 0.026
R14268 GND.n4918 GND.n4917 0.026
R14269 GND.n14084 GND.n14082 0.026
R14270 GND.n15545 GND.n15544 0.026
R14271 GND.n15750 GND.n15749 0.026
R14272 GND.n15728 GND.n15726 0.026
R14273 GND.n15862 GND.n15860 0.026
R14274 GND.n15780 GND.n15778 0.026
R14275 GND.n15773 GND.n15771 0.026
R14276 GND.n15417 GND.n15415 0.026
R14277 GND.n15334 GND.n15332 0.026
R14278 GND.n15327 GND.n15325 0.026
R14279 GND.n14933 GND.n14931 0.026
R14280 GND.n14444 GND.n14442 0.026
R14281 GND.n14452 GND.n14450 0.026
R14282 GND.n14489 GND.n14488 0.026
R14283 GND.n15447 GND.n15439 0.026
R14284 GND.n15103 GND.n15101 0.026
R14285 GND.n15026 GND.n15024 0.026
R14286 GND.n15019 GND.n15017 0.026
R14287 GND.n14722 GND.n14719 0.026
R14288 GND.n16353 GND.n16351 0.026
R14289 GND.n16614 GND.n16612 0.026
R14290 GND.n16875 GND.n16873 0.026
R14291 GND.n17136 GND.n17134 0.026
R14292 GND.n17397 GND.n17395 0.026
R14293 GND.n640 GND.n638 0.026
R14294 GND.n742 GND.n740 0.026
R14295 GND.n574 GND.n572 0.026
R14296 GND.n382 GND.n380 0.026
R14297 GND.n484 GND.n482 0.026
R14298 GND.n316 GND.n314 0.026
R14299 GND.n124 GND.n122 0.026
R14300 GND.n226 GND.n224 0.026
R14301 GND.n58 GND.n56 0.026
R14302 GND.n17739 GND.n17737 0.026
R14303 GND.n17815 GND.n17813 0.026
R14304 GND.n17894 GND.n17892 0.026
R14305 GND.n5338 GND.n5337 0.026
R14306 GND.n652 GND.n650 0.026
R14307 GND.n755 GND.n753 0.026
R14308 GND.n587 GND.n585 0.026
R14309 GND.n394 GND.n392 0.026
R14310 GND.n497 GND.n495 0.026
R14311 GND.n329 GND.n327 0.026
R14312 GND.n136 GND.n134 0.026
R14313 GND.n239 GND.n237 0.026
R14314 GND.n71 GND.n69 0.026
R14315 GND.n17751 GND.n17749 0.026
R14316 GND.n17828 GND.n17826 0.026
R14317 GND.n17907 GND.n17905 0.026
R14318 GND.n697 GND.n696 0.025
R14319 GND.n724 GND.n723 0.025
R14320 GND.n439 GND.n438 0.025
R14321 GND.n466 GND.n465 0.025
R14322 GND.n181 GND.n180 0.025
R14323 GND.n208 GND.n207 0.025
R14324 GND.n17796 GND.n17795 0.025
R14325 GND.n17718 GND.n17717 0.025
R14326 GND.n17860 GND.n17859 0.025
R14327 GND.n14863 GND.n14861 0.025
R14328 GND.n14792 GND.n14790 0.025
R14329 GND.n6283 GND.n6281 0.025
R14330 GND.n6215 GND.n6213 0.025
R14331 GND.n12651 GND.n12649 0.025
R14332 GND.n12580 GND.n12578 0.025
R14333 GND.n11264 GND.n11262 0.025
R14334 GND.n11196 GND.n11194 0.025
R14335 GND.n13671 GND.n13669 0.025
R14336 GND.n13603 GND.n13601 0.025
R14337 GND.n13387 GND.n13385 0.025
R14338 GND.n13458 GND.n13456 0.025
R14339 GND.n11987 GND.n11985 0.025
R14340 GND.n11945 GND.n11943 0.025
R14341 GND.n11893 GND.n11891 0.025
R14342 GND.n11857 GND.n11855 0.025
R14343 GND.n12237 GND.n12235 0.025
R14344 GND.n12279 GND.n12277 0.025
R14345 GND.n12330 GND.n12329 0.025
R14346 GND.n12368 GND.n12366 0.025
R14347 GND.n13092 GND.n13090 0.025
R14348 GND.n13050 GND.n13048 0.025
R14349 GND.n12998 GND.n12996 0.025
R14350 GND.n12961 GND.n12959 0.025
R14351 GND.n7726 GND.n7724 0.025
R14352 GND.n7768 GND.n7766 0.025
R14353 GND.n7819 GND.n7818 0.025
R14354 GND.n7856 GND.n7854 0.025
R14355 GND.n8099 GND.n8097 0.025
R14356 GND.n8028 GND.n8026 0.025
R14357 GND.n7037 GND.n7035 0.025
R14358 GND.n7108 GND.n7106 0.025
R14359 GND.n7326 GND.n7324 0.025
R14360 GND.n7254 GND.n7252 0.025
R14361 GND.n15980 GND.n15978 0.025
R14362 GND.n16033 GND.n16031 0.025
R14363 GND.n16087 GND.n16086 0.025
R14364 GND.n16142 GND.n16140 0.025
R14365 GND.n1091 GND.n1089 0.025
R14366 GND.n1039 GND.n1037 0.025
R14367 GND.n984 GND.n982 0.025
R14368 GND.n928 GND.n926 0.025
R14369 GND.n9680 GND.n9678 0.025
R14370 GND.n9733 GND.n9731 0.025
R14371 GND.n9787 GND.n9786 0.025
R14372 GND.n9842 GND.n9840 0.025
R14373 GND.n1271 GND.n1269 0.025
R14374 GND.n1323 GND.n1321 0.025
R14375 GND.n1377 GND.n1376 0.025
R14376 GND.n1434 GND.n1432 0.025
R14377 GND.n10260 GND.n10258 0.025
R14378 GND.n10188 GND.n10186 0.025
R14379 GND.n8824 GND.n8822 0.025
R14380 GND.n8756 GND.n8754 0.025
R14381 GND.n8530 GND.n8528 0.025
R14382 GND.n8458 GND.n8456 0.025
R14383 GND.n10085 GND.n10083 0.025
R14384 GND.n10017 GND.n10015 0.025
R14385 GND.n8979 GND.n8977 0.025
R14386 GND.n9032 GND.n9030 0.025
R14387 GND.n9086 GND.n9085 0.025
R14388 GND.n9141 GND.n9139 0.025
R14389 GND.n4452 GND.n4450 0.025
R14390 GND.n4399 GND.n4397 0.025
R14391 GND.n4344 GND.n4342 0.025
R14392 GND.n4288 GND.n4286 0.025
R14393 GND.n3231 GND.n3229 0.025
R14394 GND.n3299 GND.n3297 0.025
R14395 GND.n5047 GND.n5045 0.025
R14396 GND.n4976 GND.n4974 0.025
R14397 GND.n3385 GND.n3382 0.025
R14398 GND.n4787 GND.n4784 0.025
R14399 GND.n4701 GND.n4699 0.025
R14400 GND.n4630 GND.n4628 0.025
R14401 GND.n3031 GND.n3029 0.025
R14402 GND.n3099 GND.n3097 0.025
R14403 GND.n10455 GND.n10453 0.025
R14404 GND.n10523 GND.n10521 0.025
R14405 GND.n15599 GND.n15597 0.025
R14406 GND.n15670 GND.n15668 0.025
R14407 GND.n15162 GND.n15160 0.025
R14408 GND.n15230 GND.n15228 0.025
R14409 GND.n3872 GND.n3870 0.025
R14410 GND.n3820 GND.n3818 0.025
R14411 GND.n3765 GND.n3763 0.025
R14412 GND.n3711 GND.n3709 0.025
R14413 GND.n5710 GND.n5708 0.025
R14414 GND.n5658 GND.n5656 0.025
R14415 GND.n5603 GND.n5601 0.025
R14416 GND.n5547 GND.n5545 0.025
R14417 GND.n16425 GND.n16424 0.024
R14418 GND.n16503 GND.n16502 0.024
R14419 GND.n16686 GND.n16685 0.024
R14420 GND.n16764 GND.n16763 0.024
R14421 GND.n16947 GND.n16946 0.024
R14422 GND.n17025 GND.n17024 0.024
R14423 GND.n17208 GND.n17207 0.024
R14424 GND.n17286 GND.n17285 0.024
R14425 GND.n17469 GND.n17468 0.024
R14426 GND.n17547 GND.n17546 0.024
R14427 GND.n14498 GND.n14497 0.024
R14428 GND.n14697 GND.n14694 0.024
R14429 GND.n14371 GND.n14369 0.024
R14430 GND.n10600 GND.n10598 0.024
R14431 GND.n15510 GND.n15507 0.024
R14432 GND.n14127 GND.n14126 0.024
R14433 GND.n14322 GND.n14320 0.024
R14434 GND.n14169 GND.n14168 0.024
R14435 GND.n14239 GND.n14237 0.024
R14436 GND.n3596 GND.n3593 0.024
R14437 GND.n4812 GND.n4810 0.024
R14438 GND.n2751 GND.n2743 0.024
R14439 GND.n4070 GND.n4060 0.024
R14440 GND.n10790 GND.n10788 0.024
R14441 GND.n10855 GND.n10852 0.024
R14442 GND.n13890 GND.n13888 0.024
R14443 GND.n13974 GND.n13971 0.024
R14444 GND.n13846 GND.n13843 0.024
R14445 GND.n13748 GND.n13746 0.024
R14446 GND.n12735 GND.n12733 0.024
R14447 GND.n11451 GND.n11449 0.024
R14448 GND.n11700 GND.n11697 0.024
R14449 GND.n11512 GND.n11510 0.024
R14450 GND.n11596 GND.n11593 0.024
R14451 GND.n11088 GND.n11085 0.024
R14452 GND.n13301 GND.n13298 0.024
R14453 GND.n11344 GND.n11342 0.024
R14454 GND.n11137 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE 0.024
R14455 GND.n8184 GND.n8182 0.024
R14456 GND.n8273 GND.n8271 0.024
R14457 GND.n8362 GND.n8361 0.024
R14458 GND.n5881 GND.n5878 0.024
R14459 GND.n6010 GND.n6007 0.024
R14460 GND.n6435 GND.n6433 0.024
R14461 GND.n6922 GND.n6919 0.024
R14462 GND.n6687 GND.n6684 0.024
R14463 GND.n6732 GND.n6730 0.024
R14464 GND.n7456 GND.n7454 0.024
R14465 GND.n6571 GND.n6570 0.024
R14466 GND.n7562 GND.n7559 0.024
R14467 GND.n9317 GND.n9315 0.024
R14468 GND.n1722 GND.n1720 0.024
R14469 GND.n1676 GND.n1674 0.024
R14470 GND.n9444 GND.n9442 0.024
R14471 GND.n1590 GND.n1589 0.024
R14472 GND.n1876 GND.n1873 0.024
R14473 GND.n8676 GND.n8673 0.024
R14474 GND.n8594 GND.n8592 0.024
R14475 GND.n2515 GND.n2513 0.024
R14476 GND.n2469 GND.n2467 0.024
R14477 GND.n3425 GND.n3423 0.024
R14478 GND.n2203 GND.n2201 0.024
R14479 GND.n2353 GND.n2351 0.024
R14480 GND.n5124 GND.n5122 0.024
R14481 GND.n2011 GND.n2010 0.024
R14482 GND.n2082 GND.n2080 0.024
R14483 GND.n1968 GND.n1967 0.024
R14484 GND.n2943 GND.n2940 0.024
R14485 GND.n2856 GND.n2854 0.024
R14486 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/GATE GND.n4781 0.024
R14487 GND.n14111 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/GATE 0.024
R14488 GND.n15851 GND.n15848 0.024
R14489 GND.n15406 GND.n15403 0.024
R14490 GND.n14945 GND.n14943 0.024
R14491 GND.n15092 GND.n15089 0.024
R14492 GND.n16333 GND.n16332 0.024
R14493 GND.n16594 GND.n16593 0.024
R14494 GND.n16855 GND.n16854 0.024
R14495 GND.n17116 GND.n17115 0.024
R14496 GND.n17377 GND.n17376 0.024
R14497 GND.n691 GND.n689 0.024
R14498 GND.n563 GND.n562 0.024
R14499 GND.n556 GND.n555 0.024
R14500 GND.n433 GND.n431 0.024
R14501 GND.n305 GND.n304 0.024
R14502 GND.n298 GND.n297 0.024
R14503 GND.n175 GND.n173 0.024
R14504 GND.n47 GND.n46 0.024
R14505 GND.n40 GND.n39 0.024
R14506 GND.n17790 GND.n17788 0.024
R14507 GND.n17883 GND.n17882 0.024
R14508 GND.n17876 GND.n17875 0.024
R14509 GND.n3364 GND.n3361 0.024
R14510 GND.n14899 GND.n14897 0.023
R14511 GND.n14763 GND.n14754 0.023
R14512 GND.n6317 GND.n6315 0.023
R14513 GND.n6187 GND.n6178 0.023
R14514 GND.n12687 GND.n12685 0.023
R14515 GND.n12551 GND.n12542 0.023
R14516 GND.n11298 GND.n11296 0.023
R14517 GND.n11168 GND.n11160 0.023
R14518 GND.n13705 GND.n13703 0.023
R14519 GND.n13575 GND.n13567 0.023
R14520 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE GND.n10898 0.023
R14521 GND.n13358 GND.n13349 0.023
R14522 GND.n13494 GND.n13492 0.023
R14523 GND.n12022 GND.n12020 0.023
R14524 GND.n11931 GND.n11930 0.023
R14525 GND.n11905 GND.n11903 0.023
R14526 GND.n11828 GND.n11820 0.023
R14527 GND.n12208 GND.n12200 0.023
R14528 GND.n12292 GND.n12290 0.023
R14529 GND.n12318 GND.n12317 0.023
R14530 GND.n12404 GND.n12402 0.023
R14531 GND.n13126 GND.n13124 0.023
R14532 GND.n13036 GND.n13035 0.023
R14533 GND.n13010 GND.n13008 0.023
R14534 GND.n12932 GND.n12923 0.023
R14535 GND.n7698 GND.n7690 0.023
R14536 GND.n7781 GND.n7779 0.023
R14537 GND.n7807 GND.n7806 0.023
R14538 GND.n7891 GND.n7889 0.023
R14539 GND.n8135 GND.n8133 0.023
R14540 GND.n7999 GND.n7990 0.023
R14541 GND.n7008 GND.n6999 0.023
R14542 GND.n7144 GND.n7142 0.023
R14543 GND.n7361 GND.n7359 0.023
R14544 GND.n7225 GND.n7217 0.023
R14545 GND.n15951 GND.n15943 0.023
R14546 GND.n16055 GND.n16053 0.023
R14547 GND.n16075 GND.n16074 0.023
R14548 GND.n16177 GND.n16175 0.023
R14549 GND.n1125 GND.n1123 0.023
R14550 GND.n1019 GND.n1015 0.023
R14551 GND.n996 GND.n994 0.023
R14552 GND.n899 GND.n890 0.023
R14553 GND.n9651 GND.n9643 0.023
R14554 GND.n9755 GND.n9753 0.023
R14555 GND.n9775 GND.n9774 0.023
R14556 GND.n9877 GND.n9875 0.023
R14557 GND.n1243 GND.n1235 0.023
R14558 GND.n1345 GND.n1343 0.023
R14559 GND.n1365 GND.n1364 0.023
R14560 GND.n1470 GND.n1468 0.023
R14561 GND.n10295 GND.n10293 0.023
R14562 GND.n10159 GND.n10151 0.023
R14563 GND.n8858 GND.n8856 0.023
R14564 GND.n8728 GND.n8720 0.023
R14565 GND.n8565 GND.n8563 0.023
R14566 GND.n8429 GND.n8421 0.023
R14567 GND.n10119 GND.n10117 0.023
R14568 GND.n9989 GND.n9980 0.023
R14569 GND.n8950 GND.n8942 0.023
R14570 GND.n9054 GND.n9052 0.023
R14571 GND.n9074 GND.n9073 0.023
R14572 GND.n9176 GND.n9174 0.023
R14573 GND.n4487 GND.n4485 0.023
R14574 GND.n4379 GND.n4375 0.023
R14575 GND.n4356 GND.n4354 0.023
R14576 GND.n4259 GND.n4250 0.023
R14577 GND.n3203 GND.n3195 0.023
R14578 GND.n3334 GND.n3332 0.023
R14579 GND.n5083 GND.n5081 0.023
R14580 GND.n4947 GND.n4938 0.023
R14581 GND.n3393 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/GATE 0.023
R14582 GND.n4737 GND.n4735 0.023
R14583 GND.n4601 GND.n4592 0.023
R14584 GND.n3003 GND.n2995 0.023
R14585 GND.n3134 GND.n3132 0.023
R14586 GND.n10427 GND.n10419 0.023
R14587 GND.n10557 GND.n10555 0.023
R14588 GND.n15570 GND.n15561 0.023
R14589 GND.n15706 GND.n15704 0.023
R14590 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/GATE GND.n15305 0.023
R14591 GND.n15134 GND.n15126 0.023
R14592 GND.n15265 GND.n15263 0.023
R14593 GND.n3906 GND.n3904 0.023
R14594 GND.n3800 GND.n3796 0.023
R14595 GND.n3777 GND.n3775 0.023
R14596 GND.n3683 GND.n3674 0.023
R14597 GND.n5744 GND.n5742 0.023
R14598 GND.n5638 GND.n5634 0.023
R14599 GND.n5615 GND.n5613 0.023
R14600 GND.n5518 GND.n5509 0.023
R14601 GND.n5366 GND.n5365 0.023
R14602 GND.n16426 GND.n16425 0.023
R14603 GND.n16502 GND.n16501 0.023
R14604 GND.n16687 GND.n16686 0.023
R14605 GND.n16763 GND.n16762 0.023
R14606 GND.n16948 GND.n16947 0.023
R14607 GND.n17024 GND.n17023 0.023
R14608 GND.n17209 GND.n17208 0.023
R14609 GND.n17285 GND.n17284 0.023
R14610 GND.n17470 GND.n17469 0.023
R14611 GND.n17546 GND.n17545 0.023
R14612 GND.n696 GND.n695 0.022
R14613 GND.n723 GND.n722 0.022
R14614 GND.n438 GND.n437 0.022
R14615 GND.n465 GND.n464 0.022
R14616 GND.n180 GND.n179 0.022
R14617 GND.n207 GND.n206 0.022
R14618 GND.n17795 GND.n17794 0.022
R14619 GND.n17717 GND.n17716 0.022
R14620 GND.n9533 GND.n9532 0.022
R14621 GND.n3379 GND.n3376 0.022
R14622 GND.n12829 GND.n12532 0.021
R14623 GND.n14001 GND.n14000 0.021
R14624 GND.n13330 GND.n13329 0.021
R14625 GND.n11319 GND.n11145 0.021
R14626 GND.n3361 GND.n3356 0.021
R14627 GND.n5217 GND.n1924 0.021
R14628 GND.n2969 GND.n2968 0.021
R14629 GND.n4766 GND.n4761 0.021
R14630 GND.n15872 GND.n10400 0.021
R14631 GND.n15536 GND.n15535 0.021
R14632 GND.n14728 GND.n14727 0.021
R14633 GND.n15291 GND.n15286 0.021
R14634 GND.n14655 GND.n14654 0.021
R14635 GND.n14701 GND.n14699 0.021
R14636 GND.n14589 GND.n14588 0.021
R14637 GND.n14386 GND.n14384 0.021
R14638 GND.n10595 GND.n10593 0.021
R14639 GND.n10644 GND.n10637 0.021
R14640 GND.n15514 GND.n15512 0.021
R14641 GND.n15470 GND.n15469 0.021
R14642 GND.n14314 GND.n14313 0.021
R14643 GND.n10698 GND.n10696 0.021
R14644 GND.n14278 GND.n14277 0.021
R14645 GND.n14234 GND.n14232 0.021
R14646 GND.n14876 GND.n14874 0.021
R14647 GND.n14779 GND.n14777 0.021
R14648 GND.n3600 GND.n3598 0.021
R14649 GND.n3556 GND.n3555 0.021
R14650 GND.n4807 GND.n4805 0.021
R14651 GND.n4855 GND.n4849 0.021
R14652 GND.n6295 GND.n6293 0.021
R14653 GND.n6203 GND.n6201 0.021
R14654 GND.n12664 GND.n12662 0.021
R14655 GND.n12567 GND.n12565 0.021
R14656 GND.n10769 GND.n10768 0.021
R14657 GND.n10859 GND.n10857 0.021
R14658 GND.n13933 GND.n13932 0.021
R14659 GND.n13978 GND.n13976 0.021
R14660 GND.n13850 GND.n13848 0.021
R14661 GND.n13806 GND.n13805 0.021
R14662 GND.n13743 GND.n13741 0.021
R14663 GND.n13789 GND.n13784 0.021
R14664 GND.n11276 GND.n11274 0.021
R14665 GND.n11184 GND.n11182 0.021
R14666 GND.n13683 GND.n13681 0.021
R14667 GND.n13591 GND.n13589 0.021
R14668 GND.n10904 GND.n10901 0.021
R14669 GND.n12730 GND.n12728 0.021
R14670 GND.n12778 GND.n12772 0.021
R14671 GND.n11659 GND.n11658 0.021
R14672 GND.n11704 GND.n11702 0.021
R14673 GND.n11555 GND.n11554 0.021
R14674 GND.n11600 GND.n11598 0.021
R14675 GND.n11092 GND.n11090 0.021
R14676 GND.n11048 GND.n11047 0.021
R14677 GND.n13305 GND.n13303 0.021
R14678 GND.n13261 GND.n13260 0.021
R14679 GND.n11339 GND.n11337 0.021
R14680 GND.n11385 GND.n11380 0.021
R14681 GND.n13374 GND.n13372 0.021
R14682 GND.n13471 GND.n13469 0.021
R14683 GND.n11129 GND.n11126 0.021
R14684 GND.n11999 GND.n11997 0.021
R14685 GND.n11940 GND.n11938 0.021
R14686 GND.n11897 GND.n11895 0.021
R14687 GND.n11845 GND.n11843 0.021
R14688 GND.n12225 GND.n12223 0.021
R14689 GND.n12284 GND.n12282 0.021
R14690 GND.n12326 GND.n12325 0.021
R14691 GND.n12381 GND.n12379 0.021
R14692 GND.n13104 GND.n13102 0.021
R14693 GND.n13045 GND.n13043 0.021
R14694 GND.n13002 GND.n13000 0.021
R14695 GND.n12948 GND.n12946 0.021
R14696 GND.n7714 GND.n7712 0.021
R14697 GND.n7773 GND.n7771 0.021
R14698 GND.n7815 GND.n7814 0.021
R14699 GND.n7868 GND.n7866 0.021
R14700 GND.n8179 GND.n8177 0.021
R14701 GND.n8226 GND.n8221 0.021
R14702 GND.n8268 GND.n8266 0.021
R14703 GND.n8317 GND.n8310 0.021
R14704 GND.n5885 GND.n5883 0.021
R14705 GND.n5969 GND.n5968 0.021
R14706 GND.n6014 GND.n6012 0.021
R14707 GND.n6472 GND.n6471 0.021
R14708 GND.n6430 GND.n6428 0.021
R14709 GND.n8112 GND.n8110 0.021
R14710 GND.n8015 GND.n8013 0.021
R14711 GND.n6050 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE 0.021
R14712 GND.n7024 GND.n7022 0.021
R14713 GND.n7121 GND.n7119 0.021
R14714 GND.n6881 GND.n6880 0.021
R14715 GND.n6926 GND.n6924 0.021
R14716 GND.n6646 GND.n6645 0.021
R14717 GND.n6691 GND.n6689 0.021
R14718 GND.n6727 GND.n6725 0.021
R14719 GND.n6776 GND.n6769 0.021
R14720 GND.n7451 GND.n7449 0.021
R14721 GND.n7499 GND.n7493 0.021
R14722 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE GND.n7397 0.021
R14723 GND.n7566 GND.n7564 0.021
R14724 GND.n7522 GND.n7521 0.021
R14725 GND.n7338 GND.n7336 0.021
R14726 GND.n7242 GND.n7240 0.021
R14727 GND.n15968 GND.n15966 0.021
R14728 GND.n16041 GND.n16039 0.021
R14729 GND.n16083 GND.n16082 0.021
R14730 GND.n16154 GND.n16152 0.021
R14731 GND.n1103 GND.n1101 0.021
R14732 GND.n1031 GND.n1029 0.021
R14733 GND.n988 GND.n986 0.021
R14734 GND.n915 GND.n913 0.021
R14735 GND.n9668 GND.n9666 0.021
R14736 GND.n9741 GND.n9739 0.021
R14737 GND.n9783 GND.n9782 0.021
R14738 GND.n9854 GND.n9852 0.021
R14739 GND.n1259 GND.n1257 0.021
R14740 GND.n1331 GND.n1329 0.021
R14741 GND.n1373 GND.n1372 0.021
R14742 GND.n1447 GND.n1445 0.021
R14743 GND.n10272 GND.n10270 0.021
R14744 GND.n10176 GND.n10174 0.021
R14745 GND.n8836 GND.n8834 0.021
R14746 GND.n8744 GND.n8742 0.021
R14747 GND.n8542 GND.n8540 0.021
R14748 GND.n8446 GND.n8444 0.021
R14749 GND.n9312 GND.n9310 0.021
R14750 GND.n9359 GND.n9354 0.021
R14751 GND.n1717 GND.n1715 0.021
R14752 GND.n1766 GND.n1759 0.021
R14753 GND.n9483 GND.n9482 0.021
R14754 GND.n9439 GND.n9437 0.021
R14755 GND.n1834 GND.n1833 0.021
R14756 GND.n1880 GND.n1878 0.021
R14757 GND.n8680 GND.n8678 0.021
R14758 GND.n8636 GND.n8635 0.021
R14759 GND.n10097 GND.n10095 0.021
R14760 GND.n10005 GND.n10003 0.021
R14761 GND.n9281 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE 0.021
R14762 GND.n8967 GND.n8965 0.021
R14763 GND.n9040 GND.n9038 0.021
R14764 GND.n9082 GND.n9081 0.021
R14765 GND.n9153 GND.n9151 0.021
R14766 GND.n4464 GND.n4462 0.021
R14767 GND.n4391 GND.n4389 0.021
R14768 GND.n4348 GND.n4346 0.021
R14769 GND.n4275 GND.n4273 0.021
R14770 GND.n2510 GND.n2508 0.021
R14771 GND.n2558 GND.n2552 0.021
R14772 GND.n3219 GND.n3217 0.021
R14773 GND.n3311 GND.n3309 0.021
R14774 GND.n3464 GND.n3463 0.021
R14775 GND.n3420 GND.n3418 0.021
R14776 GND.n2416 GND.n2415 0.021
R14777 GND.n2615 GND.n2613 0.021
R14778 GND.n2348 GND.n2346 0.021
R14779 GND.n5060 GND.n5058 0.021
R14780 GND.n4963 GND.n4961 0.021
R14781 GND.n3366 GND.n3364 0.021
R14782 GND.n5226 GND.n5225 0.021
R14783 GND.n5119 GND.n5117 0.021
R14784 GND.n5166 GND.n5161 0.021
R14785 GND.n2121 GND.n2120 0.021
R14786 GND.n2077 GND.n2075 0.021
R14787 GND.n2157 GND.n2156 0.021
R14788 GND.n2642 GND.n2640 0.021
R14789 GND.n2947 GND.n2945 0.021
R14790 GND.n2903 GND.n2902 0.021
R14791 GND.n1959 GND.n1957 0.021
R14792 GND.n4757 GND.n4752 0.021
R14793 GND.n4714 GND.n4712 0.021
R14794 GND.n4617 GND.n4615 0.021
R14795 GND.n3019 GND.n3017 0.021
R14796 GND.n3111 GND.n3109 0.021
R14797 GND.n10443 GND.n10441 0.021
R14798 GND.n10535 GND.n10533 0.021
R14799 GND.n14103 GND.n14100 0.021
R14800 GND.n15586 GND.n15584 0.021
R14801 GND.n15683 GND.n15681 0.021
R14802 GND.n15855 GND.n15853 0.021
R14803 GND.n15811 GND.n15810 0.021
R14804 GND.n15410 GND.n15408 0.021
R14805 GND.n15366 GND.n15365 0.021
R14806 GND.n14940 GND.n14938 0.021
R14807 GND.n14987 GND.n14981 0.021
R14808 GND.n15096 GND.n15094 0.021
R14809 GND.n15052 GND.n15051 0.021
R14810 GND.n15312 GND.n15308 0.021
R14811 GND.n15150 GND.n15148 0.021
R14812 GND.n15242 GND.n15240 0.021
R14813 GND.n3884 GND.n3882 0.021
R14814 GND.n3812 GND.n3810 0.021
R14815 GND.n3769 GND.n3767 0.021
R14816 GND.n3699 GND.n3697 0.021
R14817 GND.n5722 GND.n5720 0.021
R14818 GND.n5650 GND.n5648 0.021
R14819 GND.n5607 GND.n5605 0.021
R14820 GND.n5534 GND.n5532 0.021
R14821 GND.n16451 GND.n16447 0.021
R14822 GND.n16565 GND.n16561 0.021
R14823 GND.n16391 GND.n16387 0.021
R14824 GND.n16330 GND.n16329 0.021
R14825 GND.n16712 GND.n16708 0.021
R14826 GND.n16826 GND.n16822 0.021
R14827 GND.n16652 GND.n16648 0.021
R14828 GND.n16591 GND.n16590 0.021
R14829 GND.n16973 GND.n16969 0.021
R14830 GND.n17087 GND.n17083 0.021
R14831 GND.n16913 GND.n16909 0.021
R14832 GND.n16852 GND.n16851 0.021
R14833 GND.n17234 GND.n17230 0.021
R14834 GND.n17348 GND.n17344 0.021
R14835 GND.n17174 GND.n17170 0.021
R14836 GND.n17113 GND.n17112 0.021
R14837 GND.n17495 GND.n17491 0.021
R14838 GND.n17609 GND.n17605 0.021
R14839 GND.n17435 GND.n17431 0.021
R14840 GND.n17374 GND.n17373 0.021
R14841 GND.n678 GND.n674 0.021
R14842 GND.n781 GND.n777 0.021
R14843 GND.n612 GND.n608 0.021
R14844 GND.n420 GND.n416 0.021
R14845 GND.n523 GND.n519 0.021
R14846 GND.n354 GND.n350 0.021
R14847 GND.n162 GND.n158 0.021
R14848 GND.n265 GND.n261 0.021
R14849 GND.n96 GND.n92 0.021
R14850 GND.n17777 GND.n17773 0.021
R14851 GND.n17854 GND.n17850 0.021
R14852 GND.n17932 GND.n17928 0.021
R14853 GND.n6117 GND.n6116 0.021
R14854 GND.n7583 GND.n6154 0.021
R14855 GND.n9414 GND.n9409 0.021
R14856 GND.n17803 GND.n17802 0.021
R14857 GND.n567 GND.n566 0.021
R14858 GND.n309 GND.n308 0.021
R14859 GND.n51 GND.n50 0.021
R14860 GND.n17887 GND.n17886 0.021
R14861 GND.n16529 GND.n16528 0.019
R14862 GND.n16482 GND.n16442 0.019
R14863 GND.n16790 GND.n16789 0.019
R14864 GND.n16743 GND.n16703 0.019
R14865 GND.n17051 GND.n17050 0.019
R14866 GND.n17004 GND.n16964 0.019
R14867 GND.n17312 GND.n17311 0.019
R14868 GND.n17265 GND.n17225 0.019
R14869 GND.n17573 GND.n17572 0.019
R14870 GND.n17526 GND.n17486 0.019
R14871 GND.n5351 GND.n5350 0.019
R14872 GND.n14526 GND.n14524 0.019
R14873 GND.n14648 GND.n14646 0.019
R14874 GND.n14657 GND.n14655 0.019
R14875 GND.n14661 GND.n14660 0.019
R14876 GND.n14704 GND.n14701 0.019
R14877 GND.n14547 GND.n14546 0.019
R14878 GND.n14582 GND.n14580 0.019
R14879 GND.n14627 GND.n14626 0.019
R14880 GND.n14389 GND.n14386 0.019
R14881 GND.n10593 GND.n10591 0.019
R14882 GND.n10637 GND.n10636 0.019
R14883 GND.n10649 GND.n10647 0.019
R14884 GND.n15517 GND.n15514 0.019
R14885 GND.n15472 GND.n15470 0.019
R14886 GND.n14077 GND.n14076 0.019
R14887 GND.n14136 GND.n14135 0.019
R14888 GND.n14305 GND.n14303 0.019
R14889 GND.n14355 GND.n14354 0.019
R14890 GND.n10701 GND.n10698 0.019
R14891 GND.n14189 GND.n14188 0.019
R14892 GND.n14283 GND.n14281 0.019
R14893 GND.n14277 GND.n14276 0.019
R14894 GND.n14272 GND.n14271 0.019
R14895 GND.n14232 GND.n14230 0.019
R14896 GND.n14886 GND.n14884 0.019
R14897 GND.n14775 GND.n14767 0.019
R14898 GND.n3603 GND.n3600 0.019
R14899 GND.n3558 GND.n3556 0.019
R14900 GND.n3549 GND.n3548 0.019
R14901 GND.n4805 GND.n4803 0.019
R14902 GND.n4849 GND.n4848 0.019
R14903 GND.n4860 GND.n4858 0.019
R14904 GND.n6305 GND.n6303 0.019
R14905 GND.n6199 GND.n6191 0.019
R14906 GND.n12674 GND.n12672 0.019
R14907 GND.n12563 GND.n12555 0.019
R14908 GND.n10831 GND.n10829 0.019
R14909 GND.n10768 GND.n10767 0.019
R14910 GND.n10862 GND.n10859 0.019
R14911 GND.n13930 GND.n13928 0.019
R14912 GND.n13935 GND.n13933 0.019
R14913 GND.n13981 GND.n13978 0.019
R14914 GND.n13853 GND.n13850 0.019
R14915 GND.n13808 GND.n13806 0.019
R14916 GND.n10949 GND.n10948 0.019
R14917 GND.n13741 GND.n13739 0.019
R14918 GND.n13784 GND.n13783 0.019
R14919 GND.n10998 GND.n10997 0.019
R14920 GND.n11286 GND.n11284 0.019
R14921 GND.n11180 GND.n11172 0.019
R14922 GND.n13693 GND.n13691 0.019
R14923 GND.n13587 GND.n13579 0.019
R14924 GND.n12728 GND.n12726 0.019
R14925 GND.n12772 GND.n12771 0.019
R14926 GND.n12783 GND.n12781 0.019
R14927 GND.n11492 GND.n11490 0.019
R14928 GND.n11661 GND.n11659 0.019
R14929 GND.n11707 GND.n11704 0.019
R14930 GND.n11552 GND.n11550 0.019
R14931 GND.n11557 GND.n11555 0.019
R14932 GND.n11603 GND.n11600 0.019
R14933 GND.n11095 GND.n11092 0.019
R14934 GND.n11050 GND.n11048 0.019
R14935 GND.n11028 GND.n11027 0.019
R14936 GND.n13308 GND.n13305 0.019
R14937 GND.n13263 GND.n13261 0.019
R14938 GND.n13253 GND.n13252 0.019
R14939 GND.n11337 GND.n11335 0.019
R14940 GND.n11380 GND.n11379 0.019
R14941 GND.n11390 GND.n11388 0.019
R14942 GND.n13370 GND.n13362 0.019
R14943 GND.n13481 GND.n13479 0.019
R14944 GND.n12010 GND.n12008 0.019
R14945 GND.n11936 GND.n11935 0.019
R14946 GND.n11900 GND.n11898 0.019
R14947 GND.n11841 GND.n11832 0.019
R14948 GND.n12221 GND.n12212 0.019
R14949 GND.n12287 GND.n12285 0.019
R14950 GND.n12323 GND.n12322 0.019
R14951 GND.n12391 GND.n12389 0.019
R14952 GND.n13114 GND.n13112 0.019
R14953 GND.n13041 GND.n13040 0.019
R14954 GND.n13005 GND.n13003 0.019
R14955 GND.n12944 GND.n12936 0.019
R14956 GND.n7710 GND.n7702 0.019
R14957 GND.n7776 GND.n7774 0.019
R14958 GND.n7812 GND.n7811 0.019
R14959 GND.n7879 GND.n7877 0.019
R14960 GND.n8177 GND.n8175 0.019
R14961 GND.n8221 GND.n8220 0.019
R14962 GND.n6061 GND.n5831 0.019
R14963 GND.n8266 GND.n8264 0.019
R14964 GND.n8310 GND.n8309 0.019
R14965 GND.n8322 GND.n8320 0.019
R14966 GND.n6382 GND.n6380 0.019
R14967 GND.n6356 GND.n6354 0.019
R14968 GND.n5888 GND.n5885 0.019
R14969 GND.n5961 GND.n5959 0.019
R14970 GND.n5971 GND.n5969 0.019
R14971 GND.n6017 GND.n6014 0.019
R14972 GND.n6477 GND.n6475 0.019
R14973 GND.n6471 GND.n6470 0.019
R14974 GND.n6428 GND.n6426 0.019
R14975 GND.n8122 GND.n8120 0.019
R14976 GND.n8011 GND.n8003 0.019
R14977 GND.n7020 GND.n7012 0.019
R14978 GND.n7131 GND.n7129 0.019
R14979 GND.n6874 GND.n6872 0.019
R14980 GND.n6883 GND.n6881 0.019
R14981 GND.n6929 GND.n6926 0.019
R14982 GND.n6639 GND.n6637 0.019
R14983 GND.n6648 GND.n6646 0.019
R14984 GND.n6694 GND.n6691 0.019
R14985 GND.n6725 GND.n6723 0.019
R14986 GND.n6769 GND.n6768 0.019
R14987 GND.n6781 GND.n6779 0.019
R14988 GND.n7449 GND.n7447 0.019
R14989 GND.n7493 GND.n7492 0.019
R14990 GND.n6531 GND.n6163 0.019
R14991 GND.n7569 GND.n7566 0.019
R14992 GND.n7524 GND.n7522 0.019
R14993 GND.n7519 GND.n7518 0.019
R14994 GND.n7349 GND.n7347 0.019
R14995 GND.n7238 GND.n7229 0.019
R14996 GND.n15964 GND.n15955 0.019
R14997 GND.n16047 GND.n16045 0.019
R14998 GND.n16080 GND.n16079 0.019
R14999 GND.n16164 GND.n16162 0.019
R15000 GND.n1113 GND.n1111 0.019
R15001 GND.n1027 GND.n1023 0.019
R15002 GND.n991 GND.n989 0.019
R15003 GND.n911 GND.n903 0.019
R15004 GND.n9664 GND.n9655 0.019
R15005 GND.n9747 GND.n9745 0.019
R15006 GND.n9780 GND.n9779 0.019
R15007 GND.n9864 GND.n9862 0.019
R15008 GND.n1255 GND.n1247 0.019
R15009 GND.n1337 GND.n1335 0.019
R15010 GND.n1370 GND.n1369 0.019
R15011 GND.n1457 GND.n1455 0.019
R15012 GND.n10283 GND.n10281 0.019
R15013 GND.n10172 GND.n10163 0.019
R15014 GND.n8846 GND.n8844 0.019
R15015 GND.n8740 GND.n8732 0.019
R15016 GND.n8553 GND.n8551 0.019
R15017 GND.n8442 GND.n8433 0.019
R15018 GND.n9310 GND.n9308 0.019
R15019 GND.n9354 GND.n9353 0.019
R15020 GND.n9364 GND.n9362 0.019
R15021 GND.n1715 GND.n1713 0.019
R15022 GND.n1759 GND.n1758 0.019
R15023 GND.n1771 GND.n1769 0.019
R15024 GND.n1667 GND.n1665 0.019
R15025 GND.n9488 GND.n9486 0.019
R15026 GND.n9482 GND.n9481 0.019
R15027 GND.n9477 GND.n9476 0.019
R15028 GND.n9437 GND.n9435 0.019
R15029 GND.n1611 GND.n1610 0.019
R15030 GND.n1827 GND.n1825 0.019
R15031 GND.n1836 GND.n1834 0.019
R15032 GND.n1840 GND.n1839 0.019
R15033 GND.n1883 GND.n1880 0.019
R15034 GND.n8683 GND.n8680 0.019
R15035 GND.n8638 GND.n8636 0.019
R15036 GND.n8633 GND.n8632 0.019
R15037 GND.n10107 GND.n10105 0.019
R15038 GND.n10001 GND.n9993 0.019
R15039 GND.n8963 GND.n8954 0.019
R15040 GND.n9046 GND.n9044 0.019
R15041 GND.n9079 GND.n9078 0.019
R15042 GND.n9163 GND.n9161 0.019
R15043 GND.n4475 GND.n4473 0.019
R15044 GND.n4387 GND.n4383 0.019
R15045 GND.n4351 GND.n4349 0.019
R15046 GND.n4271 GND.n4263 0.019
R15047 GND.n2508 GND.n2506 0.019
R15048 GND.n2552 GND.n2551 0.019
R15049 GND.n2563 GND.n2561 0.019
R15050 GND.n3215 GND.n3207 0.019
R15051 GND.n3321 GND.n3319 0.019
R15052 GND.n2244 GND.n2243 0.019
R15053 GND.n3469 GND.n3467 0.019
R15054 GND.n3463 GND.n3462 0.019
R15055 GND.n3458 GND.n3457 0.019
R15056 GND.n3418 GND.n3416 0.019
R15057 GND.n2215 GND.n2214 0.019
R15058 GND.n2406 GND.n2404 0.019
R15059 GND.n2454 GND.n2453 0.019
R15060 GND.n2618 GND.n2615 0.019
R15061 GND.n2346 GND.n2344 0.019
R15062 GND.n2333 GND.n2331 0.019
R15063 GND.n2290 GND.n2289 0.019
R15064 GND.n5070 GND.n5068 0.019
R15065 GND.n4959 GND.n4951 0.019
R15066 GND.n5117 GND.n5115 0.019
R15067 GND.n5161 GND.n5160 0.019
R15068 GND.n5171 GND.n5169 0.019
R15069 GND.n2031 GND.n2030 0.019
R15070 GND.n2126 GND.n2124 0.019
R15071 GND.n2120 GND.n2119 0.019
R15072 GND.n2115 GND.n2114 0.019
R15073 GND.n2075 GND.n2073 0.019
R15074 GND.n1978 GND.n1977 0.019
R15075 GND.n2148 GND.n2146 0.019
R15076 GND.n2195 GND.n2194 0.019
R15077 GND.n2645 GND.n2642 0.019
R15078 GND.n2950 GND.n2947 0.019
R15079 GND.n2905 GND.n2903 0.019
R15080 GND.n2895 GND.n2894 0.019
R15081 GND.n4724 GND.n4722 0.019
R15082 GND.n4613 GND.n4605 0.019
R15083 GND.n3015 GND.n3007 0.019
R15084 GND.n3121 GND.n3119 0.019
R15085 GND.n10439 GND.n10431 0.019
R15086 GND.n10545 GND.n10543 0.019
R15087 GND.n15582 GND.n15574 0.019
R15088 GND.n15693 GND.n15691 0.019
R15089 GND.n15858 GND.n15855 0.019
R15090 GND.n15813 GND.n15811 0.019
R15091 GND.n15803 GND.n15802 0.019
R15092 GND.n15413 GND.n15410 0.019
R15093 GND.n15368 GND.n15366 0.019
R15094 GND.n15357 GND.n15356 0.019
R15095 GND.n14938 GND.n14936 0.019
R15096 GND.n14981 GND.n14980 0.019
R15097 GND.n14420 GND.n14413 0.019
R15098 GND.n15099 GND.n15096 0.019
R15099 GND.n15054 GND.n15052 0.019
R15100 GND.n15049 GND.n15048 0.019
R15101 GND.n15146 GND.n15138 0.019
R15102 GND.n15253 GND.n15251 0.019
R15103 GND.n3894 GND.n3892 0.019
R15104 GND.n3808 GND.n3804 0.019
R15105 GND.n3772 GND.n3770 0.019
R15106 GND.n3695 GND.n3687 0.019
R15107 GND.n5732 GND.n5730 0.019
R15108 GND.n5646 GND.n5642 0.019
R15109 GND.n5610 GND.n5608 0.019
R15110 GND.n5530 GND.n5522 0.019
R15111 GND.n16447 GND.n16446 0.019
R15112 GND.n16456 GND.n16454 0.019
R15113 GND.n16435 GND.n16434 0.019
R15114 GND.n16561 GND.n16560 0.019
R15115 GND.n16553 GND.n16552 0.019
R15116 GND.n16521 GND.n16520 0.019
R15117 GND.n16387 GND.n16386 0.019
R15118 GND.n16379 GND.n16377 0.019
R15119 GND.n16344 GND.n16343 0.019
R15120 GND.n16708 GND.n16707 0.019
R15121 GND.n16717 GND.n16715 0.019
R15122 GND.n16696 GND.n16695 0.019
R15123 GND.n16822 GND.n16821 0.019
R15124 GND.n16814 GND.n16813 0.019
R15125 GND.n16782 GND.n16781 0.019
R15126 GND.n16648 GND.n16647 0.019
R15127 GND.n16640 GND.n16638 0.019
R15128 GND.n16605 GND.n16604 0.019
R15129 GND.n16969 GND.n16968 0.019
R15130 GND.n16978 GND.n16976 0.019
R15131 GND.n16957 GND.n16956 0.019
R15132 GND.n17083 GND.n17082 0.019
R15133 GND.n17075 GND.n17074 0.019
R15134 GND.n17043 GND.n17042 0.019
R15135 GND.n16909 GND.n16908 0.019
R15136 GND.n16901 GND.n16899 0.019
R15137 GND.n16866 GND.n16865 0.019
R15138 GND.n17230 GND.n17229 0.019
R15139 GND.n17239 GND.n17237 0.019
R15140 GND.n17218 GND.n17217 0.019
R15141 GND.n17344 GND.n17343 0.019
R15142 GND.n17336 GND.n17335 0.019
R15143 GND.n17304 GND.n17303 0.019
R15144 GND.n17170 GND.n17169 0.019
R15145 GND.n17162 GND.n17160 0.019
R15146 GND.n17127 GND.n17126 0.019
R15147 GND.n17491 GND.n17490 0.019
R15148 GND.n17500 GND.n17498 0.019
R15149 GND.n17479 GND.n17478 0.019
R15150 GND.n17605 GND.n17604 0.019
R15151 GND.n17597 GND.n17596 0.019
R15152 GND.n17565 GND.n17564 0.019
R15153 GND.n17431 GND.n17430 0.019
R15154 GND.n17423 GND.n17421 0.019
R15155 GND.n17388 GND.n17387 0.019
R15156 GND.n674 GND.n673 0.019
R15157 GND.n666 GND.n665 0.019
R15158 GND.n777 GND.n776 0.019
R15159 GND.n769 GND.n768 0.019
R15160 GND.n608 GND.n607 0.019
R15161 GND.n600 GND.n599 0.019
R15162 GND.n416 GND.n415 0.019
R15163 GND.n408 GND.n407 0.019
R15164 GND.n519 GND.n518 0.019
R15165 GND.n511 GND.n510 0.019
R15166 GND.n350 GND.n349 0.019
R15167 GND.n342 GND.n341 0.019
R15168 GND.n158 GND.n157 0.019
R15169 GND.n150 GND.n149 0.019
R15170 GND.n261 GND.n260 0.019
R15171 GND.n253 GND.n252 0.019
R15172 GND.n92 GND.n91 0.019
R15173 GND.n84 GND.n83 0.019
R15174 GND.n17773 GND.n17772 0.019
R15175 GND.n17765 GND.n17764 0.019
R15176 GND.n17850 GND.n17849 0.019
R15177 GND.n17842 GND.n17841 0.019
R15178 GND.n17928 GND.n17927 0.019
R15179 GND.n17920 GND.n17919 0.019
R15180 GND.n9551 GND.n9549 0.019
R15181 GND.n12532 GND.n12527 0.019
R15182 GND.n13329 GND.n13328 0.019
R15183 GND.n14082 GND.n10400 0.019
R15184 GND.n14727 GND.n14722 0.019
R15185 GND.n4055 GND.n4054 0.018
R15186 GND.n4054 GND.n4053 0.018
R15187 GND.n4158 GND.n4157 0.018
R15188 GND.n3955 GND.n3954 0.018
R15189 GND.n17660 GND.n17659 0.018
R15190 GND.n732 GND.n731 0.018
R15191 GND.n701 GND.n685 0.018
R15192 GND.n474 GND.n473 0.018
R15193 GND.n443 GND.n427 0.018
R15194 GND.n216 GND.n215 0.018
R15195 GND.n185 GND.n169 0.018
R15196 GND.n17726 GND.n17725 0.018
R15197 GND.n17800 GND.n17784 0.018
R15198 GND.n14888 GND.n14886 0.017
R15199 GND.n14847 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SUBSTRATE
+ 0.017
R15200 GND.n14767 GND.n14765 0.017
R15201 GND.n6307 GND.n6305 0.017
R15202 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE GND.n6235
+ 0.017
R15203 GND.n6191 GND.n6189 0.017
R15204 GND.n12676 GND.n12674 0.017
R15205 GND.n12635 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE
+ 0.017
R15206 GND.n12555 GND.n12553 0.017
R15207 GND.n11288 GND.n11286 0.017
R15208 GND.n11172 GND.n11170 0.017
R15209 GND.n13695 GND.n13693 0.017
R15210 GND.n13579 GND.n13577 0.017
R15211 GND.n12832 GND.n12829 0.017
R15212 GND.n10890 GND.n10887 0.017
R15213 GND.n13362 GND.n13360 0.017
R15214 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE GND.n13408
+ 0.017
R15215 GND.n13483 GND.n13481 0.017
R15216 GND.n13333 GND.n13330 0.017
R15217 GND.n11123 GND.n11120 0.017
R15218 GND.n12012 GND.n12010 0.017
R15219 GND.n11970 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE
+ 0.017
R15220 GND.n11935 GND.n11933 0.017
R15221 GND.n11902 GND.n11900 0.017
R15222 GND.n11870 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.017
R15223 GND.n11832 GND.n11830 0.017
R15224 GND.n12212 GND.n12210 0.017
R15225 GND.n12289 GND.n12287 0.017
R15226 GND.n12322 GND.n12320 0.017
R15227 GND.n12393 GND.n12391 0.017
R15228 GND.n13116 GND.n13114 0.017
R15229 GND.n13040 GND.n13038 0.017
R15230 GND.n13007 GND.n13005 0.017
R15231 GND.n12936 GND.n12934 0.017
R15232 GND.n7702 GND.n7700 0.017
R15233 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE GND.n7751
+ 0.017
R15234 GND.n7778 GND.n7776 0.017
R15235 GND.n7811 GND.n7809 0.017
R15236 GND.n7840 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE
+ 0.017
R15237 GND.n7881 GND.n7879 0.017
R15238 GND.n8124 GND.n8122 0.017
R15239 GND.n8003 GND.n8001 0.017
R15240 GND.n7012 GND.n7010 0.017
R15241 GND.n7133 GND.n7131 0.017
R15242 GND.n7351 GND.n7349 0.017
R15243 GND.n7309 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE
+ 0.017
R15244 GND.n7229 GND.n7227 0.017
R15245 GND.n15955 GND.n15953 0.017
R15246 GND.n16049 GND.n16047 0.017
R15247 GND.n16079 GND.n16077 0.017
R15248 GND.n16166 GND.n16164 0.017
R15249 GND.n1115 GND.n1113 0.017
R15250 GND.n1075 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SUBSTRATE
+ 0.017
R15251 GND.n1023 GND.n1021 0.017
R15252 GND.n993 GND.n991 0.017
R15253 GND.n978 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SUBSTRATE
+ 0.017
R15254 GND.n903 GND.n901 0.017
R15255 GND.n9655 GND.n9653 0.017
R15256 GND.n9749 GND.n9747 0.017
R15257 GND.n9779 GND.n9777 0.017
R15258 GND.n9866 GND.n9864 0.017
R15259 GND.n1247 GND.n1245 0.017
R15260 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SUBSTRATE GND.n1296
+ 0.017
R15261 GND.n1339 GND.n1337 0.017
R15262 GND.n1369 GND.n1367 0.017
R15263 GND.n1381 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SUBSTRATE
+ 0.017
R15264 GND.n1459 GND.n1457 0.017
R15265 GND.n10285 GND.n10283 0.017
R15266 GND.n10163 GND.n10161 0.017
R15267 GND.n8848 GND.n8846 0.017
R15268 GND.n8808 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SUBSTRATE
+ 0.017
R15269 GND.n8732 GND.n8730 0.017
R15270 GND.n8555 GND.n8553 0.017
R15271 GND.n8513 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SUBSTRATE
+ 0.017
R15272 GND.n8433 GND.n8431 0.017
R15273 GND.n10109 GND.n10107 0.017
R15274 GND.n9993 GND.n9991 0.017
R15275 GND.n8954 GND.n8952 0.017
R15276 GND.n9048 GND.n9046 0.017
R15277 GND.n9078 GND.n9076 0.017
R15278 GND.n9165 GND.n9163 0.017
R15279 GND.n4477 GND.n4475 0.017
R15280 GND.n4383 GND.n4381 0.017
R15281 GND.n4353 GND.n4351 0.017
R15282 GND.n4263 GND.n4261 0.017
R15283 GND.n3207 GND.n3205 0.017
R15284 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SUBSTRATE GND.n3251
+ 0.017
R15285 GND.n3323 GND.n3321 0.017
R15286 GND.n5072 GND.n5070 0.017
R15287 GND.n4951 GND.n4949 0.017
R15288 GND.n4726 GND.n4724 0.017
R15289 GND.n4605 GND.n4603 0.017
R15290 GND.n3007 GND.n3005 0.017
R15291 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SUBSTRATE GND.n3051
+ 0.017
R15292 GND.n3123 GND.n3121 0.017
R15293 GND.n10431 GND.n10429 0.017
R15294 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SUBSTRATE GND.n10475
+ 0.017
R15295 GND.n10547 GND.n10545 0.017
R15296 GND.n15875 GND.n15872 0.017
R15297 GND.n14097 GND.n14094 0.017
R15298 GND.n15574 GND.n15572 0.017
R15299 GND.n15695 GND.n15693 0.017
R15300 GND.n14731 GND.n14728 0.017
R15301 GND.n14472 GND.n14379 0.017
R15302 GND.n15138 GND.n15136 0.017
R15303 GND.n15255 GND.n15253 0.017
R15304 GND.n3896 GND.n3894 0.017
R15305 GND.n3856 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SUBSTRATE
+ 0.017
R15306 GND.n3804 GND.n3802 0.017
R15307 GND.n3774 GND.n3772 0.017
R15308 GND.n3759 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SUBSTRATE
+ 0.017
R15309 GND.n3687 GND.n3685 0.017
R15310 GND.n5734 GND.n5732 0.017
R15311 GND.n5694 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SUBSTRATE
+ 0.017
R15312 GND.n5642 GND.n5640 0.017
R15313 GND.n5612 GND.n5610 0.017
R15314 GND.n5597 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SUBSTRATE
+ 0.017
R15315 GND.n5522 GND.n5520 0.017
R15316 GND.n16307 GND.n16306 0.017
R15317 GND.n14637 GND.n14636 0.016
R15318 GND.n14694 GND.n14692 0.016
R15319 GND.n14571 GND.n14570 0.016
R15320 GND.n14596 GND.n14594 0.016
R15321 GND.n10602 GND.n10600 0.016
R15322 GND.n15507 GND.n15505 0.016
R15323 GND.n14293 GND.n14292 0.016
R15324 GND.n14324 GND.n14322 0.016
R15325 GND.n14291 GND.n14290 0.016
R15326 GND.n14241 GND.n14239 0.016
R15327 GND.n3593 GND.n3591 0.016
R15328 GND.n4814 GND.n4812 0.016
R15329 GND.n10852 GND.n10850 0.016
R15330 GND.n13971 GND.n13969 0.016
R15331 GND.n13843 GND.n13841 0.016
R15332 GND.n13750 GND.n13748 0.016
R15333 GND.n12737 GND.n12735 0.016
R15334 GND.n11697 GND.n11695 0.016
R15335 GND.n11593 GND.n11591 0.016
R15336 GND.n11085 GND.n11083 0.016
R15337 GND.n13298 GND.n13296 0.016
R15338 GND.n11346 GND.n11344 0.016
R15339 GND.n8186 GND.n8184 0.016
R15340 GND.n8275 GND.n8273 0.016
R15341 GND.n5878 GND.n5876 0.016
R15342 GND.n6007 GND.n6005 0.016
R15343 GND.n6437 GND.n6435 0.016
R15344 GND.n6919 GND.n6917 0.016
R15345 GND.n6684 GND.n6682 0.016
R15346 GND.n6734 GND.n6732 0.016
R15347 GND.n7458 GND.n7456 0.016
R15348 GND.n7559 GND.n7557 0.016
R15349 GND.n9577 GND.n9576 0.016
R15350 GND.n9570 GND.n9567 0.016
R15351 GND.n9561 GND.n9557 0.016
R15352 GND.n1537 GND.n1535 0.016
R15353 GND.n1537 GND.n1536 0.016
R15354 GND.n1560 GND.n1559 0.016
R15355 GND.n16247 GND.n804 0.016
R15356 GND.n16260 GND.n16257 0.016
R15357 GND.n16300 GND.n16298 0.016
R15358 GND.n16269 GND.n16267 0.016
R15359 GND.n16269 GND.n16268 0.016
R15360 GND.n16287 GND.n16285 0.016
R15361 GND.n16287 GND.n16286 0.016
R15362 GND.n16274 GND.n16273 0.016
R15363 GND.n9319 GND.n9317 0.016
R15364 GND.n1724 GND.n1722 0.016
R15365 GND.n9496 GND.n9495 0.016
R15366 GND.n9446 GND.n9444 0.016
R15367 GND.n1816 GND.n1634 0.016
R15368 GND.n1873 GND.n1871 0.016
R15369 GND.n8673 GND.n8671 0.016
R15370 GND.n5308 GND.n5291 0.016
R15371 GND.n5319 GND.n5316 0.016
R15372 GND.n5334 GND.n5330 0.016
R15373 GND.n5258 GND.n5256 0.016
R15374 GND.n5258 GND.n5257 0.016
R15375 GND.n5285 GND.n5284 0.016
R15376 GND.n2517 GND.n2515 0.016
R15377 GND.n3477 GND.n3476 0.016
R15378 GND.n3427 GND.n3425 0.016
R15379 GND.n2394 GND.n2238 0.016
R15380 GND.n2423 GND.n2421 0.016
R15381 GND.n2355 GND.n2353 0.016
R15382 GND.n5126 GND.n5124 0.016
R15383 GND.n2134 GND.n2133 0.016
R15384 GND.n2084 GND.n2082 0.016
R15385 GND.n2136 GND.n2135 0.016
R15386 GND.n2164 GND.n2162 0.016
R15387 GND.n2940 GND.n2938 0.016
R15388 GND.n15848 GND.n15846 0.016
R15389 GND.n15403 GND.n15401 0.016
R15390 GND.n14947 GND.n14945 0.016
R15391 GND.n15089 GND.n15087 0.016
R15392 GND.n5424 GND.n5250 0.016
R15393 GND.n5382 GND.n5381 0.016
R15394 GND.n5397 GND.n5395 0.016
R15395 GND.n5397 GND.n5396 0.016
R15396 GND.n5405 GND.n5404 0.016
R15397 GND.n5405 GND.n5403 0.016
R15398 GND.n5417 GND.n5416 0.016
R15399 GND.n5417 GND.n5415 0.016
R15400 GND.n5370 GND.n5369 0.016
R15401 GND.n16335 GND.n16334 0.016
R15402 GND.n16596 GND.n16595 0.016
R15403 GND.n16857 GND.n16856 0.016
R15404 GND.n17118 GND.n17117 0.016
R15405 GND.n17379 GND.n17378 0.016
R15406 GND.n16511 GND.n16510 0.016
R15407 GND.n16772 GND.n16771 0.016
R15408 GND.n17033 GND.n17032 0.016
R15409 GND.n17294 GND.n17293 0.016
R15410 GND.n17555 GND.n17554 0.016
R15411 GND.n558 GND.n557 0.015
R15412 GND.n300 GND.n299 0.015
R15413 GND.n42 GND.n41 0.015
R15414 GND.n17878 GND.n17877 0.015
R15415 GND.n14874 GND.n14872 0.015
R15416 GND.n14788 GND.n14779 0.015
R15417 GND.n6293 GND.n6291 0.015
R15418 GND.n6211 GND.n6203 0.015
R15419 GND.n12662 GND.n12660 0.015
R15420 GND.n12576 GND.n12567 0.015
R15421 GND.n11274 GND.n11272 0.015
R15422 GND.n11192 GND.n11184 0.015
R15423 GND.n13681 GND.n13679 0.015
R15424 GND.n13599 GND.n13591 0.015
R15425 GND.n13383 GND.n13374 0.015
R15426 GND.n13469 GND.n13467 0.015
R15427 GND.n11997 GND.n11995 0.015
R15428 GND.n11941 GND.n11940 0.015
R15429 GND.n11895 GND.n11894 0.015
R15430 GND.n11853 GND.n11845 0.015
R15431 GND.n12233 GND.n12225 0.015
R15432 GND.n12282 GND.n12280 0.015
R15433 GND.n12327 GND.n12326 0.015
R15434 GND.n12379 GND.n12377 0.015
R15435 GND.n13102 GND.n13100 0.015
R15436 GND.n13046 GND.n13045 0.015
R15437 GND.n13000 GND.n12999 0.015
R15438 GND.n12957 GND.n12948 0.015
R15439 GND.n7722 GND.n7714 0.015
R15440 GND.n7771 GND.n7769 0.015
R15441 GND.n7816 GND.n7815 0.015
R15442 GND.n7866 GND.n7864 0.015
R15443 GND.n8110 GND.n8108 0.015
R15444 GND.n8024 GND.n8015 0.015
R15445 GND.n7033 GND.n7024 0.015
R15446 GND.n7119 GND.n7117 0.015
R15447 GND.n7336 GND.n7334 0.015
R15448 GND.n7250 GND.n7242 0.015
R15449 GND.n15976 GND.n15968 0.015
R15450 GND.n16039 GND.n16037 0.015
R15451 GND.n16084 GND.n16083 0.015
R15452 GND.n16152 GND.n16150 0.015
R15453 GND.n1101 GND.n1099 0.015
R15454 GND.n1035 GND.n1031 0.015
R15455 GND.n986 GND.n985 0.015
R15456 GND.n924 GND.n915 0.015
R15457 GND.n9676 GND.n9668 0.015
R15458 GND.n9739 GND.n9737 0.015
R15459 GND.n9784 GND.n9783 0.015
R15460 GND.n9852 GND.n9850 0.015
R15461 GND.n1267 GND.n1259 0.015
R15462 GND.n1329 GND.n1327 0.015
R15463 GND.n1374 GND.n1373 0.015
R15464 GND.n1445 GND.n1443 0.015
R15465 GND.n10270 GND.n10268 0.015
R15466 GND.n10184 GND.n10176 0.015
R15467 GND.n8834 GND.n8832 0.015
R15468 GND.n8752 GND.n8744 0.015
R15469 GND.n8540 GND.n8538 0.015
R15470 GND.n8454 GND.n8446 0.015
R15471 GND.n10095 GND.n10093 0.015
R15472 GND.n10013 GND.n10005 0.015
R15473 GND.n9241 GND.n9240 0.015
R15474 GND.n8975 GND.n8967 0.015
R15475 GND.n9038 GND.n9036 0.015
R15476 GND.n9083 GND.n9082 0.015
R15477 GND.n9151 GND.n9149 0.015
R15478 GND.n4462 GND.n4460 0.015
R15479 GND.n4395 GND.n4391 0.015
R15480 GND.n4346 GND.n4345 0.015
R15481 GND.n4284 GND.n4275 0.015
R15482 GND.n3227 GND.n3219 0.015
R15483 GND.n3309 GND.n3307 0.015
R15484 GND.n5058 GND.n5056 0.015
R15485 GND.n4972 GND.n4963 0.015
R15486 GND.n3400 GND.n3398 0.015
R15487 GND.n4771 GND.n4769 0.015
R15488 GND.n4712 GND.n4710 0.015
R15489 GND.n4626 GND.n4617 0.015
R15490 GND.n3027 GND.n3019 0.015
R15491 GND.n3109 GND.n3107 0.015
R15492 GND.n10451 GND.n10443 0.015
R15493 GND.n10533 GND.n10531 0.015
R15494 GND.n15595 GND.n15586 0.015
R15495 GND.n15681 GND.n15679 0.015
R15496 GND.n15158 GND.n15150 0.015
R15497 GND.n15240 GND.n15238 0.015
R15498 GND.n3882 GND.n3880 0.015
R15499 GND.n3816 GND.n3812 0.015
R15500 GND.n3767 GND.n3766 0.015
R15501 GND.n3707 GND.n3699 0.015
R15502 GND.n4544 GND.n4543 0.015
R15503 GND.n5720 GND.n5718 0.015
R15504 GND.n5654 GND.n5650 0.015
R15505 GND.n5605 GND.n5604 0.015
R15506 GND.n5543 GND.n5534 0.015
R15507 GND.n5437 GND.n5432 0.015
R15508 GND.n9526 GND.n9525 0.014
R15509 GND.n14521 GND.n14518 0.014
R15510 GND.n14517 GND.n14515 0.014
R15511 GND.n14659 GND.n14657 0.014
R15512 GND.n14711 GND.n14708 0.014
R15513 GND.n14554 GND.n14552 0.014
R15514 GND.n14558 GND.n14556 0.014
R15515 GND.n14628 GND.n14591 0.014
R15516 GND.n14396 GND.n14393 0.014
R15517 GND.n10586 GND.n10584 0.014
R15518 GND.n10636 GND.n10634 0.014
R15519 GND.n10671 GND.n10669 0.014
R15520 GND.n10676 GND.n10673 0.014
R15521 GND.n15524 GND.n15521 0.014
R15522 GND.n15473 GND.n15472 0.014
R15523 GND.n14056 GND.n14054 0.014
R15524 GND.n14052 GND.n14051 0.014
R15525 GND.n14143 GND.n14141 0.014
R15526 GND.n14147 GND.n14145 0.014
R15527 GND.n14357 GND.n14317 0.014
R15528 GND.n10708 GND.n10705 0.014
R15529 GND.n14196 GND.n14194 0.014
R15530 GND.n14200 GND.n14198 0.014
R15531 GND.n14276 GND.n14274 0.014
R15532 GND.n14225 GND.n14223 0.014
R15533 GND.n3610 GND.n3607 0.014
R15534 GND.n3559 GND.n3558 0.014
R15535 GND.n3528 GND.n3526 0.014
R15536 GND.n3524 GND.n3522 0.014
R15537 GND.n4798 GND.n4796 0.014
R15538 GND.n4848 GND.n4846 0.014
R15539 GND.n4882 GND.n4880 0.014
R15540 GND.n4887 GND.n4884 0.014
R15541 GND.n10805 GND.n10803 0.014
R15542 GND.n10809 GND.n10807 0.014
R15543 GND.n10767 GND.n10765 0.014
R15544 GND.n10869 GND.n10866 0.014
R15545 GND.n13904 GND.n13902 0.014
R15546 GND.n13908 GND.n13906 0.014
R15547 GND.n13937 GND.n13935 0.014
R15548 GND.n13988 GND.n13985 0.014
R15549 GND.n13860 GND.n13857 0.014
R15550 GND.n13809 GND.n13808 0.014
R15551 GND.n10928 GND.n10926 0.014
R15552 GND.n10924 GND.n10923 0.014
R15553 GND.n13734 GND.n13732 0.014
R15554 GND.n13783 GND.n13781 0.014
R15555 GND.n10977 GND.n10975 0.014
R15556 GND.n10973 GND.n10972 0.014
R15557 GND.n12721 GND.n12719 0.014
R15558 GND.n12771 GND.n12769 0.014
R15559 GND.n12805 GND.n12803 0.014
R15560 GND.n12810 GND.n12807 0.014
R15561 GND.n11466 GND.n11464 0.014
R15562 GND.n11470 GND.n11468 0.014
R15563 GND.n11663 GND.n11661 0.014
R15564 GND.n11714 GND.n11711 0.014
R15565 GND.n11526 GND.n11524 0.014
R15566 GND.n11530 GND.n11528 0.014
R15567 GND.n11559 GND.n11557 0.014
R15568 GND.n11610 GND.n11607 0.014
R15569 GND.n11102 GND.n11099 0.014
R15570 GND.n11051 GND.n11050 0.014
R15571 GND.n11630 GND.n11628 0.014
R15572 GND.n11635 GND.n11632 0.014
R15573 GND.n13315 GND.n13312 0.014
R15574 GND.n13264 GND.n13263 0.014
R15575 GND.n13232 GND.n13230 0.014
R15576 GND.n13228 GND.n13227 0.014
R15577 GND.n11330 GND.n11328 0.014
R15578 GND.n11379 GND.n11377 0.014
R15579 GND.n11412 GND.n11410 0.014
R15580 GND.n11417 GND.n11414 0.014
R15581 GND.n8170 GND.n8168 0.014
R15582 GND.n8220 GND.n8218 0.014
R15583 GND.n6083 GND.n6081 0.014
R15584 GND.n6088 GND.n6085 0.014
R15585 GND.n8259 GND.n8257 0.014
R15586 GND.n8309 GND.n8307 0.014
R15587 GND.n8344 GND.n8342 0.014
R15588 GND.n8349 GND.n8346 0.014
R15589 GND.n6398 GND.n6395 0.014
R15590 GND.n6394 GND.n6392 0.014
R15591 GND.n6358 GND.n6356 0.014
R15592 GND.n5895 GND.n5892 0.014
R15593 GND.n5935 GND.n5933 0.014
R15594 GND.n5939 GND.n5937 0.014
R15595 GND.n5973 GND.n5971 0.014
R15596 GND.n6024 GND.n6021 0.014
R15597 GND.n6501 GND.n6498 0.014
R15598 GND.n6497 GND.n6495 0.014
R15599 GND.n6470 GND.n6468 0.014
R15600 GND.n6421 GND.n6419 0.014
R15601 GND.n6848 GND.n6846 0.014
R15602 GND.n6852 GND.n6850 0.014
R15603 GND.n6885 GND.n6883 0.014
R15604 GND.n6936 GND.n6933 0.014
R15605 GND.n6613 GND.n6611 0.014
R15606 GND.n6617 GND.n6615 0.014
R15607 GND.n6650 GND.n6648 0.014
R15608 GND.n6701 GND.n6698 0.014
R15609 GND.n6718 GND.n6716 0.014
R15610 GND.n6768 GND.n6766 0.014
R15611 GND.n6803 GND.n6801 0.014
R15612 GND.n6808 GND.n6805 0.014
R15613 GND.n7442 GND.n7440 0.014
R15614 GND.n7492 GND.n7490 0.014
R15615 GND.n6553 GND.n6551 0.014
R15616 GND.n6558 GND.n6555 0.014
R15617 GND.n7576 GND.n7573 0.014
R15618 GND.n7525 GND.n7524 0.014
R15619 GND.n6962 GND.n6960 0.014
R15620 GND.n6967 GND.n6964 0.014
R15621 GND.n9303 GND.n9301 0.014
R15622 GND.n9353 GND.n9351 0.014
R15623 GND.n9386 GND.n9384 0.014
R15624 GND.n9391 GND.n9388 0.014
R15625 GND.n1708 GND.n1706 0.014
R15626 GND.n1758 GND.n1756 0.014
R15627 GND.n1793 GND.n1791 0.014
R15628 GND.n1798 GND.n1795 0.014
R15629 GND.n1662 GND.n1659 0.014
R15630 GND.n1658 GND.n1656 0.014
R15631 GND.n9481 GND.n9479 0.014
R15632 GND.n9430 GND.n9428 0.014
R15633 GND.n1618 GND.n1616 0.014
R15634 GND.n1622 GND.n1620 0.014
R15635 GND.n1838 GND.n1836 0.014
R15636 GND.n1890 GND.n1887 0.014
R15637 GND.n8690 GND.n8687 0.014
R15638 GND.n8639 GND.n8638 0.014
R15639 GND.n8612 GND.n8610 0.014
R15640 GND.n8608 GND.n8606 0.014
R15641 GND.n2501 GND.n2499 0.014
R15642 GND.n2551 GND.n2549 0.014
R15643 GND.n2585 GND.n2583 0.014
R15644 GND.n2590 GND.n2587 0.014
R15645 GND.n2251 GND.n2249 0.014
R15646 GND.n2255 GND.n2253 0.014
R15647 GND.n3462 GND.n3460 0.014
R15648 GND.n3411 GND.n3409 0.014
R15649 GND.n2222 GND.n2220 0.014
R15650 GND.n2226 GND.n2224 0.014
R15651 GND.n2456 GND.n2419 0.014
R15652 GND.n2625 GND.n2622 0.014
R15653 GND.n2339 GND.n2337 0.014
R15654 GND.n2334 GND.n2333 0.014
R15655 GND.n2323 GND.n2321 0.014
R15656 GND.n2328 GND.n2325 0.014
R15657 GND.n5110 GND.n5108 0.014
R15658 GND.n5160 GND.n5158 0.014
R15659 GND.n5193 GND.n5191 0.014
R15660 GND.n5198 GND.n5195 0.014
R15661 GND.n2038 GND.n2036 0.014
R15662 GND.n2042 GND.n2040 0.014
R15663 GND.n2119 GND.n2117 0.014
R15664 GND.n2068 GND.n2066 0.014
R15665 GND.n1985 GND.n1983 0.014
R15666 GND.n1989 GND.n1987 0.014
R15667 GND.n2197 GND.n2160 0.014
R15668 GND.n2652 GND.n2649 0.014
R15669 GND.n2957 GND.n2954 0.014
R15670 GND.n2906 GND.n2905 0.014
R15671 GND.n2874 GND.n2872 0.014
R15672 GND.n2870 GND.n2868 0.014
R15673 GND.n15865 GND.n15862 0.014
R15674 GND.n15814 GND.n15813 0.014
R15675 GND.n15782 GND.n15780 0.014
R15676 GND.n15778 GND.n15777 0.014
R15677 GND.n15420 GND.n15417 0.014
R15678 GND.n15369 GND.n15368 0.014
R15679 GND.n15336 GND.n15334 0.014
R15680 GND.n15332 GND.n15331 0.014
R15681 GND.n14931 GND.n14929 0.014
R15682 GND.n14980 GND.n14978 0.014
R15683 GND.n14442 GND.n14440 0.014
R15684 GND.n14447 GND.n14444 0.014
R15685 GND.n15106 GND.n15103 0.014
R15686 GND.n15055 GND.n15054 0.014
R15687 GND.n15028 GND.n15026 0.014
R15688 GND.n15024 GND.n15023 0.014
R15689 GND.n16446 GND.n16444 0.014
R15690 GND.n16481 GND.n16479 0.014
R15691 GND.n16430 GND.n16429 0.014
R15692 GND.n16560 GND.n16558 0.014
R15693 GND.n16516 GND.n16514 0.014
R15694 GND.n16500 GND.n16497 0.014
R15695 GND.n16386 GND.n16384 0.014
R15696 GND.n16355 GND.n16353 0.014
R15697 GND.n16339 GND.n16338 0.014
R15698 GND.n16707 GND.n16705 0.014
R15699 GND.n16742 GND.n16740 0.014
R15700 GND.n16691 GND.n16690 0.014
R15701 GND.n16821 GND.n16819 0.014
R15702 GND.n16777 GND.n16775 0.014
R15703 GND.n16761 GND.n16758 0.014
R15704 GND.n16647 GND.n16645 0.014
R15705 GND.n16616 GND.n16614 0.014
R15706 GND.n16600 GND.n16599 0.014
R15707 GND.n16968 GND.n16966 0.014
R15708 GND.n17003 GND.n17001 0.014
R15709 GND.n16952 GND.n16951 0.014
R15710 GND.n17082 GND.n17080 0.014
R15711 GND.n17038 GND.n17036 0.014
R15712 GND.n17022 GND.n17019 0.014
R15713 GND.n16908 GND.n16906 0.014
R15714 GND.n16877 GND.n16875 0.014
R15715 GND.n16861 GND.n16860 0.014
R15716 GND.n17229 GND.n17227 0.014
R15717 GND.n17264 GND.n17262 0.014
R15718 GND.n17213 GND.n17212 0.014
R15719 GND.n17343 GND.n17341 0.014
R15720 GND.n17299 GND.n17297 0.014
R15721 GND.n17283 GND.n17280 0.014
R15722 GND.n17169 GND.n17167 0.014
R15723 GND.n17138 GND.n17136 0.014
R15724 GND.n17122 GND.n17121 0.014
R15725 GND.n17490 GND.n17488 0.014
R15726 GND.n17525 GND.n17523 0.014
R15727 GND.n17474 GND.n17473 0.014
R15728 GND.n17604 GND.n17602 0.014
R15729 GND.n17560 GND.n17558 0.014
R15730 GND.n17544 GND.n17541 0.014
R15731 GND.n17430 GND.n17428 0.014
R15732 GND.n17399 GND.n17397 0.014
R15733 GND.n17383 GND.n17382 0.014
R15734 GND.n673 GND.n671 0.014
R15735 GND.n694 GND.n691 0.014
R15736 GND.n776 GND.n774 0.014
R15737 GND.n721 GND.n718 0.014
R15738 GND.n607 GND.n605 0.014
R15739 GND.n562 GND.n561 0.014
R15740 GND.n415 GND.n413 0.014
R15741 GND.n436 GND.n433 0.014
R15742 GND.n518 GND.n516 0.014
R15743 GND.n463 GND.n460 0.014
R15744 GND.n349 GND.n347 0.014
R15745 GND.n304 GND.n303 0.014
R15746 GND.n157 GND.n155 0.014
R15747 GND.n178 GND.n175 0.014
R15748 GND.n260 GND.n258 0.014
R15749 GND.n205 GND.n202 0.014
R15750 GND.n91 GND.n89 0.014
R15751 GND.n46 GND.n45 0.014
R15752 GND.n17772 GND.n17770 0.014
R15753 GND.n17793 GND.n17790 0.014
R15754 GND.n17849 GND.n17847 0.014
R15755 GND.n17715 GND.n17712 0.014
R15756 GND.n17927 GND.n17925 0.014
R15757 GND.n17882 GND.n17881 0.014
R15758 GND.n3356 GND.n3355 0.013
R15759 GND.n2972 GND.n2969 0.013
R15760 GND.n17669 GND.n17668 0.013
R15761 GND.n17668 GND.n17667 0.013
R15762 GND.n9544 GND.n9533 0.013
R15763 GND.n718 GND.n716 0.012
R15764 GND.n553 GND.n552 0.012
R15765 GND.n716 GND.n715 0.012
R15766 GND.n552 GND.n551 0.012
R15767 GND.n460 GND.n458 0.012
R15768 GND.n295 GND.n294 0.012
R15769 GND.n458 GND.n457 0.012
R15770 GND.n294 GND.n293 0.012
R15771 GND.n202 GND.n200 0.012
R15772 GND.n37 GND.n36 0.012
R15773 GND.n200 GND.n199 0.012
R15774 GND.n36 GND.n35 0.012
R15775 GND.n17712 GND.n17710 0.012
R15776 GND.n17873 GND.n17872 0.012
R15777 GND.n17710 GND.n17709 0.012
R15778 GND.n17872 GND.n17871 0.012
R15779 GND.n14185 GND.n14173 0.012
R15780 GND.n1672 GND.n1669 0.012
R15781 GND.n2465 GND.n2205 0.012
R15782 GND.n2027 GND.n2015 0.012
R15783 GND.n14528 GND.n14502 0.012
R15784 GND.n14522 GND.n14521 0.012
R15785 GND.n14687 GND.n14685 0.012
R15786 GND.n14552 GND.n14549 0.012
R15787 GND.n14603 GND.n14601 0.012
R15788 GND.n10609 GND.n10607 0.012
R15789 GND.n15500 GND.n15498 0.012
R15790 GND.n14141 GND.n14138 0.012
R15791 GND.n14331 GND.n14329 0.012
R15792 GND.n14194 GND.n14191 0.012
R15793 GND.n14248 GND.n14246 0.012
R15794 GND.n14901 GND.n14899 0.012
R15795 GND.n14754 GND.n14752 0.012
R15796 GND.n3586 GND.n3584 0.012
R15797 GND.n4821 GND.n4819 0.012
R15798 GND.n6319 GND.n6317 0.012
R15799 GND.n6178 GND.n6176 0.012
R15800 GND.n12689 GND.n12687 0.012
R15801 GND.n12542 GND.n12540 0.012
R15802 GND.n10741 GND.n10739 0.012
R15803 GND.n13964 GND.n13962 0.012
R15804 GND.n13836 GND.n13834 0.012
R15805 GND.n13757 GND.n13755 0.012
R15806 GND.n11300 GND.n11298 0.012
R15807 GND.n11160 GND.n11158 0.012
R15808 GND.n13707 GND.n13705 0.012
R15809 GND.n13567 GND.n13565 0.012
R15810 GND.n12744 GND.n12742 0.012
R15811 GND.n11690 GND.n11688 0.012
R15812 GND.n11586 GND.n11584 0.012
R15813 GND.n11078 GND.n11076 0.012
R15814 GND.n13291 GND.n13289 0.012
R15815 GND.n11353 GND.n11351 0.012
R15816 GND.n13349 GND.n13347 0.012
R15817 GND.n13496 GND.n13494 0.012
R15818 GND.n12024 GND.n12022 0.012
R15819 GND.n11930 GND.n11928 0.012
R15820 GND.n11907 GND.n11905 0.012
R15821 GND.n11820 GND.n11818 0.012
R15822 GND.n12200 GND.n12198 0.012
R15823 GND.n12294 GND.n12292 0.012
R15824 GND.n12317 GND.n12315 0.012
R15825 GND.n12406 GND.n12404 0.012
R15826 GND.n13128 GND.n13126 0.012
R15827 GND.n13035 GND.n13033 0.012
R15828 GND.n13012 GND.n13010 0.012
R15829 GND.n12923 GND.n12921 0.012
R15830 GND.n7690 GND.n7688 0.012
R15831 GND.n7783 GND.n7781 0.012
R15832 GND.n7806 GND.n7804 0.012
R15833 GND.n7893 GND.n7891 0.012
R15834 GND.n8193 GND.n8191 0.012
R15835 GND.n8282 GND.n8280 0.012
R15836 GND.n5871 GND.n5869 0.012
R15837 GND.n6000 GND.n5998 0.012
R15838 GND.n6444 GND.n6442 0.012
R15839 GND.n8137 GND.n8135 0.012
R15840 GND.n7990 GND.n7988 0.012
R15841 GND.n6999 GND.n6997 0.012
R15842 GND.n7146 GND.n7144 0.012
R15843 GND.n6912 GND.n6910 0.012
R15844 GND.n6677 GND.n6675 0.012
R15845 GND.n6741 GND.n6739 0.012
R15846 GND.n7465 GND.n7463 0.012
R15847 GND.n7552 GND.n7550 0.012
R15848 GND.n7363 GND.n7361 0.012
R15849 GND.n7217 GND.n7215 0.012
R15850 GND.n15943 GND.n15941 0.012
R15851 GND.n16057 GND.n16055 0.012
R15852 GND.n16074 GND.n16072 0.012
R15853 GND.n16179 GND.n16177 0.012
R15854 GND.n1127 GND.n1125 0.012
R15855 GND.n1015 GND.n1013 0.012
R15856 GND.n998 GND.n996 0.012
R15857 GND.n890 GND.n888 0.012
R15858 GND.n9643 GND.n9641 0.012
R15859 GND.n9757 GND.n9755 0.012
R15860 GND.n9774 GND.n9772 0.012
R15861 GND.n9879 GND.n9877 0.012
R15862 GND.n1235 GND.n1233 0.012
R15863 GND.n1347 GND.n1345 0.012
R15864 GND.n1364 GND.n1362 0.012
R15865 GND.n1472 GND.n1470 0.012
R15866 GND.n10297 GND.n10295 0.012
R15867 GND.n10151 GND.n10149 0.012
R15868 GND.n8860 GND.n8858 0.012
R15869 GND.n8720 GND.n8718 0.012
R15870 GND.n8567 GND.n8565 0.012
R15871 GND.n8421 GND.n8419 0.012
R15872 GND.n9326 GND.n9324 0.012
R15873 GND.n1731 GND.n1729 0.012
R15874 GND.n1663 GND.n1662 0.012
R15875 GND.n9453 GND.n9451 0.012
R15876 GND.n1616 GND.n1613 0.012
R15877 GND.n1866 GND.n1864 0.012
R15878 GND.n8666 GND.n8664 0.012
R15879 GND.n10121 GND.n10119 0.012
R15880 GND.n9980 GND.n9978 0.012
R15881 GND.n8942 GND.n8940 0.012
R15882 GND.n9056 GND.n9054 0.012
R15883 GND.n9073 GND.n9071 0.012
R15884 GND.n9178 GND.n9176 0.012
R15885 GND.n4489 GND.n4487 0.012
R15886 GND.n4375 GND.n4373 0.012
R15887 GND.n4358 GND.n4356 0.012
R15888 GND.n4250 GND.n4248 0.012
R15889 GND.n2524 GND.n2522 0.012
R15890 GND.n3195 GND.n3193 0.012
R15891 GND.n3336 GND.n3334 0.012
R15892 GND.n2249 GND.n2246 0.012
R15893 GND.n3434 GND.n3432 0.012
R15894 GND.n2220 GND.n2217 0.012
R15895 GND.n2430 GND.n2428 0.012
R15896 GND.n2362 GND.n2360 0.012
R15897 GND.n5085 GND.n5083 0.012
R15898 GND.n4938 GND.n4936 0.012
R15899 GND.n5133 GND.n5131 0.012
R15900 GND.n2036 GND.n2033 0.012
R15901 GND.n2091 GND.n2089 0.012
R15902 GND.n1983 GND.n1980 0.012
R15903 GND.n2171 GND.n2169 0.012
R15904 GND.n2933 GND.n2931 0.012
R15905 GND.n2979 GND.n2978 0.012
R15906 GND.n4739 GND.n4737 0.012
R15907 GND.n4592 GND.n4590 0.012
R15908 GND.n2995 GND.n2993 0.012
R15909 GND.n3136 GND.n3134 0.012
R15910 GND.n10419 GND.n10417 0.012
R15911 GND.n10559 GND.n10557 0.012
R15912 GND.n15561 GND.n15559 0.012
R15913 GND.n15708 GND.n15706 0.012
R15914 GND.n15841 GND.n15839 0.012
R15915 GND.n15396 GND.n15394 0.012
R15916 GND.n14954 GND.n14952 0.012
R15917 GND.n15082 GND.n15080 0.012
R15918 GND.n15126 GND.n15124 0.012
R15919 GND.n15267 GND.n15265 0.012
R15920 GND.n3908 GND.n3906 0.012
R15921 GND.n3796 GND.n3794 0.012
R15922 GND.n3779 GND.n3777 0.012
R15923 GND.n3674 GND.n3672 0.012
R15924 GND.n5746 GND.n5744 0.012
R15925 GND.n5634 GND.n5632 0.012
R15926 GND.n5617 GND.n5615 0.012
R15927 GND.n5509 GND.n5507 0.012
R15928 GND.n643 GND.n641 0.012
R15929 GND.n745 GND.n743 0.012
R15930 GND.n577 GND.n575 0.012
R15931 GND.n385 GND.n383 0.012
R15932 GND.n487 GND.n485 0.012
R15933 GND.n319 GND.n317 0.012
R15934 GND.n127 GND.n125 0.012
R15935 GND.n229 GND.n227 0.012
R15936 GND.n61 GND.n59 0.012
R15937 GND.n17742 GND.n17740 0.012
R15938 GND.n17818 GND.n17816 0.012
R15939 GND.n17897 GND.n17895 0.012
R15940 GND.n5265 GND.n5264 0.012
R15941 GND.n14542 GND.n14541 0.011
R15942 GND.n14132 GND.n14131 0.011
R15943 GND.n1606 GND.n1594 0.011
R15944 GND.n2210 GND.n2209 0.011
R15945 GND.n1973 GND.n1972 0.011
R15946 GND.n8382 GND.n8381 0.011
R15947 GND.n7431 GND.n7430 0.011
R15948 GND.n9246 GND.n9245 0.011
R15949 GND.n10330 GND.n10325 0.011
R15950 GND.n637 GND.n636 0.011
R15951 GND.n739 GND.n738 0.011
R15952 GND.n571 GND.n570 0.011
R15953 GND.n379 GND.n378 0.011
R15954 GND.n481 GND.n480 0.011
R15955 GND.n313 GND.n312 0.011
R15956 GND.n121 GND.n120 0.011
R15957 GND.n223 GND.n222 0.011
R15958 GND.n55 GND.n54 0.011
R15959 GND.n17736 GND.n17735 0.011
R15960 GND.n17812 GND.n17811 0.011
R15961 GND.n17891 GND.n17890 0.011
R15962 GND.n16432 GND.n16431 0.011
R15963 GND.n16420 GND.n16419 0.011
R15964 GND.n16497 GND.n16495 0.011
R15965 GND.n16340 GND.n16339 0.011
R15966 GND.n16421 GND.n16420 0.011
R15967 GND.n16341 GND.n16340 0.011
R15968 GND.n16431 GND.n16430 0.011
R15969 GND.n16693 GND.n16692 0.011
R15970 GND.n16681 GND.n16680 0.011
R15971 GND.n16758 GND.n16756 0.011
R15972 GND.n16601 GND.n16600 0.011
R15973 GND.n16682 GND.n16681 0.011
R15974 GND.n16602 GND.n16601 0.011
R15975 GND.n16692 GND.n16691 0.011
R15976 GND.n16954 GND.n16953 0.011
R15977 GND.n16942 GND.n16941 0.011
R15978 GND.n17019 GND.n17017 0.011
R15979 GND.n16862 GND.n16861 0.011
R15980 GND.n16943 GND.n16942 0.011
R15981 GND.n16863 GND.n16862 0.011
R15982 GND.n16953 GND.n16952 0.011
R15983 GND.n17215 GND.n17214 0.011
R15984 GND.n17203 GND.n17202 0.011
R15985 GND.n17280 GND.n17278 0.011
R15986 GND.n17123 GND.n17122 0.011
R15987 GND.n17204 GND.n17203 0.011
R15988 GND.n17124 GND.n17123 0.011
R15989 GND.n17214 GND.n17213 0.011
R15990 GND.n17476 GND.n17475 0.011
R15991 GND.n17464 GND.n17463 0.011
R15992 GND.n17541 GND.n17539 0.011
R15993 GND.n17384 GND.n17383 0.011
R15994 GND.n17465 GND.n17464 0.011
R15995 GND.n17385 GND.n17384 0.011
R15996 GND.n17475 GND.n17474 0.011
R15997 GND.n9531 GND.n1567 0.01
R15998 GND.n9540 GND.n9539 0.01
R15999 GND.n14861 GND.n14859 0.01
R16000 GND.n14800 GND.n14792 0.01
R16001 GND.n6281 GND.n6279 0.01
R16002 GND.n6223 GND.n6215 0.01
R16003 GND.n12649 GND.n12647 0.01
R16004 GND.n12588 GND.n12580 0.01
R16005 GND.n11262 GND.n11260 0.01
R16006 GND.n11204 GND.n11196 0.01
R16007 GND.n13669 GND.n13667 0.01
R16008 GND.n13611 GND.n13603 0.01
R16009 GND.n12836 GND.n12835 0.01
R16010 GND.n10879 GND.n10877 0.01
R16011 GND.n10901 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE 0.01
R16012 GND.n13996 GND.n10724 0.01
R16013 GND.n13999 GND.n13996 0.01
R16014 GND.n13395 GND.n13387 0.01
R16015 GND.n13456 GND.n13454 0.01
R16016 GND.n13337 GND.n13336 0.01
R16017 GND.n11112 GND.n11110 0.01
R16018 GND.n11141 GND.n11139 0.01
R16019 GND.n11144 GND.n11141 0.01
R16020 GND.n11985 GND.n11983 0.01
R16021 GND.n11946 GND.n11945 0.01
R16022 GND.n11891 GND.n11890 0.01
R16023 GND.n11865 GND.n11857 0.01
R16024 GND.n12246 GND.n12237 0.01
R16025 GND.n12277 GND.n12275 0.01
R16026 GND.n12331 GND.n12330 0.01
R16027 GND.n12366 GND.n12364 0.01
R16028 GND.n13090 GND.n13088 0.01
R16029 GND.n13051 GND.n13050 0.01
R16030 GND.n12996 GND.n12995 0.01
R16031 GND.n12969 GND.n12961 0.01
R16032 GND.n7734 GND.n7726 0.01
R16033 GND.n7766 GND.n7764 0.01
R16034 GND.n7820 GND.n7819 0.01
R16035 GND.n7854 GND.n7852 0.01
R16036 GND.n8097 GND.n8095 0.01
R16037 GND.n8036 GND.n8028 0.01
R16038 GND.n6108 GND.n6059 0.01
R16039 GND.n7045 GND.n7037 0.01
R16040 GND.n7106 GND.n7104 0.01
R16041 GND.n7386 GND.n7384 0.01
R16042 GND.n7324 GND.n7322 0.01
R16043 GND.n7263 GND.n7254 0.01
R16044 GND.n15989 GND.n15980 0.01
R16045 GND.n16031 GND.n16029 0.01
R16046 GND.n16088 GND.n16087 0.01
R16047 GND.n16140 GND.n16138 0.01
R16048 GND.n1089 GND.n1087 0.01
R16049 GND.n1043 GND.n1039 0.01
R16050 GND.n982 GND.n981 0.01
R16051 GND.n936 GND.n928 0.01
R16052 GND.n9689 GND.n9680 0.01
R16053 GND.n9731 GND.n9729 0.01
R16054 GND.n9788 GND.n9787 0.01
R16055 GND.n9840 GND.n9838 0.01
R16056 GND.n1279 GND.n1271 0.01
R16057 GND.n1321 GND.n1319 0.01
R16058 GND.n1378 GND.n1377 0.01
R16059 GND.n1432 GND.n1430 0.01
R16060 GND.n10258 GND.n10256 0.01
R16061 GND.n10197 GND.n10188 0.01
R16062 GND.n8822 GND.n8820 0.01
R16063 GND.n8764 GND.n8756 0.01
R16064 GND.n8528 GND.n8526 0.01
R16065 GND.n8467 GND.n8458 0.01
R16066 GND.n10083 GND.n10081 0.01
R16067 GND.n10025 GND.n10017 0.01
R16068 GND.n9419 GND.n9291 0.01
R16069 GND.n8988 GND.n8979 0.01
R16070 GND.n9030 GND.n9028 0.01
R16071 GND.n9087 GND.n9086 0.01
R16072 GND.n9139 GND.n9137 0.01
R16073 GND.n4450 GND.n4448 0.01
R16074 GND.n4403 GND.n4399 0.01
R16075 GND.n4342 GND.n4341 0.01
R16076 GND.n4296 GND.n4288 0.01
R16077 GND.n3239 GND.n3231 0.01
R16078 GND.n3297 GND.n3295 0.01
R16079 GND.n5045 GND.n5043 0.01
R16080 GND.n4984 GND.n4976 0.01
R16081 GND.n3368 GND.n3366 0.01
R16082 GND.n3400 GND.n3395 0.01
R16083 GND.n1959 GND.n1954 0.01
R16084 GND.n4773 GND.n4771 0.01
R16085 GND.n4699 GND.n4697 0.01
R16086 GND.n4638 GND.n4630 0.01
R16087 GND.n3039 GND.n3031 0.01
R16088 GND.n3097 GND.n3095 0.01
R16089 GND.n10463 GND.n10455 0.01
R16090 GND.n10521 GND.n10519 0.01
R16091 GND.n15881 GND.n15880 0.01
R16092 GND.n14086 GND.n14084 0.01
R16093 GND.n14118 GND.n14113 0.01
R16094 GND.n14118 GND.n14116 0.01
R16095 GND.n15607 GND.n15599 0.01
R16096 GND.n15668 GND.n15666 0.01
R16097 GND.n14737 GND.n14736 0.01
R16098 GND.n14719 GND.n14474 0.01
R16099 GND.n15308 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/GATE 0.01
R16100 GND.n15298 GND.n15296 0.01
R16101 GND.n15296 GND.n15294 0.01
R16102 GND.n15170 GND.n15162 0.01
R16103 GND.n15228 GND.n15226 0.01
R16104 GND.n3870 GND.n3868 0.01
R16105 GND.n3824 GND.n3820 0.01
R16106 GND.n3763 GND.n3762 0.01
R16107 GND.n3719 GND.n3711 0.01
R16108 GND.n5708 GND.n5706 0.01
R16109 GND.n5662 GND.n5658 0.01
R16110 GND.n5601 GND.n5600 0.01
R16111 GND.n5555 GND.n5547 0.01
R16112 GND.n14494 GND.n14492 0.009
R16113 GND.n14511 GND.n14508 0.009
R16114 GND.n14507 GND.n14476 0.009
R16115 GND.n14717 GND.n14715 0.009
R16116 GND.n15452 GND.n15450 0.009
R16117 GND.n14565 GND.n14563 0.009
R16118 GND.n14569 GND.n14567 0.009
R16119 GND.n14402 GND.n14400 0.009
R16120 GND.n10579 GND.n10577 0.009
R16121 GND.n10661 GND.n10659 0.009
R16122 GND.n10666 GND.n10663 0.009
R16123 GND.n10693 GND.n10691 0.009
R16124 GND.n15530 GND.n15528 0.009
R16125 GND.n14066 GND.n14064 0.009
R16126 GND.n14062 GND.n14060 0.009
R16127 GND.n14036 GND.n14035 0.009
R16128 GND.n14123 GND.n14121 0.009
R16129 GND.n14154 GND.n14152 0.009
R16130 GND.n14158 GND.n14156 0.009
R16131 GND.n10714 GND.n10712 0.009
R16132 GND.n14165 GND.n14163 0.009
R16133 GND.n14207 GND.n14205 0.009
R16134 GND.n14211 GND.n14209 0.009
R16135 GND.n14218 GND.n10575 0.009
R16136 GND.n3616 GND.n3614 0.009
R16137 GND.n3538 GND.n3536 0.009
R16138 GND.n3534 GND.n3532 0.009
R16139 GND.n3507 GND.n3506 0.009
R16140 GND.n4791 GND.n4789 0.009
R16141 GND.n4872 GND.n4870 0.009
R16142 GND.n4877 GND.n4874 0.009
R16143 GND.n4903 GND.n4901 0.009
R16144 GND.n10787 GND.n10785 0.009
R16145 GND.n10815 GND.n10813 0.009
R16146 GND.n10819 GND.n10817 0.009
R16147 GND.n10875 GND.n10873 0.009
R16148 GND.n13887 GND.n13885 0.009
R16149 GND.n13914 GND.n13912 0.009
R16150 GND.n13918 GND.n13916 0.009
R16151 GND.n13994 GND.n13992 0.009
R16152 GND.n13866 GND.n13864 0.009
R16153 GND.n10938 GND.n10936 0.009
R16154 GND.n10934 GND.n10932 0.009
R16155 GND.n10908 GND.n10907 0.009
R16156 GND.n13727 GND.n13725 0.009
R16157 GND.n10987 GND.n10985 0.009
R16158 GND.n10983 GND.n10981 0.009
R16159 GND.n10957 GND.n10956 0.009
R16160 GND.n12714 GND.n12712 0.009
R16161 GND.n12795 GND.n12793 0.009
R16162 GND.n12800 GND.n12797 0.009
R16163 GND.n12827 GND.n12825 0.009
R16164 GND.n11448 GND.n11446 0.009
R16165 GND.n11476 GND.n11474 0.009
R16166 GND.n11480 GND.n11478 0.009
R16167 GND.n11720 GND.n11718 0.009
R16168 GND.n11509 GND.n11507 0.009
R16169 GND.n11536 GND.n11534 0.009
R16170 GND.n11540 GND.n11538 0.009
R16171 GND.n11616 GND.n11614 0.009
R16172 GND.n11108 GND.n11106 0.009
R16173 GND.n11620 GND.n11618 0.009
R16174 GND.n11625 GND.n11622 0.009
R16175 GND.n11652 GND.n11650 0.009
R16176 GND.n13321 GND.n13319 0.009
R16177 GND.n13242 GND.n13240 0.009
R16178 GND.n13238 GND.n13236 0.009
R16179 GND.n13212 GND.n13211 0.009
R16180 GND.n11323 GND.n11321 0.009
R16181 GND.n11402 GND.n11400 0.009
R16182 GND.n11407 GND.n11404 0.009
R16183 GND.n11433 GND.n11431 0.009
R16184 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE GND.n11129 0.009
R16185 GND.n8163 GND.n8161 0.009
R16186 GND.n6073 GND.n6071 0.009
R16187 GND.n6078 GND.n6075 0.009
R16188 GND.n6105 GND.n6103 0.009
R16189 GND.n8252 GND.n8250 0.009
R16190 GND.n8334 GND.n8332 0.009
R16191 GND.n8339 GND.n8336 0.009
R16192 GND.n8366 GND.n8364 0.009
R16193 GND.n5847 GND.n5845 0.009
R16194 GND.n6389 GND.n6386 0.009
R16195 GND.n6370 GND.n6368 0.009
R16196 GND.n5901 GND.n5899 0.009
R16197 GND.n5917 GND.n5915 0.009
R16198 GND.n5945 GND.n5943 0.009
R16199 GND.n5949 GND.n5947 0.009
R16200 GND.n6030 GND.n6028 0.009
R16201 GND.n6516 GND.n6514 0.009
R16202 GND.n6492 GND.n6489 0.009
R16203 GND.n6488 GND.n6486 0.009
R16204 GND.n6414 GND.n5824 0.009
R16205 GND.n6830 GND.n6828 0.009
R16206 GND.n6858 GND.n6856 0.009
R16207 GND.n6862 GND.n6860 0.009
R16208 GND.n6942 GND.n6940 0.009
R16209 GND.n6595 GND.n6593 0.009
R16210 GND.n6623 GND.n6621 0.009
R16211 GND.n6627 GND.n6625 0.009
R16212 GND.n6707 GND.n6705 0.009
R16213 GND.n6711 GND.n6709 0.009
R16214 GND.n6793 GND.n6791 0.009
R16215 GND.n6798 GND.n6795 0.009
R16216 GND.n6825 GND.n6823 0.009
R16217 GND.n7435 GND.n7433 0.009
R16218 GND.n6543 GND.n6541 0.009
R16219 GND.n6548 GND.n6545 0.009
R16220 GND.n6575 GND.n6573 0.009
R16221 GND.n7582 GND.n7580 0.009
R16222 GND.n6952 GND.n6950 0.009
R16223 GND.n6957 GND.n6954 0.009
R16224 GND.n6984 GND.n6982 0.009
R16225 GND.n16237 GND.n16236 0.009
R16226 GND.n9296 GND.n9294 0.009
R16227 GND.n9376 GND.n9374 0.009
R16228 GND.n9381 GND.n9378 0.009
R16229 GND.n9407 GND.n9405 0.009
R16230 GND.n1701 GND.n1699 0.009
R16231 GND.n1783 GND.n1781 0.009
R16232 GND.n1788 GND.n1785 0.009
R16233 GND.n1814 GND.n1812 0.009
R16234 GND.n1680 GND.n1678 0.009
R16235 GND.n1652 GND.n1649 0.009
R16236 GND.n1648 GND.n1636 0.009
R16237 GND.n9423 GND.n9421 0.009
R16238 GND.n1586 GND.n1584 0.009
R16239 GND.n1629 GND.n1627 0.009
R16240 GND.n1633 GND.n1631 0.009
R16241 GND.n1896 GND.n1894 0.009
R16242 GND.n8696 GND.n8694 0.009
R16243 GND.n8622 GND.n8620 0.009
R16244 GND.n8618 GND.n8616 0.009
R16245 GND.n8591 GND.n8590 0.009
R16246 GND.n5307 GND.n5306 0.009
R16247 GND.n2494 GND.n2492 0.009
R16248 GND.n2575 GND.n2573 0.009
R16249 GND.n2580 GND.n2577 0.009
R16250 GND.n2607 GND.n2605 0.009
R16251 GND.n2473 GND.n2471 0.009
R16252 GND.n2262 GND.n2260 0.009
R16253 GND.n2266 GND.n2264 0.009
R16254 GND.n3404 GND.n3402 0.009
R16255 GND.n3163 GND.n3161 0.009
R16256 GND.n2233 GND.n2231 0.009
R16257 GND.n2237 GND.n2235 0.009
R16258 GND.n2631 GND.n2629 0.009
R16259 GND.n3155 GND.n3153 0.009
R16260 GND.n2280 GND.n2278 0.009
R16261 GND.n2318 GND.n2315 0.009
R16262 GND.n2302 GND.n2301 0.009
R16263 GND.n5103 GND.n5101 0.009
R16264 GND.n5183 GND.n5181 0.009
R16265 GND.n5188 GND.n5185 0.009
R16266 GND.n5215 GND.n5213 0.009
R16267 GND.n2007 GND.n2005 0.009
R16268 GND.n2049 GND.n2047 0.009
R16269 GND.n2053 GND.n2051 0.009
R16270 GND.n2061 GND.n1941 0.009
R16271 GND.n1964 GND.n1962 0.009
R16272 GND.n1996 GND.n1994 0.009
R16273 GND.n2000 GND.n1998 0.009
R16274 GND.n2658 GND.n2656 0.009
R16275 GND.n2963 GND.n2961 0.009
R16276 GND.n2884 GND.n2882 0.009
R16277 GND.n2880 GND.n2878 0.009
R16278 GND.n2853 GND.n2852 0.009
R16279 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/GATE GND.n14103 0.009
R16280 GND.n15871 GND.n15869 0.009
R16281 GND.n15792 GND.n15790 0.009
R16282 GND.n15788 GND.n15786 0.009
R16283 GND.n15762 GND.n15761 0.009
R16284 GND.n15426 GND.n15424 0.009
R16285 GND.n15346 GND.n15344 0.009
R16286 GND.n15342 GND.n15340 0.009
R16287 GND.n15316 GND.n15315 0.009
R16288 GND.n14924 GND.n14922 0.009
R16289 GND.n14432 GND.n14430 0.009
R16290 GND.n14437 GND.n14434 0.009
R16291 GND.n14463 GND.n14461 0.009
R16292 GND.n15112 GND.n15110 0.009
R16293 GND.n15038 GND.n15036 0.009
R16294 GND.n15034 GND.n15032 0.009
R16295 GND.n15008 GND.n15007 0.009
R16296 GND.n16469 GND.n16467 0.009
R16297 GND.n16475 GND.n16472 0.009
R16298 GND.n16423 GND.n16421 0.009
R16299 GND.n16419 GND.n16417 0.009
R16300 GND.n16541 GND.n16539 0.009
R16301 GND.n16536 GND.n16535 0.009
R16302 GND.n16506 GND.n16505 0.009
R16303 GND.n16366 GND.n16364 0.009
R16304 GND.n16361 GND.n16360 0.009
R16305 GND.n16332 GND.n16330 0.009
R16306 GND.n16329 GND.n16327 0.009
R16307 GND.n16730 GND.n16728 0.009
R16308 GND.n16736 GND.n16733 0.009
R16309 GND.n16684 GND.n16682 0.009
R16310 GND.n16680 GND.n16678 0.009
R16311 GND.n16802 GND.n16800 0.009
R16312 GND.n16797 GND.n16796 0.009
R16313 GND.n16767 GND.n16766 0.009
R16314 GND.n16627 GND.n16625 0.009
R16315 GND.n16622 GND.n16621 0.009
R16316 GND.n16593 GND.n16591 0.009
R16317 GND.n16590 GND.n16588 0.009
R16318 GND.n16991 GND.n16989 0.009
R16319 GND.n16997 GND.n16994 0.009
R16320 GND.n16945 GND.n16943 0.009
R16321 GND.n16941 GND.n16939 0.009
R16322 GND.n17063 GND.n17061 0.009
R16323 GND.n17058 GND.n17057 0.009
R16324 GND.n17028 GND.n17027 0.009
R16325 GND.n16888 GND.n16886 0.009
R16326 GND.n16883 GND.n16882 0.009
R16327 GND.n16854 GND.n16852 0.009
R16328 GND.n16851 GND.n16849 0.009
R16329 GND.n17252 GND.n17250 0.009
R16330 GND.n17258 GND.n17255 0.009
R16331 GND.n17206 GND.n17204 0.009
R16332 GND.n17202 GND.n17200 0.009
R16333 GND.n17324 GND.n17322 0.009
R16334 GND.n17319 GND.n17318 0.009
R16335 GND.n17289 GND.n17288 0.009
R16336 GND.n17149 GND.n17147 0.009
R16337 GND.n17144 GND.n17143 0.009
R16338 GND.n17115 GND.n17113 0.009
R16339 GND.n17112 GND.n17110 0.009
R16340 GND.n17513 GND.n17511 0.009
R16341 GND.n17519 GND.n17516 0.009
R16342 GND.n17467 GND.n17465 0.009
R16343 GND.n17463 GND.n17461 0.009
R16344 GND.n17585 GND.n17583 0.009
R16345 GND.n17580 GND.n17579 0.009
R16346 GND.n17550 GND.n17549 0.009
R16347 GND.n17410 GND.n17408 0.009
R16348 GND.n17405 GND.n17404 0.009
R16349 GND.n17376 GND.n17374 0.009
R16350 GND.n17373 GND.n17371 0.009
R16351 GND.n654 GND.n652 0.009
R16352 GND.n649 GND.n648 0.009
R16353 GND.n757 GND.n755 0.009
R16354 GND.n752 GND.n750 0.009
R16355 GND.n589 GND.n587 0.009
R16356 GND.n584 GND.n582 0.009
R16357 GND.n551 GND.n549 0.009
R16358 GND.n396 GND.n394 0.009
R16359 GND.n391 GND.n390 0.009
R16360 GND.n499 GND.n497 0.009
R16361 GND.n494 GND.n492 0.009
R16362 GND.n331 GND.n329 0.009
R16363 GND.n326 GND.n324 0.009
R16364 GND.n293 GND.n291 0.009
R16365 GND.n138 GND.n136 0.009
R16366 GND.n133 GND.n132 0.009
R16367 GND.n241 GND.n239 0.009
R16368 GND.n236 GND.n234 0.009
R16369 GND.n73 GND.n71 0.009
R16370 GND.n68 GND.n66 0.009
R16371 GND.n35 GND.n33 0.009
R16372 GND.n17753 GND.n17751 0.009
R16373 GND.n17748 GND.n17747 0.009
R16374 GND.n17830 GND.n17828 0.009
R16375 GND.n17825 GND.n17823 0.009
R16376 GND.n17909 GND.n17907 0.009
R16377 GND.n17904 GND.n17902 0.009
R16378 GND.n17871 GND.n17869 0.009
R16379 GND.n10685 GND.n10682 0.008
R16380 GND.n14044 GND.n14043 0.008
R16381 GND.n3515 GND.n3514 0.008
R16382 GND.n4896 GND.n4893 0.008
R16383 GND.n10795 GND.n10794 0.008
R16384 GND.n13895 GND.n13894 0.008
R16385 GND.n10916 GND.n10915 0.008
R16386 GND.n10965 GND.n10964 0.008
R16387 GND.n12819 GND.n12816 0.008
R16388 GND.n11456 GND.n11455 0.008
R16389 GND.n11517 GND.n11516 0.008
R16390 GND.n11644 GND.n11641 0.008
R16391 GND.n13220 GND.n13219 0.008
R16392 GND.n11426 GND.n11423 0.008
R16393 GND.n6097 GND.n6094 0.008
R16394 GND.n8358 GND.n8355 0.008
R16395 GND.n5840 GND.n5837 0.008
R16396 GND.n5925 GND.n5924 0.008
R16397 GND.n6509 GND.n6506 0.008
R16398 GND.n6838 GND.n6837 0.008
R16399 GND.n6603 GND.n6602 0.008
R16400 GND.n6817 GND.n6814 0.008
R16401 GND.n6567 GND.n6564 0.008
R16402 GND.n6976 GND.n6973 0.008
R16403 GND.n9400 GND.n9397 0.008
R16404 GND.n1807 GND.n1804 0.008
R16405 GND.n8599 GND.n8598 0.008
R16406 GND.n2599 GND.n2596 0.008
R16407 GND.n2310 GND.n2309 0.008
R16408 GND.n5207 GND.n5204 0.008
R16409 GND.n2861 GND.n2860 0.008
R16410 GND.n15770 GND.n15769 0.008
R16411 GND.n15324 GND.n15323 0.008
R16412 GND.n14456 GND.n14453 0.008
R16413 GND.n15016 GND.n15015 0.008
R16414 GND.n16441 GND.n16440 0.008
R16415 GND.n16527 GND.n16526 0.008
R16416 GND.n16350 GND.n16349 0.008
R16417 GND.n16702 GND.n16701 0.008
R16418 GND.n16788 GND.n16787 0.008
R16419 GND.n16611 GND.n16610 0.008
R16420 GND.n16963 GND.n16962 0.008
R16421 GND.n17049 GND.n17048 0.008
R16422 GND.n16872 GND.n16871 0.008
R16423 GND.n17224 GND.n17223 0.008
R16424 GND.n17310 GND.n17309 0.008
R16425 GND.n17133 GND.n17132 0.008
R16426 GND.n17485 GND.n17484 0.008
R16427 GND.n17571 GND.n17570 0.008
R16428 GND.n17394 GND.n17393 0.008
R16429 GND.n16465 GND.n16464 0.008
R16430 GND.n16368 GND.n16367 0.008
R16431 GND.n16543 GND.n16542 0.008
R16432 GND.n16726 GND.n16725 0.008
R16433 GND.n16629 GND.n16628 0.008
R16434 GND.n16804 GND.n16803 0.008
R16435 GND.n16987 GND.n16986 0.008
R16436 GND.n16890 GND.n16889 0.008
R16437 GND.n17065 GND.n17064 0.008
R16438 GND.n17248 GND.n17247 0.008
R16439 GND.n17151 GND.n17150 0.008
R16440 GND.n17326 GND.n17325 0.008
R16441 GND.n17509 GND.n17508 0.008
R16442 GND.n17412 GND.n17411 0.008
R16443 GND.n17587 GND.n17586 0.008
R16444 GND.n656 GND.n655 0.008
R16445 GND.n591 GND.n590 0.008
R16446 GND.n759 GND.n758 0.008
R16447 GND.n398 GND.n397 0.008
R16448 GND.n333 GND.n332 0.008
R16449 GND.n501 GND.n500 0.008
R16450 GND.n140 GND.n139 0.008
R16451 GND.n75 GND.n74 0.008
R16452 GND.n243 GND.n242 0.008
R16453 GND.n17755 GND.n17754 0.008
R16454 GND.n17911 GND.n17910 0.008
R16455 GND.n17832 GND.n17831 0.008
R16456 GND.n14913 GND.n14911 0.008
R16457 GND.n14741 GND.n14739 0.008
R16458 GND.n6331 GND.n6329 0.008
R16459 GND.n6165 GND.n5822 0.008
R16460 GND.n12701 GND.n12699 0.008
R16461 GND.n11312 GND.n11310 0.008
R16462 GND.n11147 GND.n11006 0.008
R16463 GND.n13719 GND.n13717 0.008
R16464 GND.n13554 GND.n10717 0.008
R16465 GND.n13508 GND.n13506 0.008
R16466 GND.n12096 GND.n12094 0.008
R16467 GND.n11925 GND.n11923 0.008
R16468 GND.n11912 GND.n11910 0.008
R16469 GND.n11750 GND.n11735 0.008
R16470 GND.n12128 GND.n12126 0.008
R16471 GND.n12299 GND.n12297 0.008
R16472 GND.n12312 GND.n12310 0.008
R16473 GND.n12480 GND.n12478 0.008
R16474 GND.n13195 GND.n13193 0.008
R16475 GND.n13030 GND.n13028 0.008
R16476 GND.n13017 GND.n13015 0.008
R16477 GND.n12849 GND.n12847 0.008
R16478 GND.n7623 GND.n7621 0.008
R16479 GND.n7788 GND.n7786 0.008
R16480 GND.n7801 GND.n7799 0.008
R16481 GND.n7963 GND.n7961 0.008
R16482 GND.n8149 GND.n8147 0.008
R16483 GND.n7977 GND.n7975 0.008
R16484 GND.n8380 GND.n8377 0.008
R16485 GND.n6987 GND.n6149 0.008
R16486 GND.n7159 GND.n7157 0.008
R16487 GND.n7429 GND.n7426 0.008
R16488 GND.n7375 GND.n7373 0.008
R16489 GND.n7204 GND.n7202 0.008
R16490 GND.n1530 GND.n1529 0.008
R16491 GND.n15894 GND.n15892 0.008
R16492 GND.n16065 GND.n16063 0.008
R16493 GND.n16069 GND.n16067 0.008
R16494 GND.n16232 GND.n16230 0.008
R16495 GND.n1172 GND.n1170 0.008
R16496 GND.n1007 GND.n1005 0.008
R16497 GND.n1003 GND.n1001 0.008
R16498 GND.n834 GND.n832 0.008
R16499 GND.n9594 GND.n1174 0.008
R16500 GND.n9765 GND.n9763 0.008
R16501 GND.n9769 GND.n9767 0.008
R16502 GND.n9932 GND.n9930 0.008
R16503 GND.n1190 GND.n1176 0.008
R16504 GND.n1355 GND.n1353 0.008
R16505 GND.n1359 GND.n1357 0.008
R16506 GND.n1528 GND.n1526 0.008
R16507 GND.n10309 GND.n10307 0.008
R16508 GND.n10138 GND.n10136 0.008
R16509 GND.n8872 GND.n8870 0.008
R16510 GND.n8707 GND.n8705 0.008
R16511 GND.n8579 GND.n8577 0.008
R16512 GND.n8408 GND.n1899 0.008
R16513 GND.n10133 GND.n10131 0.008
R16514 GND.n9967 GND.n9965 0.008
R16515 GND.n9251 GND.n9249 0.008
R16516 GND.n5314 GND.n5313 0.008
R16517 GND.n8893 GND.n8891 0.008
R16518 GND.n9064 GND.n9062 0.008
R16519 GND.n9068 GND.n9066 0.008
R16520 GND.n9231 GND.n9229 0.008
R16521 GND.n4538 GND.n4536 0.008
R16522 GND.n4367 GND.n4365 0.008
R16523 GND.n4363 GND.n4361 0.008
R16524 GND.n4194 GND.n1915 0.008
R16525 GND.n3184 GND.n3182 0.008
R16526 GND.n3349 GND.n3347 0.008
R16527 GND.n5097 GND.n5095 0.008
R16528 GND.n4925 GND.n1919 0.008
R16529 GND.n4751 GND.n4749 0.008
R16530 GND.n4579 GND.n1934 0.008
R16531 GND.n2983 GND.n2981 0.008
R16532 GND.n3148 GND.n3146 0.008
R16533 GND.n10407 GND.n10395 0.008
R16534 GND.n10572 GND.n10570 0.008
R16535 GND.n15549 GND.n15547 0.008
R16536 GND.n15279 GND.n15277 0.008
R16537 GND.n3953 GND.n3951 0.008
R16538 GND.n3788 GND.n3786 0.008
R16539 GND.n3784 GND.n3782 0.008
R16540 GND.n3621 GND.n1917 0.008
R16541 GND.n5791 GND.n5789 0.008
R16542 GND.n5626 GND.n5624 0.008
R16543 GND.n5622 GND.n5620 0.008
R16544 GND.n5453 GND.n5451 0.008
R16545 GND.n16271 GND.n16270 0.008
R16546 GND.n5407 GND.n5406 0.008
R16547 GND.n540 GND.n539 0.008
R16548 GND.n282 GND.n281 0.008
R16549 GND.n24 GND.n23 0.008
R16550 GND.n17859 GND.n17858 0.008
R16551 GND.n5357 GND.n5352 0.008
R16552 GND.n16482 GND.n16481 0.008
R16553 GND.n16529 GND.n16516 0.008
R16554 GND.n16743 GND.n16742 0.008
R16555 GND.n16790 GND.n16777 0.008
R16556 GND.n17004 GND.n17003 0.008
R16557 GND.n17051 GND.n17038 0.008
R16558 GND.n17265 GND.n17264 0.008
R16559 GND.n17312 GND.n17299 0.008
R16560 GND.n17526 GND.n17525 0.008
R16561 GND.n17573 GND.n17560 0.008
R16562 GND.n16319 GND.n16318 0.008
R16563 GND.n16580 GND.n16579 0.008
R16564 GND.n16841 GND.n16840 0.008
R16565 GND.n17102 GND.n17101 0.008
R16566 GND.n17363 GND.n17362 0.008
R16567 GND.n5346 GND.n5344 0.007
R16568 GND.n9572 GND.n9571 0.007
R16569 GND.n16256 GND.n16254 0.007
R16570 GND.n5315 GND.n5312 0.007
R16571 GND.n5399 GND.n5398 0.007
R16572 GND.n701 GND.n700 0.007
R16573 GND.n732 GND.n727 0.007
R16574 GND.n443 GND.n442 0.007
R16575 GND.n474 GND.n469 0.007
R16576 GND.n185 GND.n184 0.007
R16577 GND.n216 GND.n211 0.007
R16578 GND.n17800 GND.n17799 0.007
R16579 GND.n17726 GND.n17721 0.007
R16580 GND.n5343 GND.n5342 0.007
R16581 GND.n5357 GND.n5356 0.007
R16582 GND.n9544 GND.n9543 0.007
R16583 GND.n5349 GND.n5348 0.007
R16584 GND.n14680 GND.n14678 0.007
R16585 GND.n14610 GND.n14608 0.007
R16586 GND.n10616 GND.n10614 0.007
R16587 GND.n15493 GND.n15491 0.007
R16588 GND.n14338 GND.n14336 0.007
R16589 GND.n14180 GND.n14179 0.007
R16590 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/DRAIN GND.n14159 0.007
R16591 GND.n14255 GND.n14253 0.007
R16592 GND.n3579 GND.n3577 0.007
R16593 GND.n4828 GND.n4826 0.007
R16594 GND.n2743 GND.n2742 0.007
R16595 GND.n4060 GND.n4059 0.007
R16596 GND.n10788 GND.n10787 0.007
R16597 GND.n10748 GND.n10746 0.007
R16598 GND.n13888 GND.n13887 0.007
R16599 GND.n13957 GND.n13955 0.007
R16600 GND.n13829 GND.n13827 0.007
R16601 GND.n13764 GND.n13762 0.007
R16602 GND.n12751 GND.n12749 0.007
R16603 GND.n11449 GND.n11448 0.007
R16604 GND.n11683 GND.n11681 0.007
R16605 GND.n11510 GND.n11509 0.007
R16606 GND.n11579 GND.n11577 0.007
R16607 GND.n11071 GND.n11069 0.007
R16608 GND.n13284 GND.n13282 0.007
R16609 GND.n11360 GND.n11358 0.007
R16610 GND.n13201 GND.n13196 0.007
R16611 GND.n12845 GND.n12844 0.007
R16612 GND.n8200 GND.n8198 0.007
R16613 GND.n8289 GND.n8287 0.007
R16614 GND.n8364 GND.n8362 0.007
R16615 GND.n5864 GND.n5862 0.007
R16616 GND.n5993 GND.n5991 0.007
R16617 GND.n6451 GND.n6449 0.007
R16618 GND.n6032 GND.n5827 0.007
R16619 GND.n6905 GND.n6903 0.007
R16620 GND.n6670 GND.n6668 0.007
R16621 GND.n6748 GND.n6746 0.007
R16622 GND.n7472 GND.n7470 0.007
R16623 GND.n6573 GND.n6571 0.007
R16624 GND.n7416 GND.n7413 0.007
R16625 GND.n7545 GND.n7543 0.007
R16626 GND.n16283 GND.n16282 0.007
R16627 GND.n16233 GND.n812 0.007
R16628 GND.n9333 GND.n9331 0.007
R16629 GND.n1738 GND.n1736 0.007
R16630 GND.n9460 GND.n9458 0.007
R16631 GND.n1859 GND.n1857 0.007
R16632 GND.n1601 GND.n1600 0.007
R16633 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN GND.n1568 0.007
R16634 GND.n8659 GND.n8657 0.007
R16635 GND.n8592 GND.n8591 0.007
R16636 GND.n9264 GND.n9262 0.007
R16637 GND.n2531 GND.n2529 0.007
R16638 GND.n3441 GND.n3439 0.007
R16639 GND.n2437 GND.n2435 0.007
R16640 GND.n2369 GND.n2367 0.007
R16641 GND.n5220 GND.n5217 0.007
R16642 GND.n5140 GND.n5138 0.007
R16643 GND.n3481 GND.n3480 0.007
R16644 GND.n3478 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/DRAIN 0.007
R16645 GND.n2098 GND.n2096 0.007
R16646 GND.n2178 GND.n2176 0.007
R16647 GND.n2022 GND.n2021 0.007
R16648 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/DRAIN GND.n2001 0.007
R16649 GND.n2926 GND.n2924 0.007
R16650 GND.n2854 GND.n2853 0.007
R16651 GND.n4761 GND.n4760 0.007
R16652 GND.n15834 GND.n15832 0.007
R16653 GND.n14535 GND.n14534 0.007
R16654 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/DRAIN GND.n14537
+ 0.007
R16655 GND.n15389 GND.n15387 0.007
R16656 GND.n14961 GND.n14959 0.007
R16657 GND.n15075 GND.n15073 0.007
R16658 GND.n15890 GND.n15889 0.007
R16659 GND.n5413 GND.n5412 0.007
R16660 GND.n16484 GND.n16483 0.007
R16661 GND.n16397 GND.n16396 0.007
R16662 GND.n16745 GND.n16744 0.007
R16663 GND.n16658 GND.n16657 0.007
R16664 GND.n17006 GND.n17005 0.007
R16665 GND.n16919 GND.n16918 0.007
R16666 GND.n17267 GND.n17266 0.007
R16667 GND.n17180 GND.n17179 0.007
R16668 GND.n17528 GND.n17527 0.007
R16669 GND.n17441 GND.n17440 0.007
R16670 GND.n700 GND.n699 0.007
R16671 GND.n727 GND.n726 0.007
R16672 GND.n555 GND.n553 0.007
R16673 GND.n703 GND.n702 0.007
R16674 GND.n618 GND.n617 0.007
R16675 GND.n442 GND.n441 0.007
R16676 GND.n469 GND.n468 0.007
R16677 GND.n297 GND.n295 0.007
R16678 GND.n445 GND.n444 0.007
R16679 GND.n360 GND.n359 0.007
R16680 GND.n184 GND.n183 0.007
R16681 GND.n211 GND.n210 0.007
R16682 GND.n39 GND.n37 0.007
R16683 GND.n187 GND.n186 0.007
R16684 GND.n102 GND.n101 0.007
R16685 GND.n17799 GND.n17798 0.007
R16686 GND.n17721 GND.n17720 0.007
R16687 GND.n17875 GND.n17873 0.007
R16688 GND.n17802 GND.n17801 0.007
R16689 GND.n17861 GND.n17860 0.007
R16690 GND.n5356 GND.n5355 0.007
R16691 GND.n5343 GND.n5340 0.007
R16692 GND.n10797 GND.n10795 0.006
R16693 GND.n13896 GND.n13895 0.006
R16694 GND.n10917 GND.n10916 0.006
R16695 GND.n10966 GND.n10965 0.006
R16696 GND.n12816 GND.n12815 0.006
R16697 GND.n11458 GND.n11456 0.006
R16698 GND.n11518 GND.n11517 0.006
R16699 GND.n11641 GND.n11640 0.006
R16700 GND.n13221 GND.n13220 0.006
R16701 GND.n11423 GND.n11422 0.006
R16702 GND.n6094 GND.n6093 0.006
R16703 GND.n8355 GND.n8354 0.006
R16704 GND.n5837 GND.n5836 0.006
R16705 GND.n5927 GND.n5925 0.006
R16706 GND.n6506 GND.n6505 0.006
R16707 GND.n6840 GND.n6838 0.006
R16708 GND.n6605 GND.n6603 0.006
R16709 GND.n6814 GND.n6813 0.006
R16710 GND.n6564 GND.n6563 0.006
R16711 GND.n6973 GND.n6972 0.006
R16712 GND.n9397 GND.n9396 0.006
R16713 GND.n1804 GND.n1803 0.006
R16714 GND.n8600 GND.n8599 0.006
R16715 GND.n2596 GND.n2595 0.006
R16716 GND.n2311 GND.n2310 0.006
R16717 GND.n5204 GND.n5203 0.006
R16718 GND.n4893 GND.n4892 0.006
R16719 GND.n3516 GND.n3515 0.006
R16720 GND.n2862 GND.n2861 0.006
R16721 GND.n14045 GND.n14044 0.006
R16722 GND.n10682 GND.n10681 0.006
R16723 GND.n15771 GND.n15770 0.006
R16724 GND.n15325 GND.n15324 0.006
R16725 GND.n14453 GND.n14452 0.006
R16726 GND.n15017 GND.n15016 0.006
R16727 GND.n16351 GND.n16350 0.006
R16728 GND.n16442 GND.n16441 0.006
R16729 GND.n16528 GND.n16527 0.006
R16730 GND.n16612 GND.n16611 0.006
R16731 GND.n16703 GND.n16702 0.006
R16732 GND.n16789 GND.n16788 0.006
R16733 GND.n16873 GND.n16872 0.006
R16734 GND.n16964 GND.n16963 0.006
R16735 GND.n17050 GND.n17049 0.006
R16736 GND.n17134 GND.n17133 0.006
R16737 GND.n17225 GND.n17224 0.006
R16738 GND.n17311 GND.n17310 0.006
R16739 GND.n17395 GND.n17394 0.006
R16740 GND.n17486 GND.n17485 0.006
R16741 GND.n17572 GND.n17571 0.006
R16742 GND.n685 GND.n683 0.006
R16743 GND.n427 GND.n425 0.006
R16744 GND.n169 GND.n167 0.006
R16745 GND.n17784 GND.n17782 0.006
R16746 GND.n731 GND.n729 0.006
R16747 GND.n473 GND.n471 0.006
R16748 GND.n215 GND.n213 0.006
R16749 GND.n17725 GND.n17723 0.006
R16750 GND.n16510 GND.n16508 0.006
R16751 GND.n16771 GND.n16769 0.006
R16752 GND.n17032 GND.n17030 0.006
R16753 GND.n17293 GND.n17291 0.006
R16754 GND.n17554 GND.n17552 0.006
R16755 GND.n16302 GND.n16301 0.006
R16756 GND.n9526 GND.n9524 0.006
R16757 GND.n5388 GND.n5387 0.006
R16758 GND.n9571 GND.n1530 0.006
R16759 GND.n9553 GND.n9552 0.006
R16760 GND.n1538 GND.n1533 0.006
R16761 GND.n16256 GND.n16255 0.006
R16762 GND.n16266 GND.n16265 0.006
R16763 GND.n16284 GND.n16283 0.006
R16764 GND.n16281 GND.n16280 0.006
R16765 GND.n5315 GND.n5314 0.006
R16766 GND.n5326 GND.n5325 0.006
R16767 GND.n5259 GND.n5254 0.006
R16768 GND.n5377 GND.n5376 0.006
R16769 GND.n5402 GND.n5401 0.006
R16770 GND.n5414 GND.n5413 0.006
R16771 GND.n5411 GND.n5410 0.006
R16772 GND.n16398 GND.n16320 0.006
R16773 GND.n16659 GND.n16581 0.006
R16774 GND.n16920 GND.n16842 0.006
R16775 GND.n17181 GND.n17103 0.006
R16776 GND.n17442 GND.n17364 0.006
R16777 GND.n619 GND.n541 0.006
R16778 GND.n361 GND.n283 0.006
R16779 GND.n103 GND.n25 0.006
R16780 GND.n17705 GND.n0 0.006
R16781 GND.n9560 GND.n9559 0.006
R16782 GND.n1544 GND.n1543 0.006
R16783 GND.n1546 GND.n1545 0.006
R16784 GND.n9569 GND.n9568 0.006
R16785 GND.n16297 GND.n16296 0.006
R16786 GND.n16292 GND.n16291 0.006
R16787 GND.n16259 GND.n16258 0.006
R16788 GND.n16294 GND.n16293 0.006
R16789 GND.n5333 GND.n5332 0.006
R16790 GND.n5268 GND.n5267 0.006
R16791 GND.n5270 GND.n5269 0.006
R16792 GND.n5318 GND.n5317 0.006
R16793 GND.n5380 GND.n5379 0.006
R16794 GND.n5385 GND.n5384 0.006
R16795 GND.n799 GND.n794 0.006
R16796 GND.n16511 GND.n16506 0.006
R16797 GND.n16772 GND.n16767 0.006
R16798 GND.n17033 GND.n17028 0.006
R16799 GND.n17294 GND.n17289 0.006
R16800 GND.n17555 GND.n17550 0.006
R16801 GND.n16570 GND.n16569 0.006
R16802 GND.n16831 GND.n16830 0.006
R16803 GND.n17092 GND.n17091 0.006
R16804 GND.n17353 GND.n17352 0.006
R16805 GND.n17614 GND.n17613 0.006
R16806 GND.n786 GND.n785 0.006
R16807 GND.n528 GND.n527 0.006
R16808 GND.n270 GND.n269 0.006
R16809 GND.n17804 GND.n17803 0.006
R16810 GND.n5348 GND.n5347 0.006
R16811 GND.n14849 GND.n14847 0.006
R16812 GND.n14813 GND.n14804 0.006
R16813 GND.n6269 GND.n6267 0.006
R16814 GND.n6235 GND.n6227 0.006
R16815 GND.n12637 GND.n12635 0.006
R16816 GND.n12601 GND.n12592 0.006
R16817 GND.n11250 GND.n11248 0.006
R16818 GND.n11216 GND.n11208 0.006
R16819 GND.n13657 GND.n13655 0.006
R16820 GND.n13623 GND.n13615 0.006
R16821 GND.n13408 GND.n13399 0.006
R16822 GND.n13444 GND.n13442 0.006
R16823 GND.n11972 GND.n11970 0.006
R16824 GND.n11950 GND.n11949 0.006
R16825 GND.n11887 GND.n11886 0.006
R16826 GND.n11870 GND.n11869 0.006
R16827 GND.n12263 GND.n12250 0.006
R16828 GND.n12272 GND.n12271 0.006
R16829 GND.n12335 GND.n12334 0.006
R16830 GND.n12354 GND.n12352 0.006
R16831 GND.n13078 GND.n13076 0.006
R16832 GND.n13056 GND.n13055 0.006
R16833 GND.n12992 GND.n12991 0.006
R16834 GND.n12974 GND.n12973 0.006
R16835 GND.n7751 GND.n7738 0.006
R16836 GND.n7761 GND.n7759 0.006
R16837 GND.n7824 GND.n7823 0.006
R16838 GND.n7842 GND.n7840 0.006
R16839 GND.n8085 GND.n8083 0.006
R16840 GND.n8049 GND.n8040 0.006
R16841 GND.n7058 GND.n7049 0.006
R16842 GND.n7094 GND.n7092 0.006
R16843 GND.n7311 GND.n7309 0.006
R16844 GND.n7275 GND.n7267 0.006
R16845 GND.n9559 GND.n9558 0.006
R16846 GND.n16006 GND.n15993 0.006
R16847 GND.n16023 GND.n16021 0.006
R16848 GND.n16091 GND.n16090 0.006
R16849 GND.n16128 GND.n16126 0.006
R16850 GND.n1077 GND.n1075 0.006
R16851 GND.n1051 GND.n1047 0.006
R16852 GND.n979 GND.n978 0.006
R16853 GND.n949 GND.n940 0.006
R16854 GND.n9706 GND.n9693 0.006
R16855 GND.n9723 GND.n9721 0.006
R16856 GND.n9791 GND.n9790 0.006
R16857 GND.n9828 GND.n9826 0.006
R16858 GND.n1296 GND.n1283 0.006
R16859 GND.n1313 GND.n1311 0.006
R16860 GND.n1381 GND.n1380 0.006
R16861 GND.n1420 GND.n1418 0.006
R16862 GND.n10245 GND.n10243 0.006
R16863 GND.n10209 GND.n10201 0.006
R16864 GND.n8810 GND.n8808 0.006
R16865 GND.n8776 GND.n8768 0.006
R16866 GND.n8515 GND.n8513 0.006
R16867 GND.n8479 GND.n8471 0.006
R16868 GND.n10071 GND.n10069 0.006
R16869 GND.n10037 GND.n10029 0.006
R16870 GND.n5332 GND.n5331 0.006
R16871 GND.n9005 GND.n8992 0.006
R16872 GND.n9022 GND.n9020 0.006
R16873 GND.n9090 GND.n9089 0.006
R16874 GND.n9127 GND.n9125 0.006
R16875 GND.n4437 GND.n4435 0.006
R16876 GND.n4411 GND.n4407 0.006
R16877 GND.n4339 GND.n4338 0.006
R16878 GND.n4309 GND.n4300 0.006
R16879 GND.n3251 GND.n3243 0.006
R16880 GND.n3285 GND.n3283 0.006
R16881 GND.n5033 GND.n5031 0.006
R16882 GND.n4997 GND.n4988 0.006
R16883 GND.n4687 GND.n4685 0.006
R16884 GND.n4651 GND.n4642 0.006
R16885 GND.n3051 GND.n3043 0.006
R16886 GND.n3085 GND.n3083 0.006
R16887 GND.n10475 GND.n10467 0.006
R16888 GND.n10509 GND.n10507 0.006
R16889 GND.n15620 GND.n15611 0.006
R16890 GND.n15656 GND.n15654 0.006
R16891 GND.n15182 GND.n15174 0.006
R16892 GND.n15216 GND.n15214 0.006
R16893 GND.n3858 GND.n3856 0.006
R16894 GND.n3832 GND.n3828 0.006
R16895 GND.n3760 GND.n3759 0.006
R16896 GND.n3731 GND.n3723 0.006
R16897 GND.n5696 GND.n5694 0.006
R16898 GND.n5670 GND.n5666 0.006
R16899 GND.n5598 GND.n5597 0.006
R16900 GND.n5568 GND.n5559 0.006
R16901 GND.n5401 GND.n5400 0.006
R16902 GND.n1539 GND.n1538 0.006
R16903 GND.n5260 GND.n5259 0.006
R16904 GND.n1563 GND.n1562 0.006
R16905 GND.n5288 GND.n5287 0.006
R16906 GND.n5371 GND.n5368 0.006
R16907 GND.n16249 GND.n16248 0.006
R16908 GND.n5423 GND.n5251 0.006
R16909 GND.n9543 GND.n9542 0.006
R16910 GND.n17656 GND.n17655 0.005
R16911 GND.n17664 GND.n17663 0.005
R16912 GND.n16266 GND.n16264 0.005
R16913 GND.n16281 GND.n16278 0.005
R16914 GND.n9531 GND.n9530 0.005
R16915 GND.n9540 GND.n9538 0.005
R16916 GND.n5402 GND.n5399 0.005
R16917 GND.n5411 GND.n5409 0.005
R16918 GND.n5347 GND.n5346 0.005
R16919 GND.n5352 GND.n5349 0.005
R16920 GND.n2737 GND.n2736 0.005
R16921 GND.n4051 GND.n4050 0.005
R16922 GND.n6047 GND.n6043 0.005
R16923 GND.n7403 GND.n7400 0.005
R16924 GND.n1543 GND.n1542 0.005
R16925 GND.n16291 GND.n16290 0.005
R16926 GND.n9278 GND.n9275 0.005
R16927 GND.n5267 GND.n5266 0.005
R16928 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/GATE GND.n3385 0.005
R16929 GND.n5384 GND.n5383 0.005
R16930 GND.n650 GND.n649 0.005
R16931 GND.n645 GND.n644 0.005
R16932 GND.n579 GND.n578 0.005
R16933 GND.n585 GND.n584 0.005
R16934 GND.n747 GND.n746 0.005
R16935 GND.n753 GND.n752 0.005
R16936 GND.n392 GND.n391 0.005
R16937 GND.n387 GND.n386 0.005
R16938 GND.n321 GND.n320 0.005
R16939 GND.n327 GND.n326 0.005
R16940 GND.n489 GND.n488 0.005
R16941 GND.n495 GND.n494 0.005
R16942 GND.n134 GND.n133 0.005
R16943 GND.n129 GND.n128 0.005
R16944 GND.n63 GND.n62 0.005
R16945 GND.n69 GND.n68 0.005
R16946 GND.n231 GND.n230 0.005
R16947 GND.n237 GND.n236 0.005
R16948 GND.n17749 GND.n17748 0.005
R16949 GND.n17744 GND.n17743 0.005
R16950 GND.n17899 GND.n17898 0.005
R16951 GND.n17905 GND.n17904 0.005
R16952 GND.n17820 GND.n17819 0.005
R16953 GND.n17826 GND.n17825 0.005
R16954 GND.n5423 GND.n5422 0.005
R16955 GND.n9542 GND.n9541 0.005
R16956 GND.n798 GND.n797 0.004
R16957 GND.n16276 GND.n16275 0.004
R16958 GND.n6116 GND.n6111 0.004
R16959 GND.n7382 GND.n6154 0.004
R16960 GND.n9417 GND.n9414 0.004
R16961 GND.n14642 GND.n14640 0.004
R16962 GND.n14646 GND.n14644 0.004
R16963 GND.n14576 GND.n14574 0.004
R16964 GND.n14580 GND.n14578 0.004
R16965 GND.n10651 GND.n10649 0.004
R16966 GND.n10656 GND.n10653 0.004
R16967 GND.n14076 GND.n14074 0.004
R16968 GND.n14072 GND.n14070 0.004
R16969 GND.n14298 GND.n14296 0.004
R16970 GND.n14303 GND.n14301 0.004
R16971 GND.n14177 GND.n14176 0.004
R16972 GND.n14183 GND.n14182 0.004
R16973 GND.n14306 GND.n14299 0.004
R16974 GND.n14307 GND.n14306 0.004
R16975 GND.n14315 GND.n14307 0.004
R16976 GND.n14358 GND.n14315 0.004
R16977 GND.n14289 GND.n14286 0.004
R16978 GND.n14285 GND.n14283 0.004
R16979 GND.n3548 GND.n3546 0.004
R16980 GND.n3544 GND.n3542 0.004
R16981 GND.n4862 GND.n4860 0.004
R16982 GND.n4867 GND.n4864 0.004
R16983 GND.n10825 GND.n10823 0.004
R16984 GND.n10829 GND.n10827 0.004
R16985 GND.n13924 GND.n13922 0.004
R16986 GND.n13928 GND.n13926 0.004
R16987 GND.n10948 GND.n10946 0.004
R16988 GND.n10944 GND.n10942 0.004
R16989 GND.n10997 GND.n10995 0.004
R16990 GND.n10993 GND.n10991 0.004
R16991 GND.n12785 GND.n12783 0.004
R16992 GND.n12790 GND.n12787 0.004
R16993 GND.n11486 GND.n11484 0.004
R16994 GND.n11490 GND.n11488 0.004
R16995 GND.n11546 GND.n11544 0.004
R16996 GND.n11550 GND.n11548 0.004
R16997 GND.n11027 GND.n11025 0.004
R16998 GND.n11023 GND.n11021 0.004
R16999 GND.n13252 GND.n13250 0.004
R17000 GND.n13248 GND.n13246 0.004
R17001 GND.n11392 GND.n11390 0.004
R17002 GND.n11397 GND.n11394 0.004
R17003 GND.n6063 GND.n6061 0.004
R17004 GND.n6068 GND.n6065 0.004
R17005 GND.n8324 GND.n8322 0.004
R17006 GND.n8329 GND.n8326 0.004
R17007 GND.n6376 GND.n6374 0.004
R17008 GND.n6380 GND.n6378 0.004
R17009 GND.n5955 GND.n5953 0.004
R17010 GND.n5959 GND.n5957 0.004
R17011 GND.n6483 GND.n6480 0.004
R17012 GND.n6479 GND.n6477 0.004
R17013 GND.n7973 GND.n7972 0.004
R17014 GND.n6868 GND.n6866 0.004
R17015 GND.n6872 GND.n6870 0.004
R17016 GND.n6633 GND.n6631 0.004
R17017 GND.n6637 GND.n6635 0.004
R17018 GND.n6783 GND.n6781 0.004
R17019 GND.n6788 GND.n6785 0.004
R17020 GND.n6533 GND.n6531 0.004
R17021 GND.n6538 GND.n6535 0.004
R17022 GND.n7592 GND.n7587 0.004
R17023 GND.n7518 GND.n7516 0.004
R17024 GND.n6947 GND.n6944 0.004
R17025 GND.n1554 GND.n1547 0.004
R17026 GND.n1554 GND.n1553 0.004
R17027 GND.n1551 GND.n1550 0.004
R17028 GND.n9561 GND.n9556 0.004
R17029 GND.n1562 GND.n1561 0.004
R17030 GND.n16304 GND.n16295 0.004
R17031 GND.n16304 GND.n16303 0.004
R17032 GND.n16300 GND.n16299 0.004
R17033 GND.n16280 GND.n16279 0.004
R17034 GND.n9366 GND.n9364 0.004
R17035 GND.n9371 GND.n9368 0.004
R17036 GND.n1773 GND.n1771 0.004
R17037 GND.n1778 GND.n1775 0.004
R17038 GND.n9494 GND.n9491 0.004
R17039 GND.n9490 GND.n9488 0.004
R17040 GND.n1821 GND.n1819 0.004
R17041 GND.n1825 GND.n1823 0.004
R17042 GND.n1598 GND.n1597 0.004
R17043 GND.n1604 GND.n1603 0.004
R17044 GND.n9499 GND.n9498 0.004
R17045 GND.n9500 GND.n9499 0.004
R17046 GND.n9501 GND.n9500 0.004
R17047 GND.n9502 GND.n9501 0.004
R17048 GND.n9519 GND.n9518 0.004
R17049 GND.n8632 GND.n8630 0.004
R17050 GND.n8628 GND.n8626 0.004
R17051 GND.n9963 GND.n9962 0.004
R17052 GND.n5279 GND.n5272 0.004
R17053 GND.n5279 GND.n5278 0.004
R17054 GND.n5276 GND.n5275 0.004
R17055 GND.n5334 GND.n5329 0.004
R17056 GND.n5287 GND.n5286 0.004
R17057 GND.n2565 GND.n2563 0.004
R17058 GND.n2570 GND.n2567 0.004
R17059 GND.n3475 GND.n3472 0.004
R17060 GND.n3471 GND.n3469 0.004
R17061 GND.n2399 GND.n2397 0.004
R17062 GND.n2404 GND.n2402 0.004
R17063 GND.n2289 GND.n2287 0.004
R17064 GND.n2285 GND.n2284 0.004
R17065 GND.n5173 GND.n5171 0.004
R17066 GND.n5178 GND.n5175 0.004
R17067 GND.n2460 GND.n2393 0.004
R17068 GND.n3487 GND.n3486 0.004
R17069 GND.n3484 GND.n3483 0.004
R17070 GND.n2407 GND.n2400 0.004
R17071 GND.n2408 GND.n2407 0.004
R17072 GND.n2417 GND.n2408 0.004
R17073 GND.n2457 GND.n2417 0.004
R17074 GND.n2132 GND.n2129 0.004
R17075 GND.n2128 GND.n2126 0.004
R17076 GND.n2141 GND.n2139 0.004
R17077 GND.n2146 GND.n2144 0.004
R17078 GND.n2019 GND.n2018 0.004
R17079 GND.n2025 GND.n2024 0.004
R17080 GND.n2149 GND.n2142 0.004
R17081 GND.n2150 GND.n2149 0.004
R17082 GND.n2158 GND.n2150 0.004
R17083 GND.n2198 GND.n2158 0.004
R17084 GND.n3496 GND.n3495 0.004
R17085 GND.n2894 GND.n2892 0.004
R17086 GND.n2890 GND.n2888 0.004
R17087 GND.n4784 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/GATE 0.004
R17088 GND.n15802 GND.n15800 0.004
R17089 GND.n15798 GND.n15796 0.004
R17090 GND.n14529 GND.n14368 0.004
R17091 GND.n14532 GND.n14531 0.004
R17092 GND.n14634 GND.n14633 0.004
R17093 GND.n14633 GND.n14632 0.004
R17094 GND.n14632 GND.n14631 0.004
R17095 GND.n14631 GND.n14630 0.004
R17096 GND.n15356 GND.n15354 0.004
R17097 GND.n15352 GND.n15350 0.004
R17098 GND.n14422 GND.n14420 0.004
R17099 GND.n14427 GND.n14424 0.004
R17100 GND.n15048 GND.n15046 0.004
R17101 GND.n15044 GND.n15042 0.004
R17102 GND.n5379 GND.n5378 0.004
R17103 GND.n5391 GND.n5390 0.004
R17104 GND.n5390 GND.n5389 0.004
R17105 GND.n16458 GND.n16456 0.004
R17106 GND.n16463 GND.n16460 0.004
R17107 GND.n16434 GND.n16432 0.004
R17108 GND.n16552 GND.n16550 0.004
R17109 GND.n16548 GND.n16546 0.004
R17110 GND.n16520 GND.n16518 0.004
R17111 GND.n16377 GND.n16375 0.004
R17112 GND.n16373 GND.n16371 0.004
R17113 GND.n16343 GND.n16341 0.004
R17114 GND.n16572 GND.n16491 0.004
R17115 GND.n16573 GND.n16572 0.004
R17116 GND.n16406 GND.n16405 0.004
R17117 GND.n16405 GND.n16316 0.004
R17118 GND.n16719 GND.n16717 0.004
R17119 GND.n16724 GND.n16721 0.004
R17120 GND.n16695 GND.n16693 0.004
R17121 GND.n16813 GND.n16811 0.004
R17122 GND.n16809 GND.n16807 0.004
R17123 GND.n16781 GND.n16779 0.004
R17124 GND.n16638 GND.n16636 0.004
R17125 GND.n16634 GND.n16632 0.004
R17126 GND.n16604 GND.n16602 0.004
R17127 GND.n16833 GND.n16752 0.004
R17128 GND.n16834 GND.n16833 0.004
R17129 GND.n16667 GND.n16666 0.004
R17130 GND.n16666 GND.n16577 0.004
R17131 GND.n16980 GND.n16978 0.004
R17132 GND.n16985 GND.n16982 0.004
R17133 GND.n16956 GND.n16954 0.004
R17134 GND.n17074 GND.n17072 0.004
R17135 GND.n17070 GND.n17068 0.004
R17136 GND.n17042 GND.n17040 0.004
R17137 GND.n16899 GND.n16897 0.004
R17138 GND.n16895 GND.n16893 0.004
R17139 GND.n16865 GND.n16863 0.004
R17140 GND.n17094 GND.n17013 0.004
R17141 GND.n17095 GND.n17094 0.004
R17142 GND.n16928 GND.n16927 0.004
R17143 GND.n16927 GND.n16838 0.004
R17144 GND.n17241 GND.n17239 0.004
R17145 GND.n17246 GND.n17243 0.004
R17146 GND.n17217 GND.n17215 0.004
R17147 GND.n17335 GND.n17333 0.004
R17148 GND.n17331 GND.n17329 0.004
R17149 GND.n17303 GND.n17301 0.004
R17150 GND.n17160 GND.n17158 0.004
R17151 GND.n17156 GND.n17154 0.004
R17152 GND.n17126 GND.n17124 0.004
R17153 GND.n17355 GND.n17274 0.004
R17154 GND.n17356 GND.n17355 0.004
R17155 GND.n17189 GND.n17188 0.004
R17156 GND.n17188 GND.n17099 0.004
R17157 GND.n17502 GND.n17500 0.004
R17158 GND.n17507 GND.n17504 0.004
R17159 GND.n17478 GND.n17476 0.004
R17160 GND.n17596 GND.n17594 0.004
R17161 GND.n17592 GND.n17590 0.004
R17162 GND.n17564 GND.n17562 0.004
R17163 GND.n17421 GND.n17419 0.004
R17164 GND.n17417 GND.n17415 0.004
R17165 GND.n17387 GND.n17385 0.004
R17166 GND.n17616 GND.n17535 0.004
R17167 GND.n17617 GND.n17616 0.004
R17168 GND.n17450 GND.n17449 0.004
R17169 GND.n17449 GND.n17360 0.004
R17170 GND.n17662 GND.n17661 0.004
R17171 GND.n665 GND.n663 0.004
R17172 GND.n661 GND.n659 0.004
R17173 GND.n768 GND.n766 0.004
R17174 GND.n764 GND.n762 0.004
R17175 GND.n599 GND.n597 0.004
R17176 GND.n595 GND.n594 0.004
R17177 GND.n790 GND.n710 0.004
R17178 GND.n791 GND.n790 0.004
R17179 GND.n627 GND.n626 0.004
R17180 GND.n626 GND.n537 0.004
R17181 GND.n407 GND.n405 0.004
R17182 GND.n403 GND.n401 0.004
R17183 GND.n510 GND.n508 0.004
R17184 GND.n506 GND.n504 0.004
R17185 GND.n341 GND.n339 0.004
R17186 GND.n337 GND.n336 0.004
R17187 GND.n532 GND.n452 0.004
R17188 GND.n533 GND.n532 0.004
R17189 GND.n369 GND.n368 0.004
R17190 GND.n368 GND.n279 0.004
R17191 GND.n149 GND.n147 0.004
R17192 GND.n145 GND.n143 0.004
R17193 GND.n252 GND.n250 0.004
R17194 GND.n248 GND.n246 0.004
R17195 GND.n83 GND.n81 0.004
R17196 GND.n79 GND.n78 0.004
R17197 GND.n274 GND.n194 0.004
R17198 GND.n275 GND.n274 0.004
R17199 GND.n111 GND.n110 0.004
R17200 GND.n110 GND.n21 0.004
R17201 GND.n17764 GND.n17762 0.004
R17202 GND.n17760 GND.n17758 0.004
R17203 GND.n17841 GND.n17839 0.004
R17204 GND.n17837 GND.n17835 0.004
R17205 GND.n17919 GND.n17917 0.004
R17206 GND.n17915 GND.n17914 0.004
R17207 GND.n9 GND.n8 0.004
R17208 GND.n17700 GND.n17695 0.004
R17209 GND.n17700 GND.n17699 0.004
R17210 GND.n17667 GND 0.004
R17211 GND.n10691 GND.n10689 0.004
R17212 GND.n14037 GND.n14036 0.004
R17213 GND.n10909 GND.n10908 0.004
R17214 GND.n10958 GND.n10957 0.004
R17215 GND.n12825 GND.n12823 0.004
R17216 GND.n11650 GND.n11648 0.004
R17217 GND.n13213 GND.n13212 0.004
R17218 GND.n11431 GND.n11430 0.004
R17219 GND.n6103 GND.n6101 0.004
R17220 GND.n5845 GND.n5844 0.004
R17221 GND.n5918 GND.n5917 0.004
R17222 GND.n6514 GND.n6513 0.004
R17223 GND.n6831 GND.n6830 0.004
R17224 GND.n6596 GND.n6595 0.004
R17225 GND.n6823 GND.n6821 0.004
R17226 GND.n6982 GND.n6980 0.004
R17227 GND.n9405 GND.n9404 0.004
R17228 GND.n1812 GND.n1811 0.004
R17229 GND.n2605 GND.n2603 0.004
R17230 GND.n2303 GND.n2302 0.004
R17231 GND.n5213 GND.n5211 0.004
R17232 GND.n4901 GND.n4900 0.004
R17233 GND.n3508 GND.n3507 0.004
R17234 GND.n15763 GND.n15762 0.004
R17235 GND.n15317 GND.n15316 0.004
R17236 GND.n14461 GND.n14460 0.004
R17237 GND.n15009 GND.n15008 0.004
R17238 GND.n16477 GND.n16476 0.004
R17239 GND.n16357 GND.n16356 0.004
R17240 GND.n16362 GND.n16361 0.004
R17241 GND.n16537 GND.n16536 0.004
R17242 GND.n16472 GND.n16470 0.004
R17243 GND.n16738 GND.n16737 0.004
R17244 GND.n16618 GND.n16617 0.004
R17245 GND.n16623 GND.n16622 0.004
R17246 GND.n16798 GND.n16797 0.004
R17247 GND.n16733 GND.n16731 0.004
R17248 GND.n16999 GND.n16998 0.004
R17249 GND.n16879 GND.n16878 0.004
R17250 GND.n16884 GND.n16883 0.004
R17251 GND.n17059 GND.n17058 0.004
R17252 GND.n16994 GND.n16992 0.004
R17253 GND.n17260 GND.n17259 0.004
R17254 GND.n17140 GND.n17139 0.004
R17255 GND.n17145 GND.n17144 0.004
R17256 GND.n17320 GND.n17319 0.004
R17257 GND.n17255 GND.n17253 0.004
R17258 GND.n17521 GND.n17520 0.004
R17259 GND.n17401 GND.n17400 0.004
R17260 GND.n17406 GND.n17405 0.004
R17261 GND.n17581 GND.n17580 0.004
R17262 GND.n17516 GND.n17514 0.004
R17263 GND.n572 GND.n571 0.004
R17264 GND.n740 GND.n739 0.004
R17265 GND.n638 GND.n637 0.004
R17266 GND.n314 GND.n313 0.004
R17267 GND.n482 GND.n481 0.004
R17268 GND.n380 GND.n379 0.004
R17269 GND.n56 GND.n55 0.004
R17270 GND.n224 GND.n223 0.004
R17271 GND.n122 GND.n121 0.004
R17272 GND.n17892 GND.n17891 0.004
R17273 GND.n17813 GND.n17812 0.004
R17274 GND.n17737 GND.n17736 0.004
R17275 GND.n14186 GND.n14185 0.004
R17276 GND.n1669 GND.n1668 0.004
R17277 GND.n2241 GND.n2205 0.004
R17278 GND.n2028 GND.n2027 0.004
R17279 GND.n14528 GND.n14527 0.004
R17280 GND.n799 GND.n798 0.004
R17281 GND.n14544 GND.n14542 0.003
R17282 GND.n14133 GND.n14132 0.003
R17283 GND.n1608 GND.n1606 0.003
R17284 GND.n2212 GND.n2210 0.003
R17285 GND.n1975 GND.n1973 0.003
R17286 GND.n17665 GND.n799 0.003
R17287 GND.n14175 GND.n14174 0.003
R17288 GND.n14176 GND.n14175 0.003
R17289 GND.n14184 GND.n14177 0.003
R17290 GND.n14184 GND.n14183 0.003
R17291 GND.n14299 GND.n14078 0.003
R17292 GND.n14359 GND.n14358 0.003
R17293 GND.n10781 GND.n10779 0.003
R17294 GND.n13879 GND.n13877 0.003
R17295 GND.n13528 GND.n13520 0.003
R17296 GND.n13541 GND.n13539 0.003
R17297 GND.n8247 GND.n8245 0.003
R17298 GND.n5909 GND.n5833 0.003
R17299 GND.n8377 GND.n8375 0.003
R17300 GND.n8369 GND.n5827 0.003
R17301 GND.n7426 GND.n7424 0.003
R17302 GND.n7418 GND.n7416 0.003
R17303 GND.n7194 GND.n7192 0.003
R17304 GND.n7181 GND.n7173 0.003
R17305 GND.n9573 GND.n9572 0.003
R17306 GND.n9555 GND.n9554 0.003
R17307 GND.n1596 GND.n1595 0.003
R17308 GND.n1597 GND.n1596 0.003
R17309 GND.n1605 GND.n1598 0.003
R17310 GND.n1605 GND.n1604 0.003
R17311 GND.n9498 GND.n9497 0.003
R17312 GND.n9503 GND.n9502 0.003
R17313 GND.n1580 GND.n1578 0.003
R17314 GND.n1694 GND.n1686 0.003
R17315 GND.n9257 GND.n9251 0.003
R17316 GND.n9262 GND.n9259 0.003
R17317 GND.n5312 GND.n5311 0.003
R17318 GND.n5328 GND.n5327 0.003
R17319 GND.n3174 GND.n3172 0.003
R17320 GND.n2487 GND.n2479 0.003
R17321 GND.n3489 GND.n3488 0.003
R17322 GND.n3488 GND.n3487 0.003
R17323 GND.n3486 GND.n3485 0.003
R17324 GND.n3485 GND.n3484 0.003
R17325 GND.n2400 GND.n2239 0.003
R17326 GND.n2458 GND.n2457 0.003
R17327 GND.n2017 GND.n2016 0.003
R17328 GND.n2018 GND.n2017 0.003
R17329 GND.n2026 GND.n2019 0.003
R17330 GND.n2026 GND.n2025 0.003
R17331 GND.n2142 GND.n1944 0.003
R17332 GND.n2199 GND.n2198 0.003
R17333 GND.n2668 GND.n2666 0.003
R17334 GND.n4917 GND.n4915 0.003
R17335 GND.n15749 GND.n15747 0.003
R17336 GND.n15736 GND.n15728 0.003
R17337 GND.n15455 GND.n15454 0.003
R17338 GND.n15454 GND.n14368 0.003
R17339 GND.n14530 GND.n14529 0.003
R17340 GND.n14531 GND.n14530 0.003
R17341 GND.n14635 GND.n14634 0.003
R17342 GND.n14630 GND.n14629 0.003
R17343 GND.n14488 GND.n14486 0.003
R17344 GND.n15439 GND.n15437 0.003
R17345 GND.n5253 GND.n5252 0.003
R17346 GND.n16486 GND.n16485 0.003
R17347 GND.n16571 GND.n16492 0.003
R17348 GND.n16404 GND.n16401 0.003
R17349 GND.n16400 GND.n16399 0.003
R17350 GND.n16489 GND.n16488 0.003
R17351 GND.n16314 GND.n16313 0.003
R17352 GND.n16747 GND.n16746 0.003
R17353 GND.n16832 GND.n16753 0.003
R17354 GND.n16665 GND.n16662 0.003
R17355 GND.n16661 GND.n16660 0.003
R17356 GND.n16750 GND.n16749 0.003
R17357 GND.n16575 GND.n16574 0.003
R17358 GND.n17008 GND.n17007 0.003
R17359 GND.n17093 GND.n17014 0.003
R17360 GND.n16926 GND.n16923 0.003
R17361 GND.n16922 GND.n16921 0.003
R17362 GND.n17011 GND.n17010 0.003
R17363 GND.n16836 GND.n16835 0.003
R17364 GND.n17269 GND.n17268 0.003
R17365 GND.n17354 GND.n17275 0.003
R17366 GND.n17187 GND.n17184 0.003
R17367 GND.n17183 GND.n17182 0.003
R17368 GND.n17272 GND.n17271 0.003
R17369 GND.n17097 GND.n17096 0.003
R17370 GND.n17530 GND.n17529 0.003
R17371 GND.n17615 GND.n17536 0.003
R17372 GND.n17448 GND.n17445 0.003
R17373 GND.n17444 GND.n17443 0.003
R17374 GND.n17533 GND.n17532 0.003
R17375 GND.n17358 GND.n17357 0.003
R17376 GND.n17619 GND.n17618 0.003
R17377 GND.n17620 GND.n17619 0.003
R17378 GND.n17621 GND.n17620 0.003
R17379 GND.n17622 GND.n17621 0.003
R17380 GND.n17623 GND.n17622 0.003
R17381 GND.n17625 GND.n17624 0.003
R17382 GND.n17626 GND.n17625 0.003
R17383 GND.n17627 GND.n17626 0.003
R17384 GND.n17628 GND.n17627 0.003
R17385 GND.n17629 GND.n17628 0.003
R17386 GND.n17630 GND.n17629 0.003
R17387 GND.n17632 GND.n17631 0.003
R17388 GND.n17633 GND.n17632 0.003
R17389 GND.n17634 GND.n17633 0.003
R17390 GND.n17635 GND.n17634 0.003
R17391 GND.n17636 GND.n17635 0.003
R17392 GND.n17637 GND.n17636 0.003
R17393 GND.n17639 GND.n17638 0.003
R17394 GND.n17640 GND.n17639 0.003
R17395 GND.n17641 GND.n17640 0.003
R17396 GND.n17642 GND.n17641 0.003
R17397 GND.n17643 GND.n17642 0.003
R17398 GND.n17644 GND.n17643 0.003
R17399 GND.n17646 GND.n17645 0.003
R17400 GND.n17647 GND.n17646 0.003
R17401 GND.n17648 GND.n17647 0.003
R17402 GND.n17649 GND.n17648 0.003
R17403 GND.n17650 GND.n17649 0.003
R17404 GND.n17651 GND.n17650 0.003
R17405 GND.n17663 GND.n17662 0.003
R17406 GND.n794 GND.n792 0.003
R17407 GND.n705 GND.n704 0.003
R17408 GND.n789 GND.n711 0.003
R17409 GND.n625 GND.n622 0.003
R17410 GND.n621 GND.n620 0.003
R17411 GND.n708 GND.n707 0.003
R17412 GND.n535 GND.n534 0.003
R17413 GND.n447 GND.n446 0.003
R17414 GND.n531 GND.n453 0.003
R17415 GND.n367 GND.n364 0.003
R17416 GND.n363 GND.n362 0.003
R17417 GND.n450 GND.n449 0.003
R17418 GND.n277 GND.n276 0.003
R17419 GND.n189 GND.n188 0.003
R17420 GND.n273 GND.n195 0.003
R17421 GND.n109 GND.n106 0.003
R17422 GND.n105 GND.n104 0.003
R17423 GND.n192 GND.n191 0.003
R17424 GND.n19 GND.n18 0.003
R17425 GND.n6 GND.n5 0.003
R17426 GND.n10 GND.n7 0.003
R17427 GND.n17702 GND.n17701 0.003
R17428 GND.n17704 GND.n17703 0.003
R17429 GND.n3 GND.n2 0.003
R17430 GND.n17697 GND.n17696 0.003
R17431 GND.n17 GND.n16 0.003
R17432 GND.n17694 GND.n17 0.003
R17433 GND.n17694 GND.n17693 0.003
R17434 GND.n17693 GND.n17692 0.003
R17435 GND.n17692 GND.n17691 0.003
R17436 GND.n17690 GND.n17689 0.003
R17437 GND.n17689 GND.n17688 0.003
R17438 GND.n17688 GND.n17687 0.003
R17439 GND.n17687 GND.n17686 0.003
R17440 GND.n17686 GND.n17685 0.003
R17441 GND.n17685 GND.n17684 0.003
R17442 GND.n17683 GND.n17682 0.003
R17443 GND.n17682 GND.n17681 0.003
R17444 GND.n17681 GND.n17680 0.003
R17445 GND.n17680 GND.n17679 0.003
R17446 GND.n17679 GND.n17678 0.003
R17447 GND.n17678 GND.n17677 0.003
R17448 GND.n17676 GND.n17675 0.003
R17449 GND.n17675 GND.n17674 0.003
R17450 GND.n17674 GND.n17673 0.003
R17451 GND.n17673 GND.n17672 0.003
R17452 GND.n17672 GND.n17671 0.003
R17453 GND.n17671 GND.n17670 0.003
R17454 GND.n9566 GND.n1532 0.003
R17455 GND.n16263 GND.n16262 0.003
R17456 GND.n9529 GND.n9528 0.003
R17457 GND.n5321 GND.n5320 0.003
R17458 GND.n5394 GND.n5393 0.003
R17459 GND.n10834 GND.n10833 0.003
R17460 GND.n10836 GND.n10835 0.003
R17461 GND.n10842 GND.n10839 0.003
R17462 GND.n10841 GND.n10840 0.003
R17463 GND.n10835 GND.n10834 0.003
R17464 GND.n10837 GND.n10836 0.003
R17465 GND.n10842 GND.n10841 0.003
R17466 GND.n10839 GND.n10838 0.003
R17467 GND.n12538 GND.n12534 0.003
R17468 GND.n12537 GND.n12536 0.003
R17469 GND.n13798 GND.n10950 0.003
R17470 GND.n13797 GND.n13796 0.003
R17471 GND.n13794 GND.n13793 0.003
R17472 GND.n13792 GND.n13791 0.003
R17473 GND.n13798 GND.n13797 0.003
R17474 GND.n12535 GND.n10950 0.003
R17475 GND.n13793 GND.n13792 0.003
R17476 GND.n13795 GND.n13794 0.003
R17477 GND.n12538 GND.n12537 0.003
R17478 GND.n12534 GND.n12533 0.003
R17479 GND.n11495 GND.n11494 0.003
R17480 GND.n11497 GND.n11496 0.003
R17481 GND.n11503 GND.n11500 0.003
R17482 GND.n11502 GND.n11501 0.003
R17483 GND.n11496 GND.n11495 0.003
R17484 GND.n11498 GND.n11497 0.003
R17485 GND.n11503 GND.n11502 0.003
R17486 GND.n11500 GND.n11499 0.003
R17487 GND.n11031 GND.n11030 0.003
R17488 GND.n11033 GND.n11032 0.003
R17489 GND.n11040 GND.n11035 0.003
R17490 GND.n11039 GND.n11038 0.003
R17491 GND.n11036 GND.n11010 0.003
R17492 GND.n11009 GND.n11008 0.003
R17493 GND.n11040 GND.n11039 0.003
R17494 GND.n11035 GND.n11034 0.003
R17495 GND.n11032 GND.n11031 0.003
R17496 GND.n11030 GND.n11029 0.003
R17497 GND.n11010 GND.n11009 0.003
R17498 GND.n11037 GND.n11036 0.003
R17499 GND.n8235 GND.n5829 0.003
R17500 GND.n8234 GND.n8233 0.003
R17501 GND.n8231 GND.n8230 0.003
R17502 GND.n8229 GND.n8228 0.003
R17503 GND.n8230 GND.n8229 0.003
R17504 GND.n8232 GND.n8231 0.003
R17505 GND.n8235 GND.n8234 0.003
R17506 GND.n5829 GND.n5828 0.003
R17507 GND.n6412 GND.n6345 0.003
R17508 GND.n6411 GND.n6410 0.003
R17509 GND.n6408 GND.n6407 0.003
R17510 GND.n6406 GND.n6405 0.003
R17511 GND.n6403 GND.n6402 0.003
R17512 GND.n6361 GND.n6360 0.003
R17513 GND.n6407 GND.n6406 0.003
R17514 GND.n6409 GND.n6408 0.003
R17515 GND.n6402 GND.n6361 0.003
R17516 GND.n6404 GND.n6403 0.003
R17517 GND.n6345 GND.n6344 0.003
R17518 GND.n6412 GND.n6411 0.003
R17519 GND.n6590 GND.n6582 0.003
R17520 GND.n6589 GND.n6588 0.003
R17521 GND.n6586 GND.n6585 0.003
R17522 GND.n6584 GND.n6583 0.003
R17523 GND.n6585 GND.n6584 0.003
R17524 GND.n6587 GND.n6586 0.003
R17525 GND.n6582 GND.n6581 0.003
R17526 GND.n6590 GND.n6589 0.003
R17527 GND.n7501 GND.n6161 0.003
R17528 GND.n7503 GND.n7502 0.003
R17529 GND.n7506 GND.n7505 0.003
R17530 GND.n7508 GND.n7507 0.003
R17531 GND.n7513 GND.n7510 0.003
R17532 GND.n7512 GND.n7511 0.003
R17533 GND.n7507 GND.n7506 0.003
R17534 GND.n7505 GND.n7504 0.003
R17535 GND.n7502 GND.n7501 0.003
R17536 GND.n6161 GND.n6160 0.003
R17537 GND.n7513 GND.n7512 0.003
R17538 GND.n7510 GND.n7509 0.003
R17539 GND.n9507 GND.n9506 0.003
R17540 GND.n9509 GND.n9508 0.003
R17541 GND.n9517 GND.n9516 0.003
R17542 GND.n9514 GND.n9513 0.003
R17543 GND.n9512 GND.n9511 0.003
R17544 GND.n9513 GND.n9512 0.003
R17545 GND.n9515 GND.n9514 0.003
R17546 GND.n9518 GND.n9517 0.003
R17547 GND.n9508 GND.n9507 0.003
R17548 GND.n9506 GND.n9505 0.003
R17549 GND.n2274 GND.n2273 0.003
R17550 GND.n2387 GND.n2386 0.003
R17551 GND.n2461 GND.n2390 0.003
R17552 GND.n2391 GND.n1927 0.003
R17553 GND.n1926 GND.n1925 0.003
R17554 GND.n2392 GND.n2391 0.003
R17555 GND.n1927 GND.n1926 0.003
R17556 GND.n2390 GND.n2389 0.003
R17557 GND.n2386 GND.n2274 0.003
R17558 GND.n2388 GND.n2387 0.003
R17559 GND.n2846 GND.n2842 0.003
R17560 GND.n2845 GND.n2844 0.003
R17561 GND.n3497 GND.n1943 0.003
R17562 GND.n3493 GND.n3492 0.003
R17563 GND.n3491 GND.n3490 0.003
R17564 GND.n2843 GND.n1943 0.003
R17565 GND.n3492 GND.n3491 0.003
R17566 GND.n3494 GND.n3493 0.003
R17567 GND.n2842 GND.n2841 0.003
R17568 GND.n2846 GND.n2845 0.003
R17569 GND.n14363 GND.n14362 0.003
R17570 GND.n14365 GND.n14364 0.003
R17571 GND.n15456 GND.n14367 0.003
R17572 GND.n15458 GND.n15457 0.003
R17573 GND.n15463 GND.n15460 0.003
R17574 GND.n15462 GND.n15461 0.003
R17575 GND.n15463 GND.n15462 0.003
R17576 GND.n15460 GND.n15459 0.003
R17577 GND.n15457 GND.n15456 0.003
R17578 GND.n14367 GND.n14366 0.003
R17579 GND.n14364 GND.n14363 0.003
R17580 GND.n14362 GND.n14361 0.003
R17581 GND.n14989 GND.n14411 0.003
R17582 GND.n14991 GND.n14990 0.003
R17583 GND.n14994 GND.n14993 0.003
R17584 GND.n14996 GND.n14995 0.003
R17585 GND.n15001 GND.n14998 0.003
R17586 GND.n15000 GND.n14999 0.003
R17587 GND.n14995 GND.n14994 0.003
R17588 GND.n14993 GND.n14992 0.003
R17589 GND.n14990 GND.n14989 0.003
R17590 GND.n14411 GND.n14410 0.003
R17591 GND.n15001 GND.n15000 0.003
R17592 GND.n14998 GND.n14997 0.003
R17593 GND.n16411 GND.n16410 0.003
R17594 GND.n16413 GND.n16412 0.003
R17595 GND.n16569 GND.n16568 0.003
R17596 GND.n16395 GND.n16394 0.003
R17597 GND.n16322 GND.n16321 0.003
R17598 GND.n16394 GND.n16393 0.003
R17599 GND.n16412 GND.n16411 0.003
R17600 GND.n16483 GND.n16413 0.003
R17601 GND.n16568 GND.n16567 0.003
R17602 GND.n16318 GND.n16317 0.003
R17603 GND.n16393 GND.n16322 0.003
R17604 GND.n16672 GND.n16671 0.003
R17605 GND.n16674 GND.n16673 0.003
R17606 GND.n16830 GND.n16829 0.003
R17607 GND.n16656 GND.n16655 0.003
R17608 GND.n16583 GND.n16582 0.003
R17609 GND.n16655 GND.n16654 0.003
R17610 GND.n16673 GND.n16672 0.003
R17611 GND.n16744 GND.n16674 0.003
R17612 GND.n16829 GND.n16828 0.003
R17613 GND.n16579 GND.n16578 0.003
R17614 GND.n16654 GND.n16583 0.003
R17615 GND.n16933 GND.n16932 0.003
R17616 GND.n16935 GND.n16934 0.003
R17617 GND.n17091 GND.n17090 0.003
R17618 GND.n16917 GND.n16916 0.003
R17619 GND.n16844 GND.n16843 0.003
R17620 GND.n16916 GND.n16915 0.003
R17621 GND.n16934 GND.n16933 0.003
R17622 GND.n17005 GND.n16935 0.003
R17623 GND.n17090 GND.n17089 0.003
R17624 GND.n16840 GND.n16839 0.003
R17625 GND.n16915 GND.n16844 0.003
R17626 GND.n17194 GND.n17193 0.003
R17627 GND.n17196 GND.n17195 0.003
R17628 GND.n17352 GND.n17351 0.003
R17629 GND.n17178 GND.n17177 0.003
R17630 GND.n17105 GND.n17104 0.003
R17631 GND.n17177 GND.n17176 0.003
R17632 GND.n17195 GND.n17194 0.003
R17633 GND.n17266 GND.n17196 0.003
R17634 GND.n17351 GND.n17350 0.003
R17635 GND.n17101 GND.n17100 0.003
R17636 GND.n17176 GND.n17105 0.003
R17637 GND.n17455 GND.n17454 0.003
R17638 GND.n17457 GND.n17456 0.003
R17639 GND.n17613 GND.n17612 0.003
R17640 GND.n17439 GND.n17438 0.003
R17641 GND.n17366 GND.n17365 0.003
R17642 GND.n17438 GND.n17437 0.003
R17643 GND.n17456 GND.n17455 0.003
R17644 GND.n17527 GND.n17457 0.003
R17645 GND.n17612 GND.n17611 0.003
R17646 GND.n17362 GND.n17361 0.003
R17647 GND.n17437 GND.n17366 0.003
R17648 GND.n629 GND.n628 0.003
R17649 GND.n681 GND.n680 0.003
R17650 GND.n785 GND.n784 0.003
R17651 GND.n615 GND.n614 0.003
R17652 GND.n543 GND.n542 0.003
R17653 GND.n616 GND.n615 0.003
R17654 GND.n614 GND.n543 0.003
R17655 GND.n702 GND.n681 0.003
R17656 GND.n680 GND.n629 0.003
R17657 GND.n784 GND.n783 0.003
R17658 GND.n539 GND.n538 0.003
R17659 GND.n371 GND.n370 0.003
R17660 GND.n423 GND.n422 0.003
R17661 GND.n527 GND.n526 0.003
R17662 GND.n357 GND.n356 0.003
R17663 GND.n285 GND.n284 0.003
R17664 GND.n358 GND.n357 0.003
R17665 GND.n356 GND.n285 0.003
R17666 GND.n444 GND.n423 0.003
R17667 GND.n422 GND.n371 0.003
R17668 GND.n526 GND.n525 0.003
R17669 GND.n281 GND.n280 0.003
R17670 GND.n113 GND.n112 0.003
R17671 GND.n165 GND.n164 0.003
R17672 GND.n269 GND.n268 0.003
R17673 GND.n99 GND.n98 0.003
R17674 GND.n27 GND.n26 0.003
R17675 GND.n100 GND.n99 0.003
R17676 GND.n98 GND.n27 0.003
R17677 GND.n186 GND.n165 0.003
R17678 GND.n164 GND.n113 0.003
R17679 GND.n268 GND.n267 0.003
R17680 GND.n23 GND.n22 0.003
R17681 GND.n17728 GND.n17727 0.003
R17682 GND.n17780 GND.n17779 0.003
R17683 GND.n17805 GND.n17804 0.003
R17684 GND.n17857 GND.n17856 0.003
R17685 GND.n17934 GND.n17863 0.003
R17686 GND.n17936 GND.n17935 0.003
R17687 GND.n17863 GND.n17862 0.003
R17688 GND.n17935 GND.n17934 0.003
R17689 GND.n17801 GND.n17780 0.003
R17690 GND.n17779 GND.n17728 0.003
R17691 GND.n17856 GND.n17805 0.003
R17692 GND.n17858 GND.n17857 0.003
R17693 GND.n1564 GND.n1563 0.003
R17694 GND.n5289 GND.n5288 0.003
R17695 GND.n5372 GND.n5371 0.003
R17696 GND.n9522 GND.n9521 0.003
R17697 GND.n16250 GND.n16249 0.003
R17698 GND.n9575 GND.n9574 0.003
R17699 GND.n5310 GND.n5309 0.003
R17700 GND.n14495 GND.n14494 0.003
R17701 GND.n17658 GND.n17656 0.002
R17702 GND.n17665 GND.n17664 0.002
R17703 GND.n15453 GND.n15452 0.002
R17704 GND.n14124 GND.n14123 0.002
R17705 GND.n14166 GND.n14165 0.002
R17706 GND.n1678 GND.n1677 0.002
R17707 GND.n1587 GND.n1586 0.002
R17708 GND.n2471 GND.n2470 0.002
R17709 GND.n3161 GND.n2204 0.002
R17710 GND.n2008 GND.n2007 0.002
R17711 GND.n1965 GND.n1964 0.002
R17712 GND.n14668 GND.n14666 0.002
R17713 GND.n14673 GND.n14671 0.002
R17714 GND.n14622 GND.n14620 0.002
R17715 GND.n14617 GND.n14615 0.002
R17716 GND.n10623 GND.n10621 0.002
R17717 GND.n10628 GND.n10626 0.002
R17718 GND.n15486 GND.n15484 0.002
R17719 GND.n15482 GND.n15479 0.002
R17720 GND.n14350 GND.n14348 0.002
R17721 GND.n14345 GND.n14343 0.002
R17722 GND.n14182 GND.n14181 0.002
R17723 GND.n14181 GND.n14180 0.002
R17724 GND.n14179 GND.n14178 0.002
R17725 GND.n14178 GND.n14159 0.002
R17726 GND.n14267 GND.n14265 0.002
R17727 GND.n14263 GND.n14260 0.002
R17728 GND.n14836 GND.n14834 0.002
R17729 GND.n14826 GND.n14817 0.002
R17730 GND.n3572 GND.n3570 0.002
R17731 GND.n3568 GND.n3565 0.002
R17732 GND.n4835 GND.n4833 0.002
R17733 GND.n4840 GND.n4838 0.002
R17734 GND.n6257 GND.n6255 0.002
R17735 GND.n6247 GND.n6239 0.002
R17736 GND.n12624 GND.n12622 0.002
R17737 GND.n12614 GND.n12605 0.002
R17738 GND.n10760 GND.n10758 0.002
R17739 GND.n10755 GND.n10753 0.002
R17740 GND.n13945 GND.n13943 0.002
R17741 GND.n13950 GND.n13948 0.002
R17742 GND.n13822 GND.n13820 0.002
R17743 GND.n13818 GND.n13815 0.002
R17744 GND.n13771 GND.n13769 0.002
R17745 GND.n13776 GND.n13774 0.002
R17746 GND.n11238 GND.n11236 0.002
R17747 GND.n11228 GND.n11220 0.002
R17748 GND.n13645 GND.n13643 0.002
R17749 GND.n13635 GND.n13627 0.002
R17750 GND.n14004 GND.n14001 0.002
R17751 GND.n12758 GND.n12756 0.002
R17752 GND.n12763 GND.n12761 0.002
R17753 GND.n11671 GND.n11669 0.002
R17754 GND.n11676 GND.n11674 0.002
R17755 GND.n11567 GND.n11565 0.002
R17756 GND.n11572 GND.n11570 0.002
R17757 GND.n11064 GND.n11062 0.002
R17758 GND.n11060 GND.n11057 0.002
R17759 GND.n13277 GND.n13275 0.002
R17760 GND.n13273 GND.n13270 0.002
R17761 GND.n11367 GND.n11365 0.002
R17762 GND.n11372 GND.n11370 0.002
R17763 GND.n13420 GND.n13412 0.002
R17764 GND.n13431 GND.n13429 0.002
R17765 GND.n11319 GND.n11318 0.002
R17766 GND.n11956 GND.n11955 0.002
R17767 GND.n11954 GND.n11953 0.002
R17768 GND.n11883 GND.n11882 0.002
R17769 GND.n11881 GND.n11880 0.002
R17770 GND.n12266 GND.n12265 0.002
R17771 GND.n12268 GND.n12267 0.002
R17772 GND.n12339 GND.n12338 0.002
R17773 GND.n12341 GND.n12340 0.002
R17774 GND.n13062 GND.n13061 0.002
R17775 GND.n13060 GND.n13059 0.002
R17776 GND.n12988 GND.n12987 0.002
R17777 GND.n12986 GND.n12985 0.002
R17778 GND.n7754 GND.n7753 0.002
R17779 GND.n7756 GND.n7755 0.002
R17780 GND.n7828 GND.n7827 0.002
R17781 GND.n7830 GND.n7829 0.002
R17782 GND.n8207 GND.n8205 0.002
R17783 GND.n8212 GND.n8210 0.002
R17784 GND.n8296 GND.n8294 0.002
R17785 GND.n8301 GND.n8299 0.002
R17786 GND.n6350 GND.n6348 0.002
R17787 GND.n5857 GND.n5855 0.002
R17788 GND.n5981 GND.n5979 0.002
R17789 GND.n5986 GND.n5984 0.002
R17790 GND.n6463 GND.n6461 0.002
R17791 GND.n6459 GND.n6456 0.002
R17792 GND.n8072 GND.n8070 0.002
R17793 GND.n8061 GND.n8053 0.002
R17794 GND.n6057 GND.n6050 0.002
R17795 GND.n7070 GND.n7062 0.002
R17796 GND.n7081 GND.n7079 0.002
R17797 GND.n6893 GND.n6891 0.002
R17798 GND.n6898 GND.n6896 0.002
R17799 GND.n6658 GND.n6656 0.002
R17800 GND.n6663 GND.n6661 0.002
R17801 GND.n6755 GND.n6753 0.002
R17802 GND.n6760 GND.n6758 0.002
R17803 GND.n7479 GND.n7477 0.002
R17804 GND.n7484 GND.n7482 0.002
R17805 GND.n7397 GND.n7394 0.002
R17806 GND.n7538 GND.n7536 0.002
R17807 GND.n7534 GND.n7531 0.002
R17808 GND.n7299 GND.n7297 0.002
R17809 GND.n7288 GND.n7279 0.002
R17810 GND.n9574 GND.n9573 0.002
R17811 GND.n1552 GND.n1551 0.002
R17812 GND.n1564 GND.n1558 0.002
R17813 GND.n9945 GND.n9586 0.002
R17814 GND.n16250 GND.n803 0.002
R17815 GND.n16277 GND.n16276 0.002
R17816 GND.n16246 GND.n16237 0.002
R17817 GND.n16009 GND.n16008 0.002
R17818 GND.n16015 GND.n16013 0.002
R17819 GND.n16106 GND.n16098 0.002
R17820 GND.n16116 GND.n16114 0.002
R17821 GND.n1061 GND.n1060 0.002
R17822 GND.n1059 GND.n1055 0.002
R17823 GND.n972 GND.n970 0.002
R17824 GND.n962 GND.n953 0.002
R17825 GND.n9709 GND.n9708 0.002
R17826 GND.n9715 GND.n9713 0.002
R17827 GND.n9806 GND.n9798 0.002
R17828 GND.n9816 GND.n9814 0.002
R17829 GND.n1299 GND.n1298 0.002
R17830 GND.n1305 GND.n1303 0.002
R17831 GND.n1396 GND.n1388 0.002
R17832 GND.n1407 GND.n1405 0.002
R17833 GND.n10233 GND.n10231 0.002
R17834 GND.n10222 GND.n10213 0.002
R17835 GND.n8798 GND.n8796 0.002
R17836 GND.n8788 GND.n8780 0.002
R17837 GND.n8503 GND.n8501 0.002
R17838 GND.n8492 GND.n8483 0.002
R17839 GND.n9340 GND.n9338 0.002
R17840 GND.n9345 GND.n9343 0.002
R17841 GND.n1745 GND.n1743 0.002
R17842 GND.n1750 GND.n1748 0.002
R17843 GND.n9523 GND.n9522 0.002
R17844 GND.n9524 GND.n9523 0.002
R17845 GND.n9537 GND.n9536 0.002
R17846 GND.n9472 GND.n9470 0.002
R17847 GND.n9468 GND.n9465 0.002
R17848 GND.n1847 GND.n1845 0.002
R17849 GND.n1852 GND.n1850 0.002
R17850 GND.n1603 GND.n1602 0.002
R17851 GND.n1602 GND.n1601 0.002
R17852 GND.n1600 GND.n1599 0.002
R17853 GND.n1599 GND.n1568 0.002
R17854 GND.n8652 GND.n8650 0.002
R17855 GND.n8648 GND.n8645 0.002
R17856 GND.n10059 GND.n10057 0.002
R17857 GND.n10049 GND.n10041 0.002
R17858 GND.n9289 GND.n9281 0.002
R17859 GND.n5311 GND.n5310 0.002
R17860 GND.n5277 GND.n5276 0.002
R17861 GND.n5289 GND.n5283 0.002
R17862 GND.n9008 GND.n9007 0.002
R17863 GND.n9014 GND.n9012 0.002
R17864 GND.n9105 GND.n9097 0.002
R17865 GND.n9115 GND.n9113 0.002
R17866 GND.n4421 GND.n4420 0.002
R17867 GND.n4419 GND.n4415 0.002
R17868 GND.n4332 GND.n4330 0.002
R17869 GND.n4322 GND.n4313 0.002
R17870 GND.n2538 GND.n2536 0.002
R17871 GND.n2543 GND.n2541 0.002
R17872 GND.n3263 GND.n3255 0.002
R17873 GND.n3273 GND.n3271 0.002
R17874 GND.n3453 GND.n3451 0.002
R17875 GND.n3449 GND.n3446 0.002
R17876 GND.n2449 GND.n2447 0.002
R17877 GND.n2444 GND.n2442 0.002
R17878 GND.n2376 GND.n2374 0.002
R17879 GND.n2381 GND.n2379 0.002
R17880 GND.n5020 GND.n5018 0.002
R17881 GND.n5010 GND.n5001 0.002
R17882 GND.n5147 GND.n5145 0.002
R17883 GND.n5152 GND.n5150 0.002
R17884 GND.n3483 GND.n3482 0.002
R17885 GND.n3482 GND.n3481 0.002
R17886 GND.n3480 GND.n3479 0.002
R17887 GND.n3479 GND.n3478 0.002
R17888 GND.n2110 GND.n2108 0.002
R17889 GND.n2106 GND.n2103 0.002
R17890 GND.n2190 GND.n2188 0.002
R17891 GND.n2185 GND.n2183 0.002
R17892 GND.n2024 GND.n2023 0.002
R17893 GND.n2023 GND.n2022 0.002
R17894 GND.n2021 GND.n2020 0.002
R17895 GND.n2020 GND.n2001 0.002
R17896 GND.n2919 GND.n2917 0.002
R17897 GND.n2915 GND.n2912 0.002
R17898 GND.n4674 GND.n4672 0.002
R17899 GND.n4664 GND.n4655 0.002
R17900 GND.n3063 GND.n3055 0.002
R17901 GND.n3073 GND.n3071 0.002
R17902 GND.n10487 GND.n10479 0.002
R17903 GND.n10497 GND.n10495 0.002
R17904 GND.n15539 GND.n15536 0.002
R17905 GND.n15632 GND.n15624 0.002
R17906 GND.n15643 GND.n15641 0.002
R17907 GND.n15827 GND.n15825 0.002
R17908 GND.n15823 GND.n15820 0.002
R17909 GND.n14533 GND.n14532 0.002
R17910 GND.n14534 GND.n14533 0.002
R17911 GND.n14536 GND.n14535 0.002
R17912 GND.n14537 GND.n14536 0.002
R17913 GND.n15382 GND.n15380 0.002
R17914 GND.n15378 GND.n15375 0.002
R17915 GND.n14968 GND.n14966 0.002
R17916 GND.n14973 GND.n14971 0.002
R17917 GND.n15068 GND.n15066 0.002
R17918 GND.n15064 GND.n15061 0.002
R17919 GND.n15286 GND.n15285 0.002
R17920 GND.n15194 GND.n15186 0.002
R17921 GND.n15204 GND.n15202 0.002
R17922 GND.n3842 GND.n3841 0.002
R17923 GND.n3840 GND.n3836 0.002
R17924 GND.n3753 GND.n3751 0.002
R17925 GND.n3743 GND.n3735 0.002
R17926 GND.n5680 GND.n5679 0.002
R17927 GND.n5678 GND.n5674 0.002
R17928 GND.n5591 GND.n5589 0.002
R17929 GND.n5581 GND.n5572 0.002
R17930 GND.n5428 GND.n5427 0.002
R17931 GND.n5422 GND.n5253 0.002
R17932 GND.n5372 GND.n5367 0.002
R17933 GND.n16571 GND.n16494 0.002
R17934 GND.n16404 GND.n16403 0.002
R17935 GND.n16401 GND.n16400 0.002
R17936 GND.n16832 GND.n16755 0.002
R17937 GND.n16665 GND.n16664 0.002
R17938 GND.n16662 GND.n16661 0.002
R17939 GND.n17093 GND.n17016 0.002
R17940 GND.n16926 GND.n16925 0.002
R17941 GND.n16923 GND.n16922 0.002
R17942 GND.n17354 GND.n17277 0.002
R17943 GND.n17187 GND.n17186 0.002
R17944 GND.n17184 GND.n17183 0.002
R17945 GND.n17615 GND.n17538 0.002
R17946 GND.n17448 GND.n17447 0.002
R17947 GND.n17445 GND.n17444 0.002
R17948 GND.n641 GND.n640 0.002
R17949 GND.n689 GND.n688 0.002
R17950 GND.n743 GND.n742 0.002
R17951 GND.n715 GND.n714 0.002
R17952 GND.n575 GND.n574 0.002
R17953 GND.n565 GND.n563 0.002
R17954 GND.n789 GND.n788 0.002
R17955 GND.n625 GND.n624 0.002
R17956 GND.n622 GND.n621 0.002
R17957 GND.n383 GND.n382 0.002
R17958 GND.n431 GND.n430 0.002
R17959 GND.n485 GND.n484 0.002
R17960 GND.n457 GND.n456 0.002
R17961 GND.n317 GND.n316 0.002
R17962 GND.n307 GND.n305 0.002
R17963 GND.n531 GND.n530 0.002
R17964 GND.n367 GND.n366 0.002
R17965 GND.n364 GND.n363 0.002
R17966 GND.n125 GND.n124 0.002
R17967 GND.n173 GND.n172 0.002
R17968 GND.n227 GND.n226 0.002
R17969 GND.n199 GND.n198 0.002
R17970 GND.n59 GND.n58 0.002
R17971 GND.n49 GND.n47 0.002
R17972 GND.n273 GND.n272 0.002
R17973 GND.n109 GND.n108 0.002
R17974 GND.n106 GND.n105 0.002
R17975 GND.n17740 GND.n17739 0.002
R17976 GND.n17788 GND.n17787 0.002
R17977 GND.n17816 GND.n17815 0.002
R17978 GND.n17709 GND.n17708 0.002
R17979 GND.n17895 GND.n17894 0.002
R17980 GND.n17885 GND.n17883 0.002
R17981 GND.n7 GND.n6 0.002
R17982 GND.n11 GND.n10 0.002
R17983 GND.n13 GND.n12 0.002
R17984 GND.n17701 GND.n14 0.002
R17985 GND.n17703 GND.n17702 0.002
R17986 GND.n5363 GND.n5362 0.002
R17987 GND.n5355 GND.n5354 0.002
R17988 GND.n17667 GND.n17666 0.002
R17989 GND.n17666 GND.n17665 0.002
R17990 GND.n9536 GND.n9535 0.002
R17991 GND.n17664 GND.n17658 0.002
R17992 GND.n16437 GND.n16436 0.001
R17993 GND.n16523 GND.n16522 0.001
R17994 GND.n16346 GND.n16345 0.001
R17995 GND.n16698 GND.n16697 0.001
R17996 GND.n16784 GND.n16783 0.001
R17997 GND.n16607 GND.n16606 0.001
R17998 GND.n16959 GND.n16958 0.001
R17999 GND.n17045 GND.n17044 0.001
R18000 GND.n16868 GND.n16867 0.001
R18001 GND.n17220 GND.n17219 0.001
R18002 GND.n17306 GND.n17305 0.001
R18003 GND.n17129 GND.n17128 0.001
R18004 GND.n17481 GND.n17480 0.001
R18005 GND.n17567 GND.n17566 0.001
R18006 GND.n17390 GND.n17389 0.001
R18007 GND.n797 GND.n796 0.001
R18008 GND.n5362 GND.n5361 0.001
R18009 GND.n5408 GND.n5375 0.001
R18010 GND.n5420 GND.n5418 0.001
R18011 GND.n5324 GND.n5323 0.001
R18012 GND.n5322 GND.n5290 0.001
R18013 GND.n5262 GND.n1566 0.001
R18014 GND.n9547 GND.n9546 0.001
R18015 GND.n9564 GND.n9563 0.001
R18016 GND.n9565 GND.n1565 0.001
R18017 GND.n16253 GND.n16252 0.001
R18018 GND.n16289 GND.n16288 0.001
R18019 GND.n16311 GND.n16310 0.001
R18020 GND.n17665 GND.n16312 0.001
R18021 GND.n5375 GND.n5374 0.001
R18022 GND.n5323 GND.n5322 0.001
R18023 GND.n9565 GND.n9564 0.001
R18024 GND.n16312 GND.n16311 0.001
R18025 GND.n16310 GND.n16309 0.001
R18026 GND.n16272 GND.n16253 0.001
R18027 GND.n16288 GND.n16272 0.001
R18028 GND.n1565 GND.n1556 0.001
R18029 GND.n9545 GND.n1566 0.001
R18030 GND.n9546 GND.n9545 0.001
R18031 GND.n5290 GND.n5281 0.001
R18032 GND.n5361 GND.n5360 0.001
R18033 GND.n5418 GND.n5408 0.001
R18034 GND.n5424 GND.n5423 0.001
R18035 GND.n9577 GND.n9575 0.001
R18036 GND.n16249 GND.n16247 0.001
R18037 GND.n5309 GND.n5308 0.001
R18038 GND.n9521 GND.n9520 0.001
R18039 GND.n5371 GND.n5370 0.001
R18040 GND.n5288 GND.n5285 0.001
R18041 GND.n1563 GND.n1560 0.001
R18042 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_9/DRAIN GND.n14078 0.001
R18043 GND.n14360 GND.n14359 0.001
R18044 GND.n10887 GND.n10879 0.001
R18045 GND.n10898 GND.n10724 0.001
R18046 GND.n10782 GND.n10771 0.001
R18047 GND.n13882 GND.n13881 0.001
R18048 GND.n13518 GND.n13517 0.001
R18049 GND.n13544 GND.n13542 0.001
R18050 GND.n11120 GND.n11112 0.001
R18051 GND.n11139 GND.n11137 0.001
R18052 GND.n8248 GND.n8237 0.001
R18053 GND.n8159 GND.n8158 0.001
R18054 GND.n8381 GND.n8380 0.001
R18055 GND.n6040 GND.n6032 0.001
R18056 GND.n6059 GND.n6057 0.001
R18057 GND.n7430 GND.n7429 0.001
R18058 GND.n7413 GND.n7411 0.001
R18059 GND.n7394 GND.n7386 0.001
R18060 GND.n7197 GND.n7195 0.001
R18061 GND.n7171 GND.n7170 0.001
R18062 GND.n1532 GND.n1531 0.001
R18063 GND.n1553 GND.n1552 0.001
R18064 GND.n9556 GND.n9555 0.001
R18065 GND.n1558 GND.n1557 0.001
R18066 GND.n16262 GND.n16261 0.001
R18067 GND.n16303 GND.n16302 0.001
R18068 GND.n16278 GND.n16277 0.001
R18069 GND.n9530 GND.n9529 0.001
R18070 GND.n9538 GND.n9537 0.001
R18071 GND.n9497 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN 0.001
R18072 GND.n9504 GND.n9503 0.001
R18073 GND.n9519 GND.n9510 0.001
R18074 GND.n1581 GND.n1570 0.001
R18075 GND.n1684 GND.n1683 0.001
R18076 GND.n9249 GND.n9246 0.001
R18077 GND.n9272 GND.n9264 0.001
R18078 GND.n9291 GND.n9289 0.001
R18079 GND.n5272 GND.n5271 0.001
R18080 GND.n5278 GND.n5277 0.001
R18081 GND.n5329 GND.n5328 0.001
R18082 GND.n5283 GND.n5282 0.001
R18083 GND.n3177 GND.n3175 0.001
R18084 GND.n2477 GND.n2476 0.001
R18085 GND.n3376 GND.n3368 0.001
R18086 GND.n3395 GND.n3393 0.001
R18087 GND.n2461 GND.n2460 0.001
R18088 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_12/DRAIN GND.n2239 0.001
R18089 GND.n2459 GND.n2458 0.001
R18090 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_11/DRAIN GND.n1944 0.001
R18091 GND.n2200 GND.n2199 0.001
R18092 GND.n3497 GND.n3496 0.001
R18093 GND.n1954 GND.n1952 0.001
R18094 GND.n4781 GND.n4773 0.001
R18095 GND.n2671 GND.n2669 0.001
R18096 GND.n4920 GND.n4918 0.001
R18097 GND.n14094 GND.n14086 0.001
R18098 GND.n14113 GND.n14111 0.001
R18099 GND.n15752 GND.n15750 0.001
R18100 GND.n15726 GND.n15725 0.001
R18101 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_13/DRAIN GND.n14635
+ 0.001
R18102 GND.n14629 GND.n14409 0.001
R18103 GND.n14489 GND.n14478 0.001
R18104 GND.n15447 GND.n15446 0.001
R18105 GND.n14474 GND.n14472 0.001
R18106 GND.n15305 GND.n15298 0.001
R18107 GND.n5393 GND.n5392 0.001
R18108 GND.n5392 GND.n5391 0.001
R18109 GND.n5389 GND.n5388 0.001
R18110 GND.n16396 GND.n16395 0.001
R18111 GND.n16494 GND.n16493 0.001
R18112 GND.n16403 GND.n16402 0.001
R18113 GND.n16490 GND.n16489 0.001
R18114 GND.n16491 GND.n16490 0.001
R18115 GND.n17648 GND.n16573 0.001
R18116 GND.n17648 GND.n16406 0.001
R18117 GND.n16316 GND.n16315 0.001
R18118 GND.n16315 GND.n16314 0.001
R18119 GND.n16657 GND.n16656 0.001
R18120 GND.n16755 GND.n16754 0.001
R18121 GND.n16664 GND.n16663 0.001
R18122 GND.n16751 GND.n16750 0.001
R18123 GND.n16752 GND.n16751 0.001
R18124 GND.n17641 GND.n16834 0.001
R18125 GND.n17641 GND.n16667 0.001
R18126 GND.n16577 GND.n16576 0.001
R18127 GND.n16576 GND.n16575 0.001
R18128 GND.n16918 GND.n16917 0.001
R18129 GND.n17016 GND.n17015 0.001
R18130 GND.n16925 GND.n16924 0.001
R18131 GND.n17012 GND.n17011 0.001
R18132 GND.n17013 GND.n17012 0.001
R18133 GND.n17634 GND.n17095 0.001
R18134 GND.n17634 GND.n16928 0.001
R18135 GND.n16838 GND.n16837 0.001
R18136 GND.n16837 GND.n16836 0.001
R18137 GND.n17179 GND.n17178 0.001
R18138 GND.n17277 GND.n17276 0.001
R18139 GND.n17186 GND.n17185 0.001
R18140 GND.n17273 GND.n17272 0.001
R18141 GND.n17274 GND.n17273 0.001
R18142 GND.n17627 GND.n17356 0.001
R18143 GND.n17627 GND.n17189 0.001
R18144 GND.n17099 GND.n17098 0.001
R18145 GND.n17098 GND.n17097 0.001
R18146 GND.n17440 GND.n17439 0.001
R18147 GND.n17538 GND.n17537 0.001
R18148 GND.n17447 GND.n17446 0.001
R18149 GND.n17534 GND.n17533 0.001
R18150 GND.n17535 GND.n17534 0.001
R18151 GND.n17620 GND.n17617 0.001
R18152 GND.n17620 GND.n17450 0.001
R18153 GND.n17360 GND.n17359 0.001
R18154 GND.n17359 GND.n17358 0.001
R18155 GND.n617 GND.n616 0.001
R18156 GND.n788 GND.n787 0.001
R18157 GND.n624 GND.n623 0.001
R18158 GND.n709 GND.n708 0.001
R18159 GND.n710 GND.n709 0.001
R18160 GND.n17673 GND.n791 0.001
R18161 GND.n17673 GND.n627 0.001
R18162 GND.n537 GND.n536 0.001
R18163 GND.n536 GND.n535 0.001
R18164 GND.n359 GND.n358 0.001
R18165 GND.n530 GND.n529 0.001
R18166 GND.n366 GND.n365 0.001
R18167 GND.n451 GND.n450 0.001
R18168 GND.n452 GND.n451 0.001
R18169 GND.n17680 GND.n533 0.001
R18170 GND.n17680 GND.n369 0.001
R18171 GND.n279 GND.n278 0.001
R18172 GND.n278 GND.n277 0.001
R18173 GND.n101 GND.n100 0.001
R18174 GND.n272 GND.n271 0.001
R18175 GND.n108 GND.n107 0.001
R18176 GND.n193 GND.n192 0.001
R18177 GND.n194 GND.n193 0.001
R18178 GND.n17687 GND.n275 0.001
R18179 GND.n17687 GND.n111 0.001
R18180 GND.n21 GND.n20 0.001
R18181 GND.n20 GND.n19 0.001
R18182 GND.n17862 GND.n17861 0.001
R18183 GND.n12 GND.n11 0.001
R18184 GND.n14 GND.n13 0.001
R18185 GND.n2 GND.n1 0.001
R18186 GND.n17694 GND.n15 0.001
R18187 GND.n17695 GND.n17694 0.001
R18188 GND.n17699 GND.n17698 0.001
R18189 GND.n17698 GND.n17697 0.001
R18190 GND.n9570 GND.n9566 0.001
R18191 GND.n5321 GND.n5319 0.001
R18192 GND.n5359 GND.n5358 0.001
R18193 GND.n5365 GND.n5364 0.001
R18194 GND.n5373 GND.n5366 0.001
R18195 GND.n5421 GND.n5338 0.001
R18196 GND.n5335 GND.n5324 0.001
R18197 GND.n5281 GND.n5280 0.001
R18198 GND.n5264 GND.n5263 0.001
R18199 GND.n9548 GND.n9547 0.001
R18200 GND.n9563 GND.n9562 0.001
R18201 GND.n1556 GND.n1555 0.001
R18202 GND.n16251 GND.n802 0.001
R18203 GND.n16305 GND.n16289 0.001
R18204 GND.n16308 GND.n16307 0.001
R18205 GND.n5374 GND.n5373 0.001
R18206 GND.n5421 GND.n5420 0.001
R18207 GND.n5394 GND.n5382 0.001
R18208 GND.n5280 GND.n5265 0.001
R18209 GND.n1555 GND.n1541 0.001
R18210 GND.n16309 GND.n16308 0.001
R18211 GND.n16306 GND.n16305 0.001
R18212 GND.n16263 GND.n16260 0.001
R18213 GND.n16252 GND.n16251 0.001
R18214 GND.n9562 GND.n9551 0.001
R18215 GND.n9549 GND.n9548 0.001
R18216 GND.n9528 GND.n9527 0.001
R18217 GND.n5263 GND.n5262 0.001
R18218 GND.n5337 GND.n5335 0.001
R18219 GND.n5364 GND.n5363 0.001
R18220 GND.n5360 GND.n5359 0.001
R18221 GND.n17531 GND.n17530 0.001
R18222 GND.n17270 GND.n17269 0.001
R18223 GND.n17009 GND.n17008 0.001
R18224 GND.n16748 GND.n16747 0.001
R18225 GND.n16487 GND.n16486 0.001
R18226 GND.n5 GND.n4 0.001
R18227 GND.n190 GND.n189 0.001
R18228 GND.n448 GND.n447 0.001
R18229 GND.n706 GND.n705 0.001
R18230 GND.n17655 GND.n17654 0.001
R18231 GND.n1550 GND.n1549 0.001
R18232 GND.n1550 GND.n1548 0.001
R18233 GND.n9570 GND.n9569 0.001
R18234 GND.n1554 GND.n1546 0.001
R18235 GND.n1554 GND.n1544 0.001
R18236 GND.n9561 GND.n9560 0.001
R18237 GND.n16300 GND.n16297 0.001
R18238 GND.n16260 GND.n16259 0.001
R18239 GND.n16304 GND.n16294 0.001
R18240 GND.n16304 GND.n16292 0.001
R18241 GND.n5275 GND.n5274 0.001
R18242 GND.n5275 GND.n5273 0.001
R18243 GND.n5319 GND.n5318 0.001
R18244 GND.n5279 GND.n5270 0.001
R18245 GND.n5279 GND.n5268 0.001
R18246 GND.n5334 GND.n5333 0.001
R18247 GND.n5382 GND.n5380 0.001
R18248 GND.n5390 GND.n5386 0.001
R18249 GND.n5390 GND.n5385 0.001
R18250 GND.n16275 GND.n16274 0.001
R18251 GND.n9571 GND.n9570 0.001
R18252 GND.n9561 GND.n9553 0.001
R18253 GND.n1538 GND.n1537 0.001
R18254 GND.n1537 GND.n1534 0.001
R18255 GND.n16260 GND.n16256 0.001
R18256 GND.n16269 GND.n16266 0.001
R18257 GND.n16270 GND.n16269 0.001
R18258 GND.n16287 GND.n16284 0.001
R18259 GND.n16287 GND.n16281 0.001
R18260 GND.n16301 GND.n16300 0.001
R18261 GND.n9533 GND.n9531 0.001
R18262 GND.n9527 GND.n9526 0.001
R18263 GND.n9541 GND.n9540 0.001
R18264 GND.n5319 GND.n5315 0.001
R18265 GND.n5334 GND.n5326 0.001
R18266 GND.n5259 GND.n5258 0.001
R18267 GND.n5258 GND.n5255 0.001
R18268 GND.n5398 GND.n5397 0.001
R18269 GND.n5382 GND.n5377 0.001
R18270 GND.n5405 GND.n5402 0.001
R18271 GND.n5406 GND.n5405 0.001
R18272 GND.n5417 GND.n5414 0.001
R18273 GND.n5417 GND.n5411 0.001
R18274 GND.n16399 GND.n16398 0.001
R18275 GND.n16660 GND.n16659 0.001
R18276 GND.n16921 GND.n16920 0.001
R18277 GND.n17182 GND.n17181 0.001
R18278 GND.n17443 GND.n17442 0.001
R18279 GND.n620 GND.n619 0.001
R18280 GND.n362 GND.n361 0.001
R18281 GND.n104 GND.n103 0.001
R18282 GND.n17705 GND.n17704 0.001
R18283 VBIAS.n1633 VBIAS.t39 846.712
R18284 VBIAS.n1571 VBIAS.t29 846.712
R18285 VBIAS.n1590 VBIAS.t16 846.712
R18286 VBIAS.n1625 VBIAS.t14 846.712
R18287 VBIAS.n1730 VBIAS.t0 846.712
R18288 VBIAS.n1668 VBIAS.t2 846.712
R18289 VBIAS.n1687 VBIAS.t4 846.712
R18290 VBIAS.n1722 VBIAS.t6 846.712
R18291 VBIAS.n1454 VBIAS.t34 846.712
R18292 VBIAS.n1799 VBIAS.t27 846.712
R18293 VBIAS.n1813 VBIAS.t23 846.712
R18294 VBIAS.n1442 VBIAS.t22 846.712
R18295 VBIAS.n1420 VBIAS.t38 846.712
R18296 VBIAS.n1866 VBIAS.t26 846.712
R18297 VBIAS.n1880 VBIAS.t25 846.712
R18298 VBIAS.n1408 VBIAS.t13 846.712
R18299 VBIAS.n1476 VBIAS.t36 846.712
R18300 VBIAS.n1538 VBIAS.t37 846.712
R18301 VBIAS.n1530 VBIAS.t24 846.712
R18302 VBIAS.n1495 VBIAS.t12 846.712
R18303 VBIAS.n669 VBIAS.t35 846.712
R18304 VBIAS.n621 VBIAS.t28 846.712
R18305 VBIAS.n607 VBIAS.t11 846.712
R18306 VBIAS.n600 VBIAS.t10 846.712
R18307 VBIAS.n770 VBIAS.t30 846.712
R18308 VBIAS.n722 VBIAS.t19 846.712
R18309 VBIAS.n708 VBIAS.t18 846.712
R18310 VBIAS.n701 VBIAS.t15 846.712
R18311 VBIAS.n871 VBIAS.t33 846.712
R18312 VBIAS.n823 VBIAS.t21 846.712
R18313 VBIAS.n809 VBIAS.t20 846.712
R18314 VBIAS.n802 VBIAS.t8 846.712
R18315 VBIAS.n515 VBIAS.t31 846.712
R18316 VBIAS.n570 VBIAS.t32 846.712
R18317 VBIAS.n563 VBIAS.t17 846.712
R18318 VBIAS.n500 VBIAS.t9 846.712
R18319 VBIAS.n1443 VBIAS.n1442 16.434
R18320 VBIAS.n1409 VBIAS.n1408 16.434
R18321 VBIAS.n1626 VBIAS.n1625 16.332
R18322 VBIAS.n1723 VBIAS.n1722 16.332
R18323 VBIAS.n178 VBIAS.n177 16.332
R18324 VBIAS.n1531 VBIAS.n1530 16.332
R18325 VBIAS.n272 VBIAS.n270 16.332
R18326 VBIAS.n368 VBIAS.n366 16.332
R18327 VBIAS.n464 VBIAS.n462 16.332
R18328 VBIAS.n601 VBIAS.n600 16.253
R18329 VBIAS.n702 VBIAS.n701 16.253
R18330 VBIAS.n803 VBIAS.n802 16.253
R18331 VBIAS.n1003 VBIAS.n1002 16.253
R18332 VBIAS.n1203 VBIAS.n1202 16.253
R18333 VBIAS.n1303 VBIAS.n1302 16.253
R18334 VBIAS.n1103 VBIAS.n1101 16.253
R18335 VBIAS.n905 VBIAS.n904 16.253
R18336 VBIAS.n564 VBIAS.n563 16.253
R18337 VBIAS.n1008 VBIAS.n1006 15.887
R18338 VBIAS.n1591 VBIAS.n1590 15.887
R18339 VBIAS.n1108 VBIAS.n1107 15.887
R18340 VBIAS.n1688 VBIAS.n1687 15.887
R18341 VBIAS.n1208 VBIAS.n1206 15.887
R18342 VBIAS.n1814 VBIAS.n1813 15.887
R18343 VBIAS.n1308 VBIAS.n1306 15.887
R18344 VBIAS.n1881 VBIAS.n1880 15.887
R18345 VBIAS.n1496 VBIAS.n1495 15.887
R18346 VBIAS.n910 VBIAS.n909 15.887
R18347 VBIAS.n238 VBIAS.n237 15.887
R18348 VBIAS.n608 VBIAS.n607 15.887
R18349 VBIAS.n334 VBIAS.n333 15.887
R18350 VBIAS.n709 VBIAS.n708 15.887
R18351 VBIAS.n430 VBIAS.n429 15.887
R18352 VBIAS.n810 VBIAS.n809 15.887
R18353 VBIAS.n502 VBIAS.n500 15.887
R18354 VBIAS.n145 VBIAS.n144 15.887
R18355 VBIAS.n1072 VBIAS.n1071 10.328
R18356 VBIAS.n1023 VBIAS.n1022 10.328
R18357 VBIAS.n1635 VBIAS.n1634 10.328
R18358 VBIAS.n1573 VBIAS.n1572 10.328
R18359 VBIAS.n1172 VBIAS.n1171 10.328
R18360 VBIAS.n1123 VBIAS.n1122 10.328
R18361 VBIAS.n1732 VBIAS.n1731 10.328
R18362 VBIAS.n1670 VBIAS.n1669 10.328
R18363 VBIAS.n1272 VBIAS.n1271 10.328
R18364 VBIAS.n1223 VBIAS.n1222 10.328
R18365 VBIAS.n1456 VBIAS.n1455 10.328
R18366 VBIAS.n1801 VBIAS.n1800 10.328
R18367 VBIAS.n1372 VBIAS.n1371 10.328
R18368 VBIAS.n1323 VBIAS.n1322 10.328
R18369 VBIAS.n1422 VBIAS.n1421 10.328
R18370 VBIAS.n1868 VBIAS.n1867 10.328
R18371 VBIAS.n1540 VBIAS.n1539 10.328
R18372 VBIAS.n1478 VBIAS.n1477 10.328
R18373 VBIAS.n974 VBIAS.n973 10.328
R18374 VBIAS.n925 VBIAS.n924 10.328
R18375 VBIAS.n281 VBIAS.n280 10.328
R18376 VBIAS.n225 VBIAS.n224 10.328
R18377 VBIAS.n671 VBIAS.n670 10.328
R18378 VBIAS.n623 VBIAS.n622 10.328
R18379 VBIAS.n377 VBIAS.n376 10.328
R18380 VBIAS.n321 VBIAS.n320 10.328
R18381 VBIAS.n772 VBIAS.n771 10.328
R18382 VBIAS.n724 VBIAS.n723 10.328
R18383 VBIAS.n473 VBIAS.n472 10.328
R18384 VBIAS.n417 VBIAS.n416 10.328
R18385 VBIAS.n873 VBIAS.n872 10.328
R18386 VBIAS.n825 VBIAS.n824 10.328
R18387 VBIAS.n572 VBIAS.n571 10.328
R18388 VBIAS.n517 VBIAS.n516 10.328
R18389 VBIAS.n187 VBIAS.n186 10.328
R18390 VBIAS.n132 VBIAS.n131 10.328
R18391 VBIAS.n66 VBIAS.n65 9.304
R18392 VBIAS.n1920 VBIAS.n1919 9.304
R18393 VBIAS.n1019 VBIAS.n1018 9.3
R18394 VBIAS.n1077 VBIAS.n1076 9.3
R18395 VBIAS.n1079 VBIAS.n1078 9.3
R18396 VBIAS.n1081 VBIAS.n1080 9.3
R18397 VBIAS.n1015 VBIAS.n1014 9.3
R18398 VBIAS.n1017 VBIAS.n1016 9.3
R18399 VBIAS.n1075 VBIAS.n1074 9.3
R18400 VBIAS.n1074 VBIAS.n1073 9.3
R18401 VBIAS.n1026 VBIAS.n1025 9.3
R18402 VBIAS.n1025 VBIAS.n1024 9.3
R18403 VBIAS.n1567 VBIAS.n1566 9.3
R18404 VBIAS.n1640 VBIAS.n1639 9.3
R18405 VBIAS.n1608 VBIAS.n1607 9.3
R18406 VBIAS.n1611 VBIAS.n1610 9.3
R18407 VBIAS.n1642 VBIAS.n1641 9.3
R18408 VBIAS.n1638 VBIAS.n1637 9.3
R18409 VBIAS.n1637 VBIAS.n1636 9.3
R18410 VBIAS.n1569 VBIAS.n1568 9.3
R18411 VBIAS.n1576 VBIAS.n1575 9.3
R18412 VBIAS.n1575 VBIAS.n1574 9.3
R18413 VBIAS.n1117 VBIAS.n1116 9.3
R18414 VBIAS.n1177 VBIAS.n1176 9.3
R18415 VBIAS.n1119 VBIAS.n1118 9.3
R18416 VBIAS.n1115 VBIAS.n1114 9.3
R18417 VBIAS.n1181 VBIAS.n1180 9.3
R18418 VBIAS.n1179 VBIAS.n1178 9.3
R18419 VBIAS.n1126 VBIAS.n1125 9.3
R18420 VBIAS.n1125 VBIAS.n1124 9.3
R18421 VBIAS.n1175 VBIAS.n1174 9.3
R18422 VBIAS.n1174 VBIAS.n1173 9.3
R18423 VBIAS.n1664 VBIAS.n1663 9.3
R18424 VBIAS.n1737 VBIAS.n1736 9.3
R18425 VBIAS.n1705 VBIAS.n1704 9.3
R18426 VBIAS.n1708 VBIAS.n1707 9.3
R18427 VBIAS.n1739 VBIAS.n1738 9.3
R18428 VBIAS.n1735 VBIAS.n1734 9.3
R18429 VBIAS.n1734 VBIAS.n1733 9.3
R18430 VBIAS.n1666 VBIAS.n1665 9.3
R18431 VBIAS.n1673 VBIAS.n1672 9.3
R18432 VBIAS.n1672 VBIAS.n1671 9.3
R18433 VBIAS.n1219 VBIAS.n1218 9.3
R18434 VBIAS.n1277 VBIAS.n1276 9.3
R18435 VBIAS.n1279 VBIAS.n1278 9.3
R18436 VBIAS.n1281 VBIAS.n1280 9.3
R18437 VBIAS.n1215 VBIAS.n1214 9.3
R18438 VBIAS.n1217 VBIAS.n1216 9.3
R18439 VBIAS.n1275 VBIAS.n1274 9.3
R18440 VBIAS.n1274 VBIAS.n1273 9.3
R18441 VBIAS.n1226 VBIAS.n1225 9.3
R18442 VBIAS.n1225 VBIAS.n1224 9.3
R18443 VBIAS.n1808 VBIAS.n1807 9.3
R18444 VBIAS.n1452 VBIAS.n1451 9.3
R18445 VBIAS.n1778 VBIAS.n1777 9.3
R18446 VBIAS.n1776 VBIAS.n1775 9.3
R18447 VBIAS.n1450 VBIAS.n1449 9.3
R18448 VBIAS.n1459 VBIAS.n1458 9.3
R18449 VBIAS.n1458 VBIAS.n1457 9.3
R18450 VBIAS.n1806 VBIAS.n1805 9.3
R18451 VBIAS.n1804 VBIAS.n1803 9.3
R18452 VBIAS.n1803 VBIAS.n1802 9.3
R18453 VBIAS.n1319 VBIAS.n1318 9.3
R18454 VBIAS.n1377 VBIAS.n1376 9.3
R18455 VBIAS.n1379 VBIAS.n1378 9.3
R18456 VBIAS.n1381 VBIAS.n1380 9.3
R18457 VBIAS.n1315 VBIAS.n1314 9.3
R18458 VBIAS.n1317 VBIAS.n1316 9.3
R18459 VBIAS.n1375 VBIAS.n1374 9.3
R18460 VBIAS.n1374 VBIAS.n1373 9.3
R18461 VBIAS.n1326 VBIAS.n1325 9.3
R18462 VBIAS.n1325 VBIAS.n1324 9.3
R18463 VBIAS.n1845 VBIAS.n1844 9.3
R18464 VBIAS.n1843 VBIAS.n1842 9.3
R18465 VBIAS.n1871 VBIAS.n1870 9.3
R18466 VBIAS.n1870 VBIAS.n1869 9.3
R18467 VBIAS.n1875 VBIAS.n1874 9.3
R18468 VBIAS.n1873 VBIAS.n1872 9.3
R18469 VBIAS.n1418 VBIAS.n1417 9.3
R18470 VBIAS.n1416 VBIAS.n1415 9.3
R18471 VBIAS.n1425 VBIAS.n1424 9.3
R18472 VBIAS.n1424 VBIAS.n1423 9.3
R18473 VBIAS.n1472 VBIAS.n1471 9.3
R18474 VBIAS.n1545 VBIAS.n1544 9.3
R18475 VBIAS.n1513 VBIAS.n1512 9.3
R18476 VBIAS.n1547 VBIAS.n1546 9.3
R18477 VBIAS.n1474 VBIAS.n1473 9.3
R18478 VBIAS.n1516 VBIAS.n1515 9.3
R18479 VBIAS.n1543 VBIAS.n1542 9.3
R18480 VBIAS.n1542 VBIAS.n1541 9.3
R18481 VBIAS.n1481 VBIAS.n1480 9.3
R18482 VBIAS.n1480 VBIAS.n1479 9.3
R18483 VBIAS.n979 VBIAS.n978 9.3
R18484 VBIAS.n983 VBIAS.n982 9.3
R18485 VBIAS.n977 VBIAS.n976 9.3
R18486 VBIAS.n976 VBIAS.n975 9.3
R18487 VBIAS.n981 VBIAS.n980 9.3
R18488 VBIAS.n928 VBIAS.n927 9.3
R18489 VBIAS.n927 VBIAS.n926 9.3
R18490 VBIAS.n921 VBIAS.n920 9.3
R18491 VBIAS.n919 VBIAS.n918 9.3
R18492 VBIAS.n917 VBIAS.n916 9.3
R18493 VBIAS.n230 VBIAS.n229 9.3
R18494 VBIAS.n232 VBIAS.n231 9.3
R18495 VBIAS.n286 VBIAS.n285 9.3
R18496 VBIAS.n288 VBIAS.n287 9.3
R18497 VBIAS.n254 VBIAS.n253 9.3
R18498 VBIAS.n284 VBIAS.n283 9.3
R18499 VBIAS.n283 VBIAS.n282 9.3
R18500 VBIAS.n257 VBIAS.n256 9.3
R18501 VBIAS.n228 VBIAS.n227 9.3
R18502 VBIAS.n227 VBIAS.n226 9.3
R18503 VBIAS.n615 VBIAS.n614 9.3
R18504 VBIAS.n617 VBIAS.n616 9.3
R18505 VBIAS.n680 VBIAS.n679 9.3
R18506 VBIAS.n678 VBIAS.n677 9.3
R18507 VBIAS.n676 VBIAS.n675 9.3
R18508 VBIAS.n674 VBIAS.n673 9.3
R18509 VBIAS.n673 VBIAS.n672 9.3
R18510 VBIAS.n619 VBIAS.n618 9.3
R18511 VBIAS.n626 VBIAS.n625 9.3
R18512 VBIAS.n625 VBIAS.n624 9.3
R18513 VBIAS.n326 VBIAS.n325 9.3
R18514 VBIAS.n328 VBIAS.n327 9.3
R18515 VBIAS.n382 VBIAS.n381 9.3
R18516 VBIAS.n384 VBIAS.n383 9.3
R18517 VBIAS.n350 VBIAS.n349 9.3
R18518 VBIAS.n380 VBIAS.n379 9.3
R18519 VBIAS.n379 VBIAS.n378 9.3
R18520 VBIAS.n353 VBIAS.n352 9.3
R18521 VBIAS.n324 VBIAS.n323 9.3
R18522 VBIAS.n323 VBIAS.n322 9.3
R18523 VBIAS.n716 VBIAS.n715 9.3
R18524 VBIAS.n718 VBIAS.n717 9.3
R18525 VBIAS.n781 VBIAS.n780 9.3
R18526 VBIAS.n779 VBIAS.n778 9.3
R18527 VBIAS.n777 VBIAS.n776 9.3
R18528 VBIAS.n775 VBIAS.n774 9.3
R18529 VBIAS.n774 VBIAS.n773 9.3
R18530 VBIAS.n720 VBIAS.n719 9.3
R18531 VBIAS.n727 VBIAS.n726 9.3
R18532 VBIAS.n726 VBIAS.n725 9.3
R18533 VBIAS.n422 VBIAS.n421 9.3
R18534 VBIAS.n424 VBIAS.n423 9.3
R18535 VBIAS.n478 VBIAS.n477 9.3
R18536 VBIAS.n480 VBIAS.n479 9.3
R18537 VBIAS.n446 VBIAS.n445 9.3
R18538 VBIAS.n476 VBIAS.n475 9.3
R18539 VBIAS.n475 VBIAS.n474 9.3
R18540 VBIAS.n449 VBIAS.n448 9.3
R18541 VBIAS.n420 VBIAS.n419 9.3
R18542 VBIAS.n419 VBIAS.n418 9.3
R18543 VBIAS.n817 VBIAS.n816 9.3
R18544 VBIAS.n819 VBIAS.n818 9.3
R18545 VBIAS.n882 VBIAS.n881 9.3
R18546 VBIAS.n880 VBIAS.n879 9.3
R18547 VBIAS.n878 VBIAS.n877 9.3
R18548 VBIAS.n876 VBIAS.n875 9.3
R18549 VBIAS.n875 VBIAS.n874 9.3
R18550 VBIAS.n821 VBIAS.n820 9.3
R18551 VBIAS.n828 VBIAS.n827 9.3
R18552 VBIAS.n827 VBIAS.n826 9.3
R18553 VBIAS.n511 VBIAS.n510 9.3
R18554 VBIAS.n579 VBIAS.n578 9.3
R18555 VBIAS.n581 VBIAS.n580 9.3
R18556 VBIAS.n577 VBIAS.n576 9.3
R18557 VBIAS.n509 VBIAS.n508 9.3
R18558 VBIAS.n513 VBIAS.n512 9.3
R18559 VBIAS.n575 VBIAS.n574 9.3
R18560 VBIAS.n574 VBIAS.n573 9.3
R18561 VBIAS.n520 VBIAS.n519 9.3
R18562 VBIAS.n519 VBIAS.n518 9.3
R18563 VBIAS.n161 VBIAS.n160 9.3
R18564 VBIAS.n194 VBIAS.n193 9.3
R18565 VBIAS.n190 VBIAS.n189 9.3
R18566 VBIAS.n189 VBIAS.n188 9.3
R18567 VBIAS.n192 VBIAS.n191 9.3
R18568 VBIAS.n164 VBIAS.n163 9.3
R18569 VBIAS.n135 VBIAS.n134 9.3
R18570 VBIAS.n134 VBIAS.n133 9.3
R18571 VBIAS.n139 VBIAS.n138 9.3
R18572 VBIAS.n137 VBIAS.n136 9.3
R18573 VBIAS.n1970 VBIAS.n1969 9.3
R18574 VBIAS.n1966 VBIAS.n1965 9.3
R18575 VBIAS.n1948 VBIAS.n1947 9.3
R18576 VBIAS.n1961 VBIAS.n1960 9.3
R18577 VBIAS.n1954 VBIAS.n1953 9.3
R18578 VBIAS.n1917 VBIAS.n1916 9.3
R18579 VBIAS.n9 VBIAS.n8 9.3
R18580 VBIAS.n1935 VBIAS.n1934 9.3
R18581 VBIAS.n1932 VBIAS.n1931 9.3
R18582 VBIAS.n1928 VBIAS.n1927 9.3
R18583 VBIAS.n3 VBIAS.n2 9.3
R18584 VBIAS.n1959 VBIAS.n1958 9.3
R18585 VBIAS.n1972 VBIAS.n1971 9.3
R18586 VBIAS.n63 VBIAS.n62 9.3
R18587 VBIAS.n43 VBIAS.n42 9.3
R18588 VBIAS.n85 VBIAS.n84 9.3
R18589 VBIAS.n79 VBIAS.n78 9.3
R18590 VBIAS.n75 VBIAS.n74 9.3
R18591 VBIAS.n31 VBIAS.n30 9.3
R18592 VBIAS.n28 VBIAS.n27 9.3
R18593 VBIAS.n36 VBIAS.n35 9.3
R18594 VBIAS.n54 VBIAS.n53 9.3
R18595 VBIAS.n52 VBIAS.n51 9.3
R18596 VBIAS.n24 VBIAS.n23 9.3
R18597 VBIAS.n48 VBIAS.n47 9.3
R18598 VBIAS.n41 VBIAS.n40 9.3
R18599 VBIAS.n1029 VBIAS.n1028 9
R18600 VBIAS.n1068 VBIAS.n1067 9
R18601 VBIAS.n1062 VBIAS.n1061 9
R18602 VBIAS.n1055 VBIAS.n1054 9
R18603 VBIAS.n1631 VBIAS.n1630 9
R18604 VBIAS.n1613 VBIAS.n1612 9
R18605 VBIAS.n1606 VBIAS.n1605 9
R18606 VBIAS.n1579 VBIAS.n1578 9
R18607 VBIAS.n1155 VBIAS.n1154 9
R18608 VBIAS.n1129 VBIAS.n1128 9
R18609 VBIAS.n1168 VBIAS.n1167 9
R18610 VBIAS.n1162 VBIAS.n1161 9
R18611 VBIAS.n1728 VBIAS.n1727 9
R18612 VBIAS.n1710 VBIAS.n1709 9
R18613 VBIAS.n1703 VBIAS.n1702 9
R18614 VBIAS.n1676 VBIAS.n1675 9
R18615 VBIAS.n1229 VBIAS.n1228 9
R18616 VBIAS.n1268 VBIAS.n1267 9
R18617 VBIAS.n1262 VBIAS.n1261 9
R18618 VBIAS.n1255 VBIAS.n1254 9
R18619 VBIAS.n1462 VBIAS.n1461 9
R18620 VBIAS.n1772 VBIAS.n1771 9
R18621 VBIAS.n1780 VBIAS.n1779 9
R18622 VBIAS.n1785 VBIAS.n1784 9
R18623 VBIAS.n1329 VBIAS.n1328 9
R18624 VBIAS.n1368 VBIAS.n1367 9
R18625 VBIAS.n1362 VBIAS.n1361 9
R18626 VBIAS.n1355 VBIAS.n1354 9
R18627 VBIAS.n1847 VBIAS.n1846 9
R18628 VBIAS.n1852 VBIAS.n1851 9
R18629 VBIAS.n1428 VBIAS.n1427 9
R18630 VBIAS.n1839 VBIAS.n1838 9
R18631 VBIAS.n1536 VBIAS.n1535 9
R18632 VBIAS.n1518 VBIAS.n1517 9
R18633 VBIAS.n1511 VBIAS.n1510 9
R18634 VBIAS.n1484 VBIAS.n1483 9
R18635 VBIAS.n931 VBIAS.n930 9
R18636 VBIAS.n970 VBIAS.n969 9
R18637 VBIAS.n957 VBIAS.n956 9
R18638 VBIAS.n964 VBIAS.n963 9
R18639 VBIAS.n277 VBIAS.n276 9
R18640 VBIAS.n259 VBIAS.n258 9
R18641 VBIAS.n252 VBIAS.n251 9
R18642 VBIAS.n221 VBIAS.n220 9
R18643 VBIAS.n629 VBIAS.n628 9
R18644 VBIAS.n661 VBIAS.n603 9
R18645 VBIAS.n655 VBIAS.n604 9
R18646 VBIAS.n667 VBIAS.n666 9
R18647 VBIAS.n373 VBIAS.n372 9
R18648 VBIAS.n355 VBIAS.n354 9
R18649 VBIAS.n348 VBIAS.n347 9
R18650 VBIAS.n317 VBIAS.n316 9
R18651 VBIAS.n730 VBIAS.n729 9
R18652 VBIAS.n762 VBIAS.n704 9
R18653 VBIAS.n756 VBIAS.n705 9
R18654 VBIAS.n768 VBIAS.n767 9
R18655 VBIAS.n469 VBIAS.n468 9
R18656 VBIAS.n451 VBIAS.n450 9
R18657 VBIAS.n444 VBIAS.n443 9
R18658 VBIAS.n413 VBIAS.n412 9
R18659 VBIAS.n831 VBIAS.n830 9
R18660 VBIAS.n863 VBIAS.n805 9
R18661 VBIAS.n857 VBIAS.n806 9
R18662 VBIAS.n869 VBIAS.n868 9
R18663 VBIAS.n523 VBIAS.n522 9
R18664 VBIAS.n550 VBIAS.n549 9
R18665 VBIAS.n543 VBIAS.n542 9
R18666 VBIAS.n568 VBIAS.n567 9
R18667 VBIAS.n128 VBIAS.n127 9
R18668 VBIAS.n183 VBIAS.n182 9
R18669 VBIAS.n165 VBIAS.n118 9
R18670 VBIAS.n159 VBIAS.n158 9
R18671 VBIAS.n1946 VBIAS.n1942 9
R18672 VBIAS.n22 VBIAS.n18 9
R18673 VBIAS.n87 VBIAS.n86 9
R18674 VBIAS.n71 VBIAS.n70 9
R18675 VBIAS.n1930 VBIAS.n1925 9
R18676 VBIAS.n11 VBIAS.n10 9
R18677 VBIAS.n1922 VBIAS.n1921 9
R18678 VBIAS.n1956 VBIAS.n1955 9
R18679 VBIAS.n56 VBIAS.n55 9
R18680 VBIAS.n50 VBIAS.n49 9
R18681 VBIAS.n38 VBIAS.n37 9
R18682 VBIAS.n68 VBIAS.n67 9
R18683 VBIAS.n1974 VBIAS.n1973 9
R18684 VBIAS.n1968 VBIAS.n1967 9
R18685 VBIAS.n1059 VBIAS.n1058 8.764
R18686 VBIAS.n1610 VBIAS.n1609 8.764
R18687 VBIAS.n1159 VBIAS.n1158 8.764
R18688 VBIAS.n1707 VBIAS.n1706 8.764
R18689 VBIAS.n1259 VBIAS.n1258 8.764
R18690 VBIAS.n1775 VBIAS.n1774 8.764
R18691 VBIAS.n1359 VBIAS.n1358 8.764
R18692 VBIAS.n1842 VBIAS.n1841 8.764
R18693 VBIAS.n1515 VBIAS.n1514 8.764
R18694 VBIAS.n961 VBIAS.n960 8.764
R18695 VBIAS.n256 VBIAS.n255 8.764
R18696 VBIAS.n659 VBIAS.n657 8.764
R18697 VBIAS.n352 VBIAS.n351 8.764
R18698 VBIAS.n760 VBIAS.n758 8.764
R18699 VBIAS.n448 VBIAS.n447 8.764
R18700 VBIAS.n861 VBIAS.n859 8.764
R18701 VBIAS.n547 VBIAS.n546 8.764
R18702 VBIAS.n163 VBIAS.n162 8.764
R18703 VBIAS.n1071 VBIAS.n1070 6.885
R18704 VBIAS.n1022 VBIAS.n1021 6.885
R18705 VBIAS.n1634 VBIAS.n1633 6.885
R18706 VBIAS.n1572 VBIAS.n1571 6.885
R18707 VBIAS.n1171 VBIAS.n1170 6.885
R18708 VBIAS.n1122 VBIAS.n1121 6.885
R18709 VBIAS.n1731 VBIAS.n1730 6.885
R18710 VBIAS.n1669 VBIAS.n1668 6.885
R18711 VBIAS.n1271 VBIAS.n1270 6.885
R18712 VBIAS.n1222 VBIAS.n1221 6.885
R18713 VBIAS.n1455 VBIAS.n1454 6.885
R18714 VBIAS.n1800 VBIAS.n1799 6.885
R18715 VBIAS.n1371 VBIAS.n1370 6.885
R18716 VBIAS.n1322 VBIAS.n1321 6.885
R18717 VBIAS.n1421 VBIAS.n1420 6.885
R18718 VBIAS.n1867 VBIAS.n1866 6.885
R18719 VBIAS.n1539 VBIAS.n1538 6.885
R18720 VBIAS.n1477 VBIAS.n1476 6.885
R18721 VBIAS.n973 VBIAS.n972 6.885
R18722 VBIAS.n924 VBIAS.n923 6.885
R18723 VBIAS.n280 VBIAS.n279 6.885
R18724 VBIAS.n224 VBIAS.n223 6.885
R18725 VBIAS.n670 VBIAS.n669 6.885
R18726 VBIAS.n622 VBIAS.n621 6.885
R18727 VBIAS.n376 VBIAS.n375 6.885
R18728 VBIAS.n320 VBIAS.n319 6.885
R18729 VBIAS.n771 VBIAS.n770 6.885
R18730 VBIAS.n723 VBIAS.n722 6.885
R18731 VBIAS.n472 VBIAS.n471 6.885
R18732 VBIAS.n416 VBIAS.n415 6.885
R18733 VBIAS.n872 VBIAS.n871 6.885
R18734 VBIAS.n824 VBIAS.n823 6.885
R18735 VBIAS.n571 VBIAS.n570 6.885
R18736 VBIAS.n516 VBIAS.n515 6.885
R18737 VBIAS.n186 VBIAS.n185 6.885
R18738 VBIAS.n131 VBIAS.n130 6.885
R18739 VBIAS.n1008 VBIAS.n1007 6.276
R18740 VBIAS.n1591 VBIAS.n1588 6.276
R18741 VBIAS.n1108 VBIAS.n1105 6.276
R18742 VBIAS.n1688 VBIAS.n1685 6.276
R18743 VBIAS.n1208 VBIAS.n1207 6.276
R18744 VBIAS.n1814 VBIAS.n1811 6.276
R18745 VBIAS.n1308 VBIAS.n1307 6.276
R18746 VBIAS.n1881 VBIAS.n1878 6.276
R18747 VBIAS.n1496 VBIAS.n1493 6.276
R18748 VBIAS.n910 VBIAS.n907 6.276
R18749 VBIAS.n238 VBIAS.n235 6.276
R18750 VBIAS.n608 VBIAS.n605 6.276
R18751 VBIAS.n334 VBIAS.n331 6.276
R18752 VBIAS.n709 VBIAS.n706 6.276
R18753 VBIAS.n430 VBIAS.n427 6.276
R18754 VBIAS.n810 VBIAS.n807 6.276
R18755 VBIAS.n502 VBIAS.n501 6.276
R18756 VBIAS.n145 VBIAS.n142 6.276
R18757 VBIAS.n564 VBIAS.n561 5.776
R18758 VBIAS.n1103 VBIAS.n1102 5.776
R18759 VBIAS.n905 VBIAS.n902 5.776
R18760 VBIAS.n1003 VBIAS.n1000 5.776
R18761 VBIAS.n1203 VBIAS.n1200 5.776
R18762 VBIAS.n1303 VBIAS.n1300 5.776
R18763 VBIAS.n601 VBIAS.n598 5.776
R18764 VBIAS.n702 VBIAS.n699 5.776
R18765 VBIAS.n803 VBIAS.n800 5.776
R18766 VBIAS.n1531 VBIAS.n1528 5.708
R18767 VBIAS.n272 VBIAS.n271 5.708
R18768 VBIAS.n368 VBIAS.n367 5.708
R18769 VBIAS.n464 VBIAS.n463 5.708
R18770 VBIAS.n178 VBIAS.n175 5.708
R18771 VBIAS.n1626 VBIAS.n1623 5.708
R18772 VBIAS.n1723 VBIAS.n1720 5.708
R18773 VBIAS.n1443 VBIAS.n1440 5.531
R18774 VBIAS.n1409 VBIAS.n1406 5.531
R18775 VBIAS.n1060 VBIAS.n1059 4.65
R18776 VBIAS.n1160 VBIAS.n1159 4.65
R18777 VBIAS.n1260 VBIAS.n1259 4.65
R18778 VBIAS.n1360 VBIAS.n1359 4.65
R18779 VBIAS.n962 VBIAS.n961 4.65
R18780 VBIAS.n660 VBIAS.n659 4.65
R18781 VBIAS.n761 VBIAS.n760 4.65
R18782 VBIAS.n862 VBIAS.n861 4.65
R18783 VBIAS.n548 VBIAS.n547 4.65
R18784 VBIAS.n26 VBIAS.n17 4.574
R18785 VBIAS.n1950 VBIAS.n1941 4.574
R18786 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE VBIAS.n1052 4.5
R18787 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE VBIAS.n1152 4.5
R18788 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE VBIAS.n1252 4.5
R18789 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE VBIAS.n1352 4.5
R18790 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE VBIAS.n954 4.5
R18791 VBIAS.n1002 VBIAS.n1001 4.131
R18792 VBIAS.n1006 VBIAS.n1005 4.131
R18793 VBIAS.n1625 VBIAS.n1624 4.131
R18794 VBIAS.n1590 VBIAS.n1589 4.131
R18795 VBIAS.n1101 VBIAS.n1100 4.131
R18796 VBIAS.n1107 VBIAS.n1106 4.131
R18797 VBIAS.n1722 VBIAS.n1721 4.131
R18798 VBIAS.n1687 VBIAS.n1686 4.131
R18799 VBIAS.n1202 VBIAS.n1201 4.131
R18800 VBIAS.n1206 VBIAS.n1205 4.131
R18801 VBIAS.n1442 VBIAS.n1441 4.131
R18802 VBIAS.n1813 VBIAS.n1812 4.131
R18803 VBIAS.n1302 VBIAS.n1301 4.131
R18804 VBIAS.n1306 VBIAS.n1305 4.131
R18805 VBIAS.n1408 VBIAS.n1407 4.131
R18806 VBIAS.n1880 VBIAS.n1879 4.131
R18807 VBIAS.n1530 VBIAS.n1529 4.131
R18808 VBIAS.n1495 VBIAS.n1494 4.131
R18809 VBIAS.n904 VBIAS.n903 4.131
R18810 VBIAS.n909 VBIAS.n908 4.131
R18811 VBIAS.n270 VBIAS.n269 4.131
R18812 VBIAS.n237 VBIAS.n236 4.131
R18813 VBIAS.n600 VBIAS.n599 4.131
R18814 VBIAS.n607 VBIAS.n606 4.131
R18815 VBIAS.n366 VBIAS.n365 4.131
R18816 VBIAS.n333 VBIAS.n332 4.131
R18817 VBIAS.n701 VBIAS.n700 4.131
R18818 VBIAS.n708 VBIAS.n707 4.131
R18819 VBIAS.n462 VBIAS.n461 4.131
R18820 VBIAS.n429 VBIAS.n428 4.131
R18821 VBIAS.n802 VBIAS.n801 4.131
R18822 VBIAS.n809 VBIAS.n808 4.131
R18823 VBIAS.n563 VBIAS.n562 4.131
R18824 VBIAS.n500 VBIAS.n499 4.131
R18825 VBIAS.n177 VBIAS.n176 4.131
R18826 VBIAS.n144 VBIAS.n143 4.131
R18827 VBIAS.n1882 VBIAS.n1881 3.48
R18828 VBIAS.n1815 VBIAS.n1814 3.48
R18829 VBIAS.n953 VBIAS.n932 3.41
R18830 VBIAS.n988 VBIAS.n987 3.41
R18831 VBIAS.n1051 VBIAS.n1030 3.41
R18832 VBIAS.n1086 VBIAS.n1085 3.41
R18833 VBIAS.n1151 VBIAS.n1130 3.41
R18834 VBIAS.n1186 VBIAS.n1185 3.41
R18835 VBIAS.n1251 VBIAS.n1230 3.41
R18836 VBIAS.n1286 VBIAS.n1285 3.41
R18837 VBIAS.n1351 VBIAS.n1330 3.41
R18838 VBIAS.n1386 VBIAS.n1385 3.41
R18839 VBIAS.n854 VBIAS.n853 3.41
R18840 VBIAS.n887 VBIAS.n886 3.41
R18841 VBIAS.n753 VBIAS.n752 3.41
R18842 VBIAS.n786 VBIAS.n785 3.41
R18843 VBIAS.n652 VBIAS.n651 3.41
R18844 VBIAS.n685 VBIAS.n684 3.41
R18845 VBIAS.n554 VBIAS.n553 3.41
R18846 VBIAS.n539 VBIAS.n538 3.41
R18847 VBIAS.n586 VBIAS.n585 3.41
R18848 VBIAS.n1784 VBIAS.n1783 3.388
R18849 VBIAS.n1851 VBIAS.n1850 3.388
R18850 VBIAS.n1941 VBIAS.n1940 3.388
R18851 VBIAS.n17 VBIAS.n16 3.388
R18852 VBIAS.n1592 VBIAS.n1591 3.348
R18853 VBIAS.n1689 VBIAS.n1688 3.348
R18854 VBIAS.n1497 VBIAS.n1496 3.348
R18855 VBIAS.n239 VBIAS.n238 3.348
R18856 VBIAS.n335 VBIAS.n334 3.348
R18857 VBIAS.n431 VBIAS.n430 3.348
R18858 VBIAS.n146 VBIAS.n145 3.348
R18859 VBIAS.n1943 VBIAS.t3 3.326
R18860 VBIAS.n1943 VBIAS.t5 3.326
R18861 VBIAS.n19 VBIAS.t7 3.326
R18862 VBIAS.n19 VBIAS.t1 3.326
R18863 VBIAS.n1028 VBIAS.n1027 3.011
R18864 VBIAS.n1578 VBIAS.n1577 3.011
R18865 VBIAS.n1128 VBIAS.n1127 3.011
R18866 VBIAS.n1675 VBIAS.n1674 3.011
R18867 VBIAS.n1228 VBIAS.n1227 3.011
R18868 VBIAS.n1328 VBIAS.n1327 3.011
R18869 VBIAS.n1483 VBIAS.n1482 3.011
R18870 VBIAS.n930 VBIAS.n929 3.011
R18871 VBIAS.n220 VBIAS.n219 3.011
R18872 VBIAS.n628 VBIAS.n627 3.011
R18873 VBIAS.n316 VBIAS.n315 3.011
R18874 VBIAS.n729 VBIAS.n728 3.011
R18875 VBIAS.n412 VBIAS.n411 3.011
R18876 VBIAS.n830 VBIAS.n829 3.011
R18877 VBIAS.n522 VBIAS.n521 3.011
R18878 VBIAS.n127 VBIAS.n126 3.011
R18879 VBIAS.n1595 VBIAS.n1594 3
R18880 VBIAS.n1646 VBIAS.n1645 3
R18881 VBIAS.n1616 VBIAS.n1615 3
R18882 VBIAS.n1603 VBIAS.n1602 3
R18883 VBIAS.n1692 VBIAS.n1691 3
R18884 VBIAS.n1743 VBIAS.n1742 3
R18885 VBIAS.n1713 VBIAS.n1712 3
R18886 VBIAS.n1700 VBIAS.n1699 3
R18887 VBIAS.n1818 VBIAS.n1817 3
R18888 VBIAS.n1788 VBIAS.n1787 3
R18889 VBIAS.n1885 VBIAS.n1884 3
R18890 VBIAS.n1855 VBIAS.n1854 3
R18891 VBIAS.n1500 VBIAS.n1499 3
R18892 VBIAS.n1551 VBIAS.n1550 3
R18893 VBIAS.n1521 VBIAS.n1520 3
R18894 VBIAS.n1508 VBIAS.n1507 3
R18895 VBIAS.n292 VBIAS.n291 3
R18896 VBIAS.n262 VBIAS.n261 3
R18897 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE VBIAS.n249 3
R18898 VBIAS.n242 VBIAS.n241 3
R18899 VBIAS.n388 VBIAS.n387 3
R18900 VBIAS.n358 VBIAS.n357 3
R18901 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE VBIAS.n345 3
R18902 VBIAS.n338 VBIAS.n337 3
R18903 VBIAS.n484 VBIAS.n483 3
R18904 VBIAS.n454 VBIAS.n453 3
R18905 VBIAS VBIAS.n441 3
R18906 VBIAS.n434 VBIAS.n433 3
R18907 VBIAS.n149 VBIAS.n148 3
R18908 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE VBIAS.n156 3
R18909 VBIAS.n168 VBIAS.n167 3
R18910 VBIAS.n198 VBIAS.n197 3
R18911 VBIAS.n179 VBIAS.n178 2.893
R18912 VBIAS.n1532 VBIAS.n1531 2.893
R18913 VBIAS.n273 VBIAS.n272 2.893
R18914 VBIAS.n369 VBIAS.n368 2.893
R18915 VBIAS.n465 VBIAS.n464 2.893
R18916 VBIAS.n1627 VBIAS.n1626 2.893
R18917 VBIAS.n1724 VBIAS.n1723 2.893
R18918 VBIAS.n1444 VBIAS.n1443 2.796
R18919 VBIAS.n1410 VBIAS.n1409 2.796
R18920 VBIAS.n609 VBIAS.n608 2.747
R18921 VBIAS.n710 VBIAS.n709 2.747
R18922 VBIAS.n811 VBIAS.n810 2.747
R18923 VBIAS.n1009 VBIAS.n1008 2.747
R18924 VBIAS.n1109 VBIAS.n1108 2.747
R18925 VBIAS.n1209 VBIAS.n1208 2.747
R18926 VBIAS.n1309 VBIAS.n1308 2.747
R18927 VBIAS.n503 VBIAS.n502 2.747
R18928 VBIAS.n911 VBIAS.n910 2.746
R18929 VBIAS.n1937 VBIAS.n1936 2.473
R18930 VBIAS.n89 VBIAS.n69 2.469
R18931 VBIAS.n89 VBIAS.n88 2.469
R18932 VBIAS.n1924 VBIAS.n12 2.469
R18933 VBIAS.n1924 VBIAS.n1923 2.469
R18934 VBIAS.n1004 VBIAS.n1003 2.382
R18935 VBIAS.n1204 VBIAS.n1203 2.382
R18936 VBIAS.n1304 VBIAS.n1303 2.382
R18937 VBIAS.n1104 VBIAS.n1103 2.382
R18938 VBIAS.n906 VBIAS.n905 2.382
R18939 VBIAS.n602 VBIAS.n601 2.381
R18940 VBIAS.n703 VBIAS.n702 2.381
R18941 VBIAS.n804 VBIAS.n803 2.381
R18942 VBIAS.n565 VBIAS.n564 2.381
R18943 VBIAS.n1067 VBIAS.n1066 2.258
R18944 VBIAS.n1630 VBIAS.n1629 2.258
R18945 VBIAS.n1167 VBIAS.n1166 2.258
R18946 VBIAS.n1727 VBIAS.n1726 2.258
R18947 VBIAS.n1267 VBIAS.n1266 2.258
R18948 VBIAS.n1367 VBIAS.n1366 2.258
R18949 VBIAS.n1535 VBIAS.n1534 2.258
R18950 VBIAS.n969 VBIAS.n968 2.258
R18951 VBIAS.n276 VBIAS.n275 2.258
R18952 VBIAS.n666 VBIAS.n665 2.258
R18953 VBIAS.n372 VBIAS.n371 2.258
R18954 VBIAS.n767 VBIAS.n766 2.258
R18955 VBIAS.n468 VBIAS.n467 2.258
R18956 VBIAS.n868 VBIAS.n867 2.258
R18957 VBIAS.n567 VBIAS.n566 2.258
R18958 VBIAS.n182 VBIAS.n181 2.258
R18959 VBIAS.n1770 VBIAS.n1769 2.25
R18960 VBIAS.n1837 VBIAS.n1836 2.25
R18961 VBIAS.n58 VBIAS.n57 2.231
R18962 VBIAS.n1976 VBIAS.n1975 2.231
R18963 VBIAS.n1461 VBIAS.n1460 1.882
R18964 VBIAS.n1427 VBIAS.n1426 1.882
R18965 VBIAS.n900 VBIAS.n497 1.713
R18966 VBIAS.n1859 VBIAS.n1858 1.705
R18967 VBIAS.n1834 VBIAS.n1833 1.705
R18968 VBIAS.n1889 VBIAS.n1888 1.705
R18969 VBIAS.n1829 VBIAS.n1828 1.705
R18970 VBIAS.n1822 VBIAS.n1821 1.705
R18971 VBIAS.n1792 VBIAS.n1791 1.705
R18972 VBIAS.n1767 VBIAS.n1766 1.705
R18973 VBIAS.n1762 VBIAS.n1761 1.705
R18974 VBIAS.n1073 VBIAS.n1072 1.377
R18975 VBIAS.n1024 VBIAS.n1023 1.377
R18976 VBIAS.n1636 VBIAS.n1635 1.377
R18977 VBIAS.n1574 VBIAS.n1573 1.377
R18978 VBIAS.n1173 VBIAS.n1172 1.377
R18979 VBIAS.n1124 VBIAS.n1123 1.377
R18980 VBIAS.n1733 VBIAS.n1732 1.377
R18981 VBIAS.n1671 VBIAS.n1670 1.377
R18982 VBIAS.n1273 VBIAS.n1272 1.377
R18983 VBIAS.n1224 VBIAS.n1223 1.377
R18984 VBIAS.n1457 VBIAS.n1456 1.377
R18985 VBIAS.n1802 VBIAS.n1801 1.377
R18986 VBIAS.n1373 VBIAS.n1372 1.377
R18987 VBIAS.n1324 VBIAS.n1323 1.377
R18988 VBIAS.n1423 VBIAS.n1422 1.377
R18989 VBIAS.n1869 VBIAS.n1868 1.377
R18990 VBIAS.n1541 VBIAS.n1540 1.377
R18991 VBIAS.n1479 VBIAS.n1478 1.377
R18992 VBIAS.n975 VBIAS.n974 1.377
R18993 VBIAS.n926 VBIAS.n925 1.377
R18994 VBIAS.n282 VBIAS.n281 1.377
R18995 VBIAS.n226 VBIAS.n225 1.377
R18996 VBIAS.n672 VBIAS.n671 1.377
R18997 VBIAS.n624 VBIAS.n623 1.377
R18998 VBIAS.n378 VBIAS.n377 1.377
R18999 VBIAS.n322 VBIAS.n321 1.377
R19000 VBIAS.n773 VBIAS.n772 1.377
R19001 VBIAS.n725 VBIAS.n724 1.377
R19002 VBIAS.n474 VBIAS.n473 1.377
R19003 VBIAS.n418 VBIAS.n417 1.377
R19004 VBIAS.n874 VBIAS.n873 1.377
R19005 VBIAS.n826 VBIAS.n825 1.377
R19006 VBIAS.n573 VBIAS.n572 1.377
R19007 VBIAS.n518 VBIAS.n517 1.377
R19008 VBIAS.n188 VBIAS.n187 1.377
R19009 VBIAS.n133 VBIAS.n132 1.377
R19010 VBIAS.n20 VBIAS.n19 1.155
R19011 VBIAS.n1944 VBIAS.n1943 1.155
R19012 VBIAS.n1649 VBIAS.n1648 1.137
R19013 VBIAS.n1188 VBIAS.n1187 1.137
R19014 VBIAS.n1746 VBIAS.n1745 1.137
R19015 VBIAS.n1088 VBIAS.n1087 1.137
R19016 VBIAS.n1288 VBIAS.n1287 1.137
R19017 VBIAS.n1388 VBIAS.n1387 1.137
R19018 VBIAS.n687 VBIAS.n686 1.137
R19019 VBIAS.n788 VBIAS.n787 1.137
R19020 VBIAS.n889 VBIAS.n888 1.137
R19021 VBIAS.n295 VBIAS.n294 1.137
R19022 VBIAS.n391 VBIAS.n390 1.137
R19023 VBIAS.n487 VBIAS.n486 1.137
R19024 VBIAS.n1913 VBIAS.n1906 1.137
R19025 VBIAS.n1913 VBIAS.n1912 1.137
R19026 VBIAS.n108 VBIAS.n107 1.137
R19027 VBIAS.n1898 VBIAS.n1897 1.137
R19028 VBIAS.n1399 VBIAS.n1398 0.967
R19029 VBIAS.n900 VBIAS.n899 0.96
R19030 VBIAS.n1891 VBIAS.n1890 0.955
R19031 VBIAS.n21 VBIAS.n20 0.921
R19032 VBIAS.n1945 VBIAS.n1944 0.921
R19033 VBIAS.n1554 VBIAS.n1553 0.897
R19034 VBIAS.n588 VBIAS.n587 0.897
R19035 VBIAS.n990 VBIAS.n989 0.897
R19036 VBIAS.n201 VBIAS.n200 0.897
R19037 VBIAS.n1891 VBIAS.n1399 0.807
R19038 VBIAS.n788 VBIAS.n697 0.787
R19039 VBIAS.n391 VBIAS.n305 0.787
R19040 VBIAS.n1074 VBIAS.n1069 0.752
R19041 VBIAS.n1025 VBIAS.n1020 0.752
R19042 VBIAS.n1637 VBIAS.n1632 0.752
R19043 VBIAS.n1575 VBIAS.n1570 0.752
R19044 VBIAS.n1174 VBIAS.n1169 0.752
R19045 VBIAS.n1125 VBIAS.n1120 0.752
R19046 VBIAS.n1734 VBIAS.n1729 0.752
R19047 VBIAS.n1672 VBIAS.n1667 0.752
R19048 VBIAS.n1274 VBIAS.n1269 0.752
R19049 VBIAS.n1225 VBIAS.n1220 0.752
R19050 VBIAS.n1458 VBIAS.n1453 0.752
R19051 VBIAS.n1803 VBIAS.n1798 0.752
R19052 VBIAS.n1374 VBIAS.n1369 0.752
R19053 VBIAS.n1325 VBIAS.n1320 0.752
R19054 VBIAS.n1424 VBIAS.n1419 0.752
R19055 VBIAS.n1870 VBIAS.n1865 0.752
R19056 VBIAS.n1542 VBIAS.n1537 0.752
R19057 VBIAS.n1480 VBIAS.n1475 0.752
R19058 VBIAS.n976 VBIAS.n971 0.752
R19059 VBIAS.n927 VBIAS.n922 0.752
R19060 VBIAS.n283 VBIAS.n278 0.752
R19061 VBIAS.n227 VBIAS.n222 0.752
R19062 VBIAS.n673 VBIAS.n668 0.752
R19063 VBIAS.n625 VBIAS.n620 0.752
R19064 VBIAS.n379 VBIAS.n374 0.752
R19065 VBIAS.n323 VBIAS.n318 0.752
R19066 VBIAS.n774 VBIAS.n769 0.752
R19067 VBIAS.n726 VBIAS.n721 0.752
R19068 VBIAS.n475 VBIAS.n470 0.752
R19069 VBIAS.n419 VBIAS.n414 0.752
R19070 VBIAS.n875 VBIAS.n870 0.752
R19071 VBIAS.n827 VBIAS.n822 0.752
R19072 VBIAS.n574 VBIAS.n569 0.752
R19073 VBIAS.n519 VBIAS.n514 0.752
R19074 VBIAS.n189 VBIAS.n184 0.752
R19075 VBIAS.n134 VBIAS.n129 0.752
R19076 VBIAS.n1941 VBIAS.n1939 0.506
R19077 VBIAS.n17 VBIAS.n15 0.506
R19078 VBIAS.n1965 VBIAS.n1964 0.476
R19079 VBIAS.n47 VBIAS.n46 0.476
R19080 VBIAS.n1953 VBIAS.n1952 0.445
R19081 VBIAS.n35 VBIAS.n34 0.445
R19082 VBIAS.n1927 VBIAS.n1926 0.414
R19083 VBIAS.n74 VBIAS.n73 0.414
R19084 VBIAS.n8 VBIAS.n7 0.382
R19085 VBIAS.n84 VBIAS.n83 0.382
R19086 VBIAS.n1059 VBIAS.n1057 0.376
R19087 VBIAS.n1159 VBIAS.n1157 0.376
R19088 VBIAS.n1259 VBIAS.n1257 0.376
R19089 VBIAS.n1359 VBIAS.n1357 0.376
R19090 VBIAS.n961 VBIAS.n959 0.376
R19091 VBIAS.n659 VBIAS.n658 0.376
R19092 VBIAS.n760 VBIAS.n759 0.376
R19093 VBIAS.n861 VBIAS.n860 0.376
R19094 VBIAS.n547 VBIAS.n545 0.376
R19095 VBIAS.n1892 VBIAS.n1891 0.341
R19096 VBIAS.n1088 VBIAS.n998 0.302
R19097 VBIAS.n1188 VBIAS.n1098 0.302
R19098 VBIAS.n1288 VBIAS.n1198 0.302
R19099 VBIAS.n1388 VBIAS.n1298 0.302
R19100 VBIAS.n1746 VBIAS.n1659 0.286
R19101 VBIAS.n1649 VBIAS.n1562 0.286
R19102 VBIAS.n889 VBIAS.n798 0.286
R19103 VBIAS.n687 VBIAS.n596 0.286
R19104 VBIAS.n295 VBIAS.n209 0.286
R19105 VBIAS.n487 VBIAS.n401 0.286
R19106 VBIAS.n1893 VBIAS.n1892 0.279
R19107 VBIAS.n1757 VBIAS.n1756 0.278
R19108 VBIAS.n1824 VBIAS.n1823 0.277
R19109 VBIAS.n1914 VBIAS.n1913 0.213
R19110 VBIAS.n1399 VBIAS.n900 0.149
R19111 VBIAS.n1935 VBIAS.n1933 0.06
R19112 VBIAS.n1962 VBIAS.n1961 0.06
R19113 VBIAS.n32 VBIAS.n31 0.06
R19114 VBIAS.n44 VBIAS.n43 0.06
R19115 VBIAS.n1832 VBIAS.n1400 0.056
R19116 VBIAS.n1765 VBIAS.n1434 0.056
R19117 VBIAS.n1751 VBIAS.n1750 0.056
R19118 VBIAS.n1654 VBIAS.n1653 0.056
R19119 VBIAS.n1557 VBIAS.n1556 0.056
R19120 VBIAS.n993 VBIAS.n992 0.056
R19121 VBIAS.n1093 VBIAS.n1092 0.056
R19122 VBIAS.n1193 VBIAS.n1192 0.056
R19123 VBIAS.n1293 VBIAS.n1292 0.056
R19124 VBIAS.n1393 VBIAS.n1392 0.056
R19125 VBIAS.n894 VBIAS.n893 0.056
R19126 VBIAS.n793 VBIAS.n792 0.056
R19127 VBIAS.n692 VBIAS.n691 0.056
R19128 VBIAS.n591 VBIAS.n590 0.056
R19129 VBIAS.n204 VBIAS.n203 0.056
R19130 VBIAS.n300 VBIAS.n299 0.056
R19131 VBIAS.n396 VBIAS.n395 0.056
R19132 VBIAS.n492 VBIAS.n491 0.056
R19133 VBIAS.n57 VBIAS.n26 0.054
R19134 VBIAS.n1975 VBIAS.n1950 0.054
R19135 VBIAS.n1975 VBIAS.n1974 0.054
R19136 VBIAS.n57 VBIAS.n56 0.054
R19137 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/DRAIN VBIAS.n1980
+ 0.054
R19138 VBIAS.n3 VBIAS.n1 0.049
R19139 VBIAS.n79 VBIAS.n77 0.049
R19140 VBIAS.n76 VBIAS.n75 0.048
R19141 VBIAS.n1892 VBIAS 0.048
R19142 VBIAS.n1048 VBIAS.n1047 0.045
R19143 VBIAS.n1598 VBIAS.n1597 0.045
R19144 VBIAS.n1148 VBIAS.n1147 0.045
R19145 VBIAS.n1695 VBIAS.n1694 0.045
R19146 VBIAS.n1248 VBIAS.n1247 0.045
R19147 VBIAS.n1796 VBIAS.n1795 0.045
R19148 VBIAS.n1348 VBIAS.n1347 0.045
R19149 VBIAS.n1863 VBIAS.n1862 0.045
R19150 VBIAS.n1503 VBIAS.n1502 0.045
R19151 VBIAS.n950 VBIAS.n949 0.045
R19152 VBIAS.n245 VBIAS.n244 0.045
R19153 VBIAS.n648 VBIAS.n647 0.045
R19154 VBIAS.n341 VBIAS.n340 0.045
R19155 VBIAS.n749 VBIAS.n748 0.045
R19156 VBIAS.n437 VBIAS.n436 0.045
R19157 VBIAS.n850 VBIAS.n849 0.045
R19158 VBIAS.n535 VBIAS.n534 0.045
R19159 VBIAS.n152 VBIAS.n151 0.045
R19160 VBIAS.n1033 VBIAS.n1032 0.043
R19161 VBIAS.n1621 VBIAS.n1620 0.043
R19162 VBIAS.n1133 VBIAS.n1132 0.043
R19163 VBIAS.n1718 VBIAS.n1717 0.043
R19164 VBIAS.n1233 VBIAS.n1232 0.043
R19165 VBIAS.n1772 VBIAS.n1770 0.043
R19166 VBIAS.n1466 VBIAS.n1465 0.043
R19167 VBIAS.n1333 VBIAS.n1332 0.043
R19168 VBIAS.n1839 VBIAS.n1837 0.043
R19169 VBIAS.n1432 VBIAS.n1431 0.043
R19170 VBIAS.n1526 VBIAS.n1525 0.043
R19171 VBIAS.n935 VBIAS.n934 0.043
R19172 VBIAS.n267 VBIAS.n266 0.043
R19173 VBIAS.n632 VBIAS.n631 0.043
R19174 VBIAS.n363 VBIAS.n362 0.043
R19175 VBIAS.n733 VBIAS.n732 0.043
R19176 VBIAS.n459 VBIAS.n458 0.043
R19177 VBIAS.n834 VBIAS.n833 0.043
R19178 VBIAS.n558 VBIAS.n557 0.043
R19179 VBIAS.n173 VBIAS.n172 0.043
R19180 VBIAS.n1954 VBIAS.n1951 0.043
R19181 VBIAS.n36 VBIAS.n33 0.043
R19182 VBIAS.n1614 VBIAS.n1613 0.041
R19183 VBIAS.n1711 VBIAS.n1710 0.041
R19184 VBIAS.n1861 VBIAS.n1860 0.041
R19185 VBIAS.n1794 VBIAS.n1793 0.041
R19186 VBIAS.n1754 VBIAS.n1753 0.041
R19187 VBIAS.n1657 VBIAS.n1656 0.041
R19188 VBIAS.n1560 VBIAS.n1559 0.041
R19189 VBIAS.n1519 VBIAS.n1518 0.041
R19190 VBIAS.n996 VBIAS.n995 0.041
R19191 VBIAS.n1096 VBIAS.n1095 0.041
R19192 VBIAS.n1196 VBIAS.n1195 0.041
R19193 VBIAS.n1296 VBIAS.n1295 0.041
R19194 VBIAS.n1396 VBIAS.n1395 0.041
R19195 VBIAS.n260 VBIAS.n259 0.041
R19196 VBIAS.n356 VBIAS.n355 0.041
R19197 VBIAS.n452 VBIAS.n451 0.041
R19198 VBIAS.n897 VBIAS.n896 0.041
R19199 VBIAS.n796 VBIAS.n795 0.041
R19200 VBIAS.n695 VBIAS.n694 0.041
R19201 VBIAS.n594 VBIAS.n593 0.041
R19202 VBIAS.n166 VBIAS.n165 0.041
R19203 VBIAS.n207 VBIAS.n206 0.041
R19204 VBIAS.n303 VBIAS.n302 0.041
R19205 VBIAS.n399 VBIAS.n398 0.041
R19206 VBIAS.n495 VBIAS.n494 0.041
R19207 VBIAS.n1831 VBIAS.n1830 0.04
R19208 VBIAS.n1764 VBIAS.n1763 0.04
R19209 VBIAS.n1748 VBIAS.n1747 0.04
R19210 VBIAS.n1651 VBIAS.n1650 0.04
R19211 VBIAS.n1090 VBIAS.n1089 0.04
R19212 VBIAS.n1190 VBIAS.n1189 0.04
R19213 VBIAS.n1290 VBIAS.n1289 0.04
R19214 VBIAS.n1390 VBIAS.n1389 0.04
R19215 VBIAS.n891 VBIAS.n890 0.04
R19216 VBIAS.n790 VBIAS.n789 0.04
R19217 VBIAS.n689 VBIAS.n688 0.04
R19218 VBIAS.n297 VBIAS.n296 0.04
R19219 VBIAS.n393 VBIAS.n392 0.04
R19220 VBIAS.n489 VBIAS.n488 0.04
R19221 VBIAS.n1966 VBIAS.n1963 0.04
R19222 VBIAS.n48 VBIAS.n45 0.04
R19223 VBIAS.n1040 VBIAS.n1039 0.039
R19224 VBIAS.n1582 VBIAS.n1581 0.039
R19225 VBIAS.n1140 VBIAS.n1139 0.039
R19226 VBIAS.n1679 VBIAS.n1678 0.039
R19227 VBIAS.n1240 VBIAS.n1239 0.039
R19228 VBIAS.n1340 VBIAS.n1339 0.039
R19229 VBIAS.n1487 VBIAS.n1486 0.039
R19230 VBIAS.n942 VBIAS.n941 0.039
R19231 VBIAS.n214 VBIAS.n213 0.039
R19232 VBIAS.n639 VBIAS.n638 0.039
R19233 VBIAS.n310 VBIAS.n309 0.039
R19234 VBIAS.n740 VBIAS.n739 0.039
R19235 VBIAS.n406 VBIAS.n405 0.039
R19236 VBIAS.n841 VBIAS.n840 0.039
R19237 VBIAS.n526 VBIAS.n525 0.039
R19238 VBIAS.n121 VBIAS.n120 0.039
R19239 VBIAS.n1437 VBIAS.n1436 0.038
R19240 VBIAS.n1403 VBIAS.n1402 0.038
R19241 VBIAS.n1606 VBIAS.n1604 0.037
R19242 VBIAS.n1703 VBIAS.n1701 0.037
R19243 VBIAS.n1463 VBIAS.n1462 0.037
R19244 VBIAS.n1429 VBIAS.n1428 0.037
R19245 VBIAS.n1511 VBIAS.n1509 0.037
R19246 VBIAS.n252 VBIAS.n250 0.037
R19247 VBIAS.n348 VBIAS.n346 0.037
R19248 VBIAS.n444 VBIAS.n442 0.037
R19249 VBIAS.n159 VBIAS.n157 0.037
R19250 VBIAS.n22 VBIAS.n21 0.036
R19251 VBIAS.n1946 VBIAS.n1945 0.036
R19252 VBIAS.n1580 VBIAS.n1579 0.035
R19253 VBIAS.n1677 VBIAS.n1676 0.035
R19254 VBIAS.n1809 VBIAS.n1808 0.035
R19255 VBIAS.n1876 VBIAS.n1875 0.035
R19256 VBIAS.n1485 VBIAS.n1484 0.035
R19257 VBIAS.n221 VBIAS.n212 0.035
R19258 VBIAS.n317 VBIAS.n308 0.035
R19259 VBIAS.n413 VBIAS.n404 0.035
R19260 VBIAS.n128 VBIAS.n119 0.035
R19261 VBIAS.n1782 VBIAS.n1781 0.034
R19262 VBIAS.n1786 VBIAS.n1785 0.034
R19263 VBIAS.n1849 VBIAS.n1848 0.034
R19264 VBIAS.n1853 VBIAS.n1852 0.034
R19265 VBIAS.n1567 VBIAS.n1565 0.032
R19266 VBIAS.n1664 VBIAS.n1662 0.032
R19267 VBIAS.n1472 VBIAS.n1470 0.032
R19268 VBIAS.n233 VBIAS.n232 0.032
R19269 VBIAS.n329 VBIAS.n328 0.032
R19270 VBIAS.n425 VBIAS.n424 0.032
R19271 VBIAS.n140 VBIAS.n139 0.032
R19272 VBIAS.n1970 VBIAS.n1968 0.031
R19273 VBIAS.n52 VBIAS.n50 0.031
R19274 VBIAS.n1 VBIAS.n0 0.03
R19275 VBIAS.n77 VBIAS.n76 0.03
R19276 VBIAS.n9 VBIAS.n6 0.029
R19277 VBIAS.n85 VBIAS.n82 0.029
R19278 VBIAS.n1039 VBIAS.n1038 0.029
R19279 VBIAS.n1581 VBIAS.n1563 0.029
R19280 VBIAS.n1139 VBIAS.n1138 0.029
R19281 VBIAS.n1678 VBIAS.n1660 0.029
R19282 VBIAS.n1239 VBIAS.n1238 0.029
R19283 VBIAS.n1339 VBIAS.n1338 0.029
R19284 VBIAS.n1486 VBIAS.n1468 0.029
R19285 VBIAS.n941 VBIAS.n940 0.029
R19286 VBIAS.n213 VBIAS.n210 0.029
R19287 VBIAS.n662 VBIAS.n661 0.029
R19288 VBIAS.n638 VBIAS.n637 0.029
R19289 VBIAS.n309 VBIAS.n306 0.029
R19290 VBIAS.n763 VBIAS.n762 0.029
R19291 VBIAS.n739 VBIAS.n738 0.029
R19292 VBIAS.n405 VBIAS.n402 0.029
R19293 VBIAS.n864 VBIAS.n863 0.029
R19294 VBIAS.n840 VBIAS.n839 0.029
R19295 VBIAS.n525 VBIAS.n524 0.029
R19296 VBIAS.n551 VBIAS.n550 0.029
R19297 VBIAS.n120 VBIAS.n116 0.029
R19298 VBIAS.n1063 VBIAS.n1062 0.028
R19299 VBIAS.n1608 VBIAS.n1606 0.028
R19300 VBIAS.n1163 VBIAS.n1162 0.028
R19301 VBIAS.n1705 VBIAS.n1703 0.028
R19302 VBIAS.n1263 VBIAS.n1262 0.028
R19303 VBIAS.n1363 VBIAS.n1362 0.028
R19304 VBIAS.n1513 VBIAS.n1511 0.028
R19305 VBIAS.n965 VBIAS.n964 0.028
R19306 VBIAS.n254 VBIAS.n252 0.028
R19307 VBIAS.n350 VBIAS.n348 0.028
R19308 VBIAS.n446 VBIAS.n444 0.028
R19309 VBIAS.n161 VBIAS.n159 0.028
R19310 VBIAS.n1914 VBIAS.n90 0.027
R19311 VBIAS.n1041 VBIAS.n1040 0.026
R19312 VBIAS.n1055 VBIAS.n1053 0.026
R19313 VBIAS.n1643 VBIAS.n1642 0.026
R19314 VBIAS.n1613 VBIAS.n1611 0.026
R19315 VBIAS.n1583 VBIAS.n1582 0.026
R19316 VBIAS.n1141 VBIAS.n1140 0.026
R19317 VBIAS.n1155 VBIAS.n1153 0.026
R19318 VBIAS.n1740 VBIAS.n1739 0.026
R19319 VBIAS.n1710 VBIAS.n1708 0.026
R19320 VBIAS.n1680 VBIAS.n1679 0.026
R19321 VBIAS.n1241 VBIAS.n1240 0.026
R19322 VBIAS.n1255 VBIAS.n1253 0.026
R19323 VBIAS.n1780 VBIAS.n1778 0.026
R19324 VBIAS.n1341 VBIAS.n1340 0.026
R19325 VBIAS.n1355 VBIAS.n1353 0.026
R19326 VBIAS.n1847 VBIAS.n1845 0.026
R19327 VBIAS.n1488 VBIAS.n1487 0.026
R19328 VBIAS.n1548 VBIAS.n1547 0.026
R19329 VBIAS.n1518 VBIAS.n1516 0.026
R19330 VBIAS.n957 VBIAS.n955 0.026
R19331 VBIAS.n943 VBIAS.n942 0.026
R19332 VBIAS.n215 VBIAS.n214 0.026
R19333 VBIAS.n289 VBIAS.n288 0.026
R19334 VBIAS.n259 VBIAS.n257 0.026
R19335 VBIAS.n655 VBIAS.n654 0.026
R19336 VBIAS.n640 VBIAS.n639 0.026
R19337 VBIAS.n311 VBIAS.n310 0.026
R19338 VBIAS.n385 VBIAS.n384 0.026
R19339 VBIAS.n355 VBIAS.n353 0.026
R19340 VBIAS.n756 VBIAS.n755 0.026
R19341 VBIAS.n741 VBIAS.n740 0.026
R19342 VBIAS.n407 VBIAS.n406 0.026
R19343 VBIAS.n481 VBIAS.n480 0.026
R19344 VBIAS.n451 VBIAS.n449 0.026
R19345 VBIAS.n857 VBIAS.n856 0.026
R19346 VBIAS.n842 VBIAS.n841 0.026
R19347 VBIAS.n527 VBIAS.n526 0.026
R19348 VBIAS.n543 VBIAS.n541 0.026
R19349 VBIAS.n195 VBIAS.n194 0.026
R19350 VBIAS.n165 VBIAS.n164 0.026
R19351 VBIAS.n122 VBIAS.n121 0.026
R19352 VBIAS.n1932 VBIAS.n1930 0.026
R19353 VBIAS.n1959 VBIAS.n1957 0.026
R19354 VBIAS.n41 VBIAS.n39 0.026
R19355 VBIAS.n667 VBIAS.n664 0.025
R19356 VBIAS.n652 VBIAS.n629 0.025
R19357 VBIAS.n768 VBIAS.n765 0.025
R19358 VBIAS.n753 VBIAS.n730 0.025
R19359 VBIAS.n869 VBIAS.n866 0.025
R19360 VBIAS.n854 VBIAS.n831 0.025
R19361 VBIAS.n539 VBIAS.n523 0.025
R19362 VBIAS.n1068 VBIAS.n1065 0.024
R19363 VBIAS.n1030 VBIAS.n1029 0.024
R19364 VBIAS.n1168 VBIAS.n1165 0.024
R19365 VBIAS.n1130 VBIAS.n1129 0.024
R19366 VBIAS.n1268 VBIAS.n1265 0.024
R19367 VBIAS.n1230 VBIAS.n1229 0.024
R19368 VBIAS.n1817 VBIAS.n1810 0.024
R19369 VBIAS.n1368 VBIAS.n1365 0.024
R19370 VBIAS.n1330 VBIAS.n1329 0.024
R19371 VBIAS.n1884 VBIAS.n1877 0.024
R19372 VBIAS.n970 VBIAS.n967 0.024
R19373 VBIAS.n932 VBIAS.n931 0.024
R19374 VBIAS.n1917 VBIAS.n1915 0.024
R19375 VBIAS.n63 VBIAS.n61 0.024
R19376 VBIAS.n1439 VBIAS.n1438 0.023
R19377 VBIAS.n1405 VBIAS.n1404 0.023
R19378 VBIAS.n6 VBIAS.n5 0.022
R19379 VBIAS.n82 VBIAS.n81 0.022
R19380 VBIAS.n1015 VBIAS.n1013 0.022
R19381 VBIAS.n1594 VBIAS.n1587 0.022
R19382 VBIAS.n1115 VBIAS.n1113 0.022
R19383 VBIAS.n1691 VBIAS.n1684 0.022
R19384 VBIAS.n1215 VBIAS.n1213 0.022
R19385 VBIAS.n1450 VBIAS.n1448 0.022
R19386 VBIAS.n1452 VBIAS.n1450 0.022
R19387 VBIAS.n1462 VBIAS.n1459 0.022
R19388 VBIAS.n1776 VBIAS.n1773 0.022
R19389 VBIAS.n1315 VBIAS.n1313 0.022
R19390 VBIAS.n1416 VBIAS.n1414 0.022
R19391 VBIAS.n1418 VBIAS.n1416 0.022
R19392 VBIAS.n1428 VBIAS.n1425 0.022
R19393 VBIAS.n1843 VBIAS.n1840 0.022
R19394 VBIAS.n1499 VBIAS.n1492 0.022
R19395 VBIAS.n917 VBIAS.n915 0.022
R19396 VBIAS.n241 VBIAS.n234 0.022
R19397 VBIAS.n615 VBIAS.n613 0.022
R19398 VBIAS.n337 VBIAS.n330 0.022
R19399 VBIAS.n716 VBIAS.n714 0.022
R19400 VBIAS.n433 VBIAS.n426 0.022
R19401 VBIAS.n817 VBIAS.n815 0.022
R19402 VBIAS.n509 VBIAS.n507 0.022
R19403 VBIAS.n148 VBIAS.n141 0.022
R19404 VBIAS.n1767 VBIAS.n1467 0.021
R19405 VBIAS.n1834 VBIAS.n1433 0.021
R19406 VBIAS.n1950 VBIAS.n1949 0.021
R19407 VBIAS.n26 VBIAS.n25 0.021
R19408 VBIAS.n1642 VBIAS.n1640 0.02
R19409 VBIAS.n1638 VBIAS.n1631 0.02
R19410 VBIAS.n1739 VBIAS.n1737 0.02
R19411 VBIAS.n1735 VBIAS.n1728 0.02
R19412 VBIAS.n1547 VBIAS.n1545 0.02
R19413 VBIAS.n1543 VBIAS.n1536 0.02
R19414 VBIAS.n288 VBIAS.n286 0.02
R19415 VBIAS.n284 VBIAS.n277 0.02
R19416 VBIAS.n384 VBIAS.n382 0.02
R19417 VBIAS.n380 VBIAS.n373 0.02
R19418 VBIAS.n480 VBIAS.n478 0.02
R19419 VBIAS.n476 VBIAS.n469 0.02
R19420 VBIAS.n194 VBIAS.n192 0.02
R19421 VBIAS.n190 VBIAS.n183 0.02
R19422 VBIAS.n1035 VBIAS.n1034 0.019
R19423 VBIAS.n1050 VBIAS.n1049 0.019
R19424 VBIAS.n1056 VBIAS.n1055 0.019
R19425 VBIAS.n1619 VBIAS.n1618 0.019
R19426 VBIAS.n1600 VBIAS.n1599 0.019
R19427 VBIAS.n1135 VBIAS.n1134 0.019
R19428 VBIAS.n1150 VBIAS.n1149 0.019
R19429 VBIAS.n1156 VBIAS.n1155 0.019
R19430 VBIAS.n1716 VBIAS.n1715 0.019
R19431 VBIAS.n1697 VBIAS.n1696 0.019
R19432 VBIAS.n1235 VBIAS.n1234 0.019
R19433 VBIAS.n1250 VBIAS.n1249 0.019
R19434 VBIAS.n1256 VBIAS.n1255 0.019
R19435 VBIAS.n1335 VBIAS.n1334 0.019
R19436 VBIAS.n1350 VBIAS.n1349 0.019
R19437 VBIAS.n1356 VBIAS.n1355 0.019
R19438 VBIAS.n1524 VBIAS.n1523 0.019
R19439 VBIAS.n1505 VBIAS.n1504 0.019
R19440 VBIAS.n958 VBIAS.n957 0.019
R19441 VBIAS.n937 VBIAS.n936 0.019
R19442 VBIAS.n952 VBIAS.n951 0.019
R19443 VBIAS.n265 VBIAS.n264 0.019
R19444 VBIAS.n247 VBIAS.n246 0.019
R19445 VBIAS.n656 VBIAS.n655 0.019
R19446 VBIAS.n634 VBIAS.n633 0.019
R19447 VBIAS.n650 VBIAS.n649 0.019
R19448 VBIAS.n361 VBIAS.n360 0.019
R19449 VBIAS.n343 VBIAS.n342 0.019
R19450 VBIAS.n757 VBIAS.n756 0.019
R19451 VBIAS.n735 VBIAS.n734 0.019
R19452 VBIAS.n751 VBIAS.n750 0.019
R19453 VBIAS.n457 VBIAS.n456 0.019
R19454 VBIAS.n439 VBIAS.n438 0.019
R19455 VBIAS.n858 VBIAS.n857 0.019
R19456 VBIAS.n836 VBIAS.n835 0.019
R19457 VBIAS.n852 VBIAS.n851 0.019
R19458 VBIAS.n556 VBIAS.n555 0.019
R19459 VBIAS.n537 VBIAS.n536 0.019
R19460 VBIAS.n544 VBIAS.n543 0.019
R19461 VBIAS.n171 VBIAS.n170 0.019
R19462 VBIAS.n154 VBIAS.n153 0.019
R19463 VBIAS.n1974 VBIAS.n1972 0.019
R19464 VBIAS.n1949 VBIAS.n1948 0.019
R19465 VBIAS.n56 VBIAS.n54 0.019
R19466 VBIAS.n25 VBIAS.n24 0.019
R19467 VBIAS.n1082 VBIAS.n1081 0.018
R19468 VBIAS.n1062 VBIAS.n1060 0.018
R19469 VBIAS.n1645 VBIAS.n1644 0.018
R19470 VBIAS.n1593 VBIAS.n1592 0.018
R19471 VBIAS.n1182 VBIAS.n1181 0.018
R19472 VBIAS.n1162 VBIAS.n1160 0.018
R19473 VBIAS.n1742 VBIAS.n1741 0.018
R19474 VBIAS.n1690 VBIAS.n1689 0.018
R19475 VBIAS.n1282 VBIAS.n1281 0.018
R19476 VBIAS.n1262 VBIAS.n1260 0.018
R19477 VBIAS.n1445 VBIAS.n1444 0.018
R19478 VBIAS.n1448 VBIAS.n1447 0.018
R19479 VBIAS.n1791 VBIAS.n1790 0.018
R19480 VBIAS.n1382 VBIAS.n1381 0.018
R19481 VBIAS.n1362 VBIAS.n1360 0.018
R19482 VBIAS.n1411 VBIAS.n1410 0.018
R19483 VBIAS.n1414 VBIAS.n1413 0.018
R19484 VBIAS.n1858 VBIAS.n1857 0.018
R19485 VBIAS.n1550 VBIAS.n1549 0.018
R19486 VBIAS.n1498 VBIAS.n1497 0.018
R19487 VBIAS.n984 VBIAS.n983 0.018
R19488 VBIAS.n964 VBIAS.n962 0.018
R19489 VBIAS.n291 VBIAS.n290 0.018
R19490 VBIAS.n234 VBIAS.n233 0.018
R19491 VBIAS.n240 VBIAS.n239 0.018
R19492 VBIAS.n681 VBIAS.n680 0.018
R19493 VBIAS.n661 VBIAS.n660 0.018
R19494 VBIAS.n387 VBIAS.n386 0.018
R19495 VBIAS.n330 VBIAS.n329 0.018
R19496 VBIAS.n336 VBIAS.n335 0.018
R19497 VBIAS.n782 VBIAS.n781 0.018
R19498 VBIAS.n762 VBIAS.n761 0.018
R19499 VBIAS.n483 VBIAS.n482 0.018
R19500 VBIAS.n426 VBIAS.n425 0.018
R19501 VBIAS.n432 VBIAS.n431 0.018
R19502 VBIAS.n883 VBIAS.n882 0.018
R19503 VBIAS.n863 VBIAS.n862 0.018
R19504 VBIAS.n582 VBIAS.n581 0.018
R19505 VBIAS.n550 VBIAS.n548 0.018
R19506 VBIAS.n197 VBIAS.n196 0.018
R19507 VBIAS.n141 VBIAS.n140 0.018
R19508 VBIAS.n147 VBIAS.n146 0.018
R19509 VBIAS.n12 VBIAS.n11 0.018
R19510 VBIAS.n69 VBIAS.n68 0.018
R19511 VBIAS.n88 VBIAS.n87 0.018
R19512 VBIAS.n1923 VBIAS.n1922 0.018
R19513 VBIAS.n1628 VBIAS.n1627 0.017
R19514 VBIAS.n1644 VBIAS.n1643 0.017
R19515 VBIAS.n1579 VBIAS.n1576 0.017
R19516 VBIAS.n1569 VBIAS.n1567 0.017
R19517 VBIAS.n1725 VBIAS.n1724 0.017
R19518 VBIAS.n1741 VBIAS.n1740 0.017
R19519 VBIAS.n1676 VBIAS.n1673 0.017
R19520 VBIAS.n1666 VBIAS.n1664 0.017
R19521 VBIAS.n1447 VBIAS.n1446 0.017
R19522 VBIAS.n1806 VBIAS.n1804 0.017
R19523 VBIAS.n1810 VBIAS.n1809 0.017
R19524 VBIAS.n1818 VBIAS.n1797 0.017
R19525 VBIAS.n1413 VBIAS.n1412 0.017
R19526 VBIAS.n1873 VBIAS.n1871 0.017
R19527 VBIAS.n1877 VBIAS.n1876 0.017
R19528 VBIAS.n1885 VBIAS.n1864 0.017
R19529 VBIAS.n1533 VBIAS.n1532 0.017
R19530 VBIAS.n1549 VBIAS.n1548 0.017
R19531 VBIAS.n1484 VBIAS.n1481 0.017
R19532 VBIAS.n1474 VBIAS.n1472 0.017
R19533 VBIAS.n274 VBIAS.n273 0.017
R19534 VBIAS.n290 VBIAS.n289 0.017
R19535 VBIAS.n228 VBIAS.n221 0.017
R19536 VBIAS.n232 VBIAS.n230 0.017
R19537 VBIAS.n370 VBIAS.n369 0.017
R19538 VBIAS.n386 VBIAS.n385 0.017
R19539 VBIAS.n324 VBIAS.n317 0.017
R19540 VBIAS.n328 VBIAS.n326 0.017
R19541 VBIAS.n466 VBIAS.n465 0.017
R19542 VBIAS.n482 VBIAS.n481 0.017
R19543 VBIAS.n420 VBIAS.n413 0.017
R19544 VBIAS.n424 VBIAS.n422 0.017
R19545 VBIAS.n180 VBIAS.n179 0.017
R19546 VBIAS.n196 VBIAS.n195 0.017
R19547 VBIAS.n135 VBIAS.n128 0.017
R19548 VBIAS.n139 VBIAS.n137 0.017
R19549 VBIAS.n1816 VBIAS.n1815 0.016
R19550 VBIAS.n1883 VBIAS.n1882 0.016
R19551 VBIAS.n1833 VBIAS.n1831 0.016
R19552 VBIAS.n1860 VBIAS.n1859 0.016
R19553 VBIAS.n1766 VBIAS.n1764 0.016
R19554 VBIAS.n1793 VBIAS.n1792 0.016
R19555 VBIAS.n1749 VBIAS.n1748 0.016
R19556 VBIAS.n1753 VBIAS.n1752 0.016
R19557 VBIAS.n1652 VBIAS.n1651 0.016
R19558 VBIAS.n1656 VBIAS.n1655 0.016
R19559 VBIAS.n1555 VBIAS.n1554 0.016
R19560 VBIAS.n1559 VBIAS.n1558 0.016
R19561 VBIAS.n991 VBIAS.n990 0.016
R19562 VBIAS.n995 VBIAS.n994 0.016
R19563 VBIAS.n1091 VBIAS.n1090 0.016
R19564 VBIAS.n1095 VBIAS.n1094 0.016
R19565 VBIAS.n1191 VBIAS.n1190 0.016
R19566 VBIAS.n1195 VBIAS.n1194 0.016
R19567 VBIAS.n1291 VBIAS.n1290 0.016
R19568 VBIAS.n1295 VBIAS.n1294 0.016
R19569 VBIAS.n1391 VBIAS.n1390 0.016
R19570 VBIAS.n1395 VBIAS.n1394 0.016
R19571 VBIAS.n892 VBIAS.n891 0.016
R19572 VBIAS.n896 VBIAS.n895 0.016
R19573 VBIAS.n791 VBIAS.n790 0.016
R19574 VBIAS.n795 VBIAS.n794 0.016
R19575 VBIAS.n690 VBIAS.n689 0.016
R19576 VBIAS.n694 VBIAS.n693 0.016
R19577 VBIAS.n589 VBIAS.n588 0.016
R19578 VBIAS.n593 VBIAS.n592 0.016
R19579 VBIAS.n202 VBIAS.n201 0.016
R19580 VBIAS.n206 VBIAS.n205 0.016
R19581 VBIAS.n298 VBIAS.n297 0.016
R19582 VBIAS.n302 VBIAS.n301 0.016
R19583 VBIAS.n394 VBIAS.n393 0.016
R19584 VBIAS.n398 VBIAS.n397 0.016
R19585 VBIAS.n490 VBIAS.n489 0.016
R19586 VBIAS.n494 VBIAS.n493 0.016
R19587 VBIAS.n1963 VBIAS.n1962 0.016
R19588 VBIAS.n45 VBIAS.n44 0.016
R19589 VBIAS.n1046 VBIAS.n1045 0.015
R19590 VBIAS.n1012 VBIAS.n1011 0.015
R19591 VBIAS.n1576 VBIAS.n1569 0.015
R19592 VBIAS.n1596 VBIAS.n1595 0.015
R19593 VBIAS.n1146 VBIAS.n1145 0.015
R19594 VBIAS.n1112 VBIAS.n1111 0.015
R19595 VBIAS.n1673 VBIAS.n1666 0.015
R19596 VBIAS.n1693 VBIAS.n1692 0.015
R19597 VBIAS.n1246 VBIAS.n1245 0.015
R19598 VBIAS.n1212 VBIAS.n1211 0.015
R19599 VBIAS.n1808 VBIAS.n1806 0.015
R19600 VBIAS.n1346 VBIAS.n1345 0.015
R19601 VBIAS.n1312 VBIAS.n1311 0.015
R19602 VBIAS.n1875 VBIAS.n1873 0.015
R19603 VBIAS.n1890 VBIAS.n1889 0.015
R19604 VBIAS.n1823 VBIAS.n1822 0.015
R19605 VBIAS.n1756 VBIAS.n1755 0.015
R19606 VBIAS.n1659 VBIAS.n1658 0.015
R19607 VBIAS.n1562 VBIAS.n1561 0.015
R19608 VBIAS.n1501 VBIAS.n1500 0.015
R19609 VBIAS.n1481 VBIAS.n1474 0.015
R19610 VBIAS.n914 VBIAS.n913 0.015
R19611 VBIAS.n948 VBIAS.n947 0.015
R19612 VBIAS.n998 VBIAS.n997 0.015
R19613 VBIAS.n1098 VBIAS.n1097 0.015
R19614 VBIAS.n1198 VBIAS.n1197 0.015
R19615 VBIAS.n1298 VBIAS.n1297 0.015
R19616 VBIAS.n1398 VBIAS.n1397 0.015
R19617 VBIAS.n243 VBIAS.n242 0.015
R19618 VBIAS.n230 VBIAS.n228 0.015
R19619 VBIAS.n612 VBIAS.n611 0.015
R19620 VBIAS.n646 VBIAS.n645 0.015
R19621 VBIAS.n339 VBIAS.n338 0.015
R19622 VBIAS.n326 VBIAS.n324 0.015
R19623 VBIAS.n713 VBIAS.n712 0.015
R19624 VBIAS.n747 VBIAS.n746 0.015
R19625 VBIAS.n435 VBIAS.n434 0.015
R19626 VBIAS.n422 VBIAS.n420 0.015
R19627 VBIAS.n814 VBIAS.n813 0.015
R19628 VBIAS.n848 VBIAS.n847 0.015
R19629 VBIAS.n899 VBIAS.n898 0.015
R19630 VBIAS.n798 VBIAS.n797 0.015
R19631 VBIAS.n697 VBIAS.n696 0.015
R19632 VBIAS.n596 VBIAS.n595 0.015
R19633 VBIAS.n533 VBIAS.n532 0.015
R19634 VBIAS.n506 VBIAS.n505 0.015
R19635 VBIAS.n137 VBIAS.n135 0.015
R19636 VBIAS.n150 VBIAS.n149 0.015
R19637 VBIAS.n209 VBIAS.n208 0.015
R19638 VBIAS.n305 VBIAS.n304 0.015
R19639 VBIAS.n401 VBIAS.n400 0.015
R19640 VBIAS.n497 VBIAS.n496 0.015
R19641 VBIAS.n1081 VBIAS.n1079 0.014
R19642 VBIAS.n1075 VBIAS.n1068 0.014
R19643 VBIAS.n1181 VBIAS.n1179 0.014
R19644 VBIAS.n1175 VBIAS.n1168 0.014
R19645 VBIAS.n1281 VBIAS.n1279 0.014
R19646 VBIAS.n1275 VBIAS.n1268 0.014
R19647 VBIAS.n1381 VBIAS.n1379 0.014
R19648 VBIAS.n1375 VBIAS.n1368 0.014
R19649 VBIAS.n983 VBIAS.n981 0.014
R19650 VBIAS.n977 VBIAS.n970 0.014
R19651 VBIAS.n680 VBIAS.n678 0.014
R19652 VBIAS.n674 VBIAS.n667 0.014
R19653 VBIAS.n781 VBIAS.n779 0.014
R19654 VBIAS.n775 VBIAS.n768 0.014
R19655 VBIAS.n882 VBIAS.n880 0.014
R19656 VBIAS.n876 VBIAS.n869 0.014
R19657 VBIAS.n581 VBIAS.n579 0.014
R19658 VBIAS.n575 VBIAS.n568 0.014
R19659 VBIAS.n11 VBIAS.n9 0.014
R19660 VBIAS.n1948 VBIAS.n1946 0.014
R19661 VBIAS.n87 VBIAS.n85 0.014
R19662 VBIAS.n24 VBIAS.n22 0.014
R19663 VBIAS.n1031 VBIAS.n999 0.013
R19664 VBIAS.n1047 VBIAS.n1046 0.013
R19665 VBIAS.n1084 VBIAS.n1083 0.013
R19666 VBIAS.n1013 VBIAS.n1012 0.013
R19667 VBIAS.n1010 VBIAS.n1009 0.013
R19668 VBIAS.n1645 VBIAS.n1628 0.013
R19669 VBIAS.n1646 VBIAS.n1622 0.013
R19670 VBIAS.n1597 VBIAS.n1596 0.013
R19671 VBIAS.n1131 VBIAS.n1099 0.013
R19672 VBIAS.n1147 VBIAS.n1146 0.013
R19673 VBIAS.n1184 VBIAS.n1183 0.013
R19674 VBIAS.n1113 VBIAS.n1112 0.013
R19675 VBIAS.n1110 VBIAS.n1109 0.013
R19676 VBIAS.n1742 VBIAS.n1725 0.013
R19677 VBIAS.n1743 VBIAS.n1719 0.013
R19678 VBIAS.n1694 VBIAS.n1693 0.013
R19679 VBIAS.n1231 VBIAS.n1199 0.013
R19680 VBIAS.n1247 VBIAS.n1246 0.013
R19681 VBIAS.n1284 VBIAS.n1283 0.013
R19682 VBIAS.n1213 VBIAS.n1212 0.013
R19683 VBIAS.n1210 VBIAS.n1209 0.013
R19684 VBIAS.n1446 VBIAS.n1445 0.013
R19685 VBIAS.n1465 VBIAS.n1464 0.013
R19686 VBIAS.n1331 VBIAS.n1299 0.013
R19687 VBIAS.n1347 VBIAS.n1346 0.013
R19688 VBIAS.n1384 VBIAS.n1383 0.013
R19689 VBIAS.n1313 VBIAS.n1312 0.013
R19690 VBIAS.n1310 VBIAS.n1309 0.013
R19691 VBIAS.n1412 VBIAS.n1411 0.013
R19692 VBIAS.n1431 VBIAS.n1430 0.013
R19693 VBIAS.n1829 VBIAS.n1824 0.013
R19694 VBIAS.n1762 VBIAS.n1757 0.013
R19695 VBIAS.n1551 VBIAS.n1527 0.013
R19696 VBIAS.n1502 VBIAS.n1501 0.013
R19697 VBIAS.n1550 VBIAS.n1533 0.013
R19698 VBIAS.n986 VBIAS.n985 0.013
R19699 VBIAS.n915 VBIAS.n914 0.013
R19700 VBIAS.n912 VBIAS.n911 0.013
R19701 VBIAS.n933 VBIAS.n901 0.013
R19702 VBIAS.n949 VBIAS.n948 0.013
R19703 VBIAS.n292 VBIAS.n268 0.013
R19704 VBIAS.n244 VBIAS.n243 0.013
R19705 VBIAS.n291 VBIAS.n274 0.013
R19706 VBIAS.n683 VBIAS.n682 0.013
R19707 VBIAS.n613 VBIAS.n612 0.013
R19708 VBIAS.n610 VBIAS.n609 0.013
R19709 VBIAS.n630 VBIAS.n597 0.013
R19710 VBIAS.n647 VBIAS.n646 0.013
R19711 VBIAS.n388 VBIAS.n364 0.013
R19712 VBIAS.n340 VBIAS.n339 0.013
R19713 VBIAS.n387 VBIAS.n370 0.013
R19714 VBIAS.n784 VBIAS.n783 0.013
R19715 VBIAS.n714 VBIAS.n713 0.013
R19716 VBIAS.n711 VBIAS.n710 0.013
R19717 VBIAS.n731 VBIAS.n698 0.013
R19718 VBIAS.n748 VBIAS.n747 0.013
R19719 VBIAS.n484 VBIAS.n460 0.013
R19720 VBIAS.n436 VBIAS.n435 0.013
R19721 VBIAS.n483 VBIAS.n466 0.013
R19722 VBIAS.n885 VBIAS.n884 0.013
R19723 VBIAS.n815 VBIAS.n814 0.013
R19724 VBIAS.n812 VBIAS.n811 0.013
R19725 VBIAS.n832 VBIAS.n799 0.013
R19726 VBIAS.n849 VBIAS.n848 0.013
R19727 VBIAS.n560 VBIAS.n559 0.013
R19728 VBIAS.n534 VBIAS.n533 0.013
R19729 VBIAS.n584 VBIAS.n583 0.013
R19730 VBIAS.n507 VBIAS.n506 0.013
R19731 VBIAS.n504 VBIAS.n503 0.013
R19732 VBIAS.n197 VBIAS.n180 0.013
R19733 VBIAS.n198 VBIAS.n174 0.013
R19734 VBIAS.n151 VBIAS.n150 0.013
R19735 VBIAS.n1936 VBIAS.n1935 0.012
R19736 VBIAS.n31 VBIAS.n29 0.012
R19737 VBIAS.n1087 VBIAS.n1086 0.011
R19738 VBIAS.n1032 VBIAS.n1031 0.011
R19739 VBIAS.n1034 VBIAS.n1033 0.011
R19740 VBIAS.n1049 VBIAS.n1048 0.011
R19741 VBIAS.n1085 VBIAS.n1004 0.011
R19742 VBIAS.n1083 VBIAS.n1082 0.011
R19743 VBIAS.n1029 VBIAS.n1026 0.011
R19744 VBIAS.n1017 VBIAS.n1015 0.011
R19745 VBIAS.n1640 VBIAS.n1638 0.011
R19746 VBIAS.n1648 VBIAS.n1647 0.011
R19747 VBIAS.n1622 VBIAS.n1621 0.011
R19748 VBIAS.n1620 VBIAS.n1619 0.011
R19749 VBIAS.n1599 VBIAS.n1598 0.011
R19750 VBIAS.n1187 VBIAS.n1186 0.011
R19751 VBIAS.n1132 VBIAS.n1131 0.011
R19752 VBIAS.n1134 VBIAS.n1133 0.011
R19753 VBIAS.n1149 VBIAS.n1148 0.011
R19754 VBIAS.n1185 VBIAS.n1104 0.011
R19755 VBIAS.n1183 VBIAS.n1182 0.011
R19756 VBIAS.n1129 VBIAS.n1126 0.011
R19757 VBIAS.n1117 VBIAS.n1115 0.011
R19758 VBIAS.n1737 VBIAS.n1735 0.011
R19759 VBIAS.n1745 VBIAS.n1744 0.011
R19760 VBIAS.n1719 VBIAS.n1718 0.011
R19761 VBIAS.n1717 VBIAS.n1716 0.011
R19762 VBIAS.n1696 VBIAS.n1695 0.011
R19763 VBIAS.n1287 VBIAS.n1286 0.011
R19764 VBIAS.n1232 VBIAS.n1231 0.011
R19765 VBIAS.n1234 VBIAS.n1233 0.011
R19766 VBIAS.n1249 VBIAS.n1248 0.011
R19767 VBIAS.n1285 VBIAS.n1204 0.011
R19768 VBIAS.n1283 VBIAS.n1282 0.011
R19769 VBIAS.n1229 VBIAS.n1226 0.011
R19770 VBIAS.n1217 VBIAS.n1215 0.011
R19771 VBIAS.n1761 VBIAS.n1760 0.011
R19772 VBIAS.n1797 VBIAS.n1796 0.011
R19773 VBIAS.n1387 VBIAS.n1386 0.011
R19774 VBIAS.n1332 VBIAS.n1331 0.011
R19775 VBIAS.n1334 VBIAS.n1333 0.011
R19776 VBIAS.n1349 VBIAS.n1348 0.011
R19777 VBIAS.n1385 VBIAS.n1304 0.011
R19778 VBIAS.n1383 VBIAS.n1382 0.011
R19779 VBIAS.n1329 VBIAS.n1326 0.011
R19780 VBIAS.n1317 VBIAS.n1315 0.011
R19781 VBIAS.n1828 VBIAS.n1827 0.011
R19782 VBIAS.n1864 VBIAS.n1863 0.011
R19783 VBIAS.n1527 VBIAS.n1526 0.011
R19784 VBIAS.n1525 VBIAS.n1524 0.011
R19785 VBIAS.n1504 VBIAS.n1503 0.011
R19786 VBIAS.n1545 VBIAS.n1543 0.011
R19787 VBIAS.n987 VBIAS.n906 0.011
R19788 VBIAS.n985 VBIAS.n984 0.011
R19789 VBIAS.n931 VBIAS.n928 0.011
R19790 VBIAS.n919 VBIAS.n917 0.011
R19791 VBIAS.n934 VBIAS.n933 0.011
R19792 VBIAS.n936 VBIAS.n935 0.011
R19793 VBIAS.n951 VBIAS.n950 0.011
R19794 VBIAS.n294 VBIAS.n293 0.011
R19795 VBIAS.n268 VBIAS.n267 0.011
R19796 VBIAS.n266 VBIAS.n265 0.011
R19797 VBIAS.n246 VBIAS.n245 0.011
R19798 VBIAS.n286 VBIAS.n284 0.011
R19799 VBIAS.n684 VBIAS.n602 0.011
R19800 VBIAS.n682 VBIAS.n681 0.011
R19801 VBIAS.n629 VBIAS.n626 0.011
R19802 VBIAS.n617 VBIAS.n615 0.011
R19803 VBIAS.n686 VBIAS.n685 0.011
R19804 VBIAS.n631 VBIAS.n630 0.011
R19805 VBIAS.n633 VBIAS.n632 0.011
R19806 VBIAS.n649 VBIAS.n648 0.011
R19807 VBIAS.n390 VBIAS.n389 0.011
R19808 VBIAS.n364 VBIAS.n363 0.011
R19809 VBIAS.n362 VBIAS.n361 0.011
R19810 VBIAS.n342 VBIAS.n341 0.011
R19811 VBIAS.n382 VBIAS.n380 0.011
R19812 VBIAS.n785 VBIAS.n703 0.011
R19813 VBIAS.n783 VBIAS.n782 0.011
R19814 VBIAS.n730 VBIAS.n727 0.011
R19815 VBIAS.n718 VBIAS.n716 0.011
R19816 VBIAS.n787 VBIAS.n786 0.011
R19817 VBIAS.n732 VBIAS.n731 0.011
R19818 VBIAS.n734 VBIAS.n733 0.011
R19819 VBIAS.n750 VBIAS.n749 0.011
R19820 VBIAS.n486 VBIAS.n485 0.011
R19821 VBIAS.n460 VBIAS.n459 0.011
R19822 VBIAS.n458 VBIAS.n457 0.011
R19823 VBIAS.n438 VBIAS.n437 0.011
R19824 VBIAS.n478 VBIAS.n476 0.011
R19825 VBIAS.n886 VBIAS.n804 0.011
R19826 VBIAS.n884 VBIAS.n883 0.011
R19827 VBIAS.n831 VBIAS.n828 0.011
R19828 VBIAS.n819 VBIAS.n817 0.011
R19829 VBIAS.n888 VBIAS.n887 0.011
R19830 VBIAS.n833 VBIAS.n832 0.011
R19831 VBIAS.n835 VBIAS.n834 0.011
R19832 VBIAS.n851 VBIAS.n850 0.011
R19833 VBIAS.n559 VBIAS.n558 0.011
R19834 VBIAS.n557 VBIAS.n556 0.011
R19835 VBIAS.n536 VBIAS.n535 0.011
R19836 VBIAS.n585 VBIAS.n565 0.011
R19837 VBIAS.n583 VBIAS.n582 0.011
R19838 VBIAS.n523 VBIAS.n520 0.011
R19839 VBIAS.n511 VBIAS.n509 0.011
R19840 VBIAS.n192 VBIAS.n190 0.011
R19841 VBIAS.n174 VBIAS.n173 0.011
R19842 VBIAS.n172 VBIAS.n171 0.011
R19843 VBIAS.n153 VBIAS.n152 0.011
R19844 VBIAS.n1929 VBIAS.n1928 0.011
R19845 VBIAS.n75 VBIAS.n72 0.011
R19846 VBIAS.n1747 VBIAS.n1746 0.011
R19847 VBIAS.n1650 VBIAS.n1649 0.011
R19848 VBIAS.n1089 VBIAS.n1088 0.011
R19849 VBIAS.n1189 VBIAS.n1188 0.011
R19850 VBIAS.n1289 VBIAS.n1288 0.011
R19851 VBIAS.n1389 VBIAS.n1388 0.011
R19852 VBIAS.n890 VBIAS.n889 0.011
R19853 VBIAS.n789 VBIAS.n788 0.011
R19854 VBIAS.n688 VBIAS.n687 0.011
R19855 VBIAS.n296 VBIAS.n295 0.011
R19856 VBIAS.n392 VBIAS.n391 0.011
R19857 VBIAS.n488 VBIAS.n487 0.011
R19858 VBIAS.n1467 VBIAS.n1466 0.01
R19859 VBIAS.n1433 VBIAS.n1432 0.01
R19860 VBIAS.n90 VBIAS.n89 0.01
R19861 VBIAS.n1086 VBIAS.n999 0.009
R19862 VBIAS.n1085 VBIAS.n1084 0.009
R19863 VBIAS.n1647 VBIAS.n1646 0.009
R19864 VBIAS.n1186 VBIAS.n1099 0.009
R19865 VBIAS.n1185 VBIAS.n1184 0.009
R19866 VBIAS.n1744 VBIAS.n1743 0.009
R19867 VBIAS.n1286 VBIAS.n1199 0.009
R19868 VBIAS.n1285 VBIAS.n1284 0.009
R19869 VBIAS.n1459 VBIAS.n1452 0.009
R19870 VBIAS.n1760 VBIAS.n1759 0.009
R19871 VBIAS.n1386 VBIAS.n1299 0.009
R19872 VBIAS.n1385 VBIAS.n1384 0.009
R19873 VBIAS.n1425 VBIAS.n1418 0.009
R19874 VBIAS.n1827 VBIAS.n1826 0.009
R19875 VBIAS.n1552 VBIAS.n1551 0.009
R19876 VBIAS.n987 VBIAS.n986 0.009
R19877 VBIAS.n988 VBIAS.n901 0.009
R19878 VBIAS.n293 VBIAS.n292 0.009
R19879 VBIAS.n684 VBIAS.n683 0.009
R19880 VBIAS.n685 VBIAS.n597 0.009
R19881 VBIAS.n389 VBIAS.n388 0.009
R19882 VBIAS.n785 VBIAS.n784 0.009
R19883 VBIAS.n786 VBIAS.n698 0.009
R19884 VBIAS.n485 VBIAS.n484 0.009
R19885 VBIAS.n886 VBIAS.n885 0.009
R19886 VBIAS.n887 VBIAS.n799 0.009
R19887 VBIAS.n586 VBIAS.n560 0.009
R19888 VBIAS.n585 VBIAS.n584 0.009
R19889 VBIAS.n199 VBIAS.n198 0.009
R19890 VBIAS.n1956 VBIAS.n1954 0.009
R19891 VBIAS.n1961 VBIAS.n1959 0.009
R19892 VBIAS.n33 VBIAS.n32 0.009
R19893 VBIAS.n38 VBIAS.n36 0.009
R19894 VBIAS.n43 VBIAS.n41 0.009
R19895 VBIAS.n989 VBIAS.n988 0.009
R19896 VBIAS.n200 VBIAS.n199 0.009
R19897 VBIAS.n1553 VBIAS.n1552 0.009
R19898 VBIAS.n587 VBIAS.n586 0.009
R19899 VBIAS.n1924 VBIAS.n1914 0.007
R19900 VBIAS.n1923 VBIAS.n1918 0.007
R19901 VBIAS.n69 VBIAS.n64 0.007
R19902 VBIAS.n12 VBIAS.n4 0.007
R19903 VBIAS.n88 VBIAS.n80 0.007
R19904 VBIAS.n1044 VBIAS.n1043 0.007
R19905 VBIAS.n1019 VBIAS.n1017 0.007
R19906 VBIAS.n1594 VBIAS.n1593 0.007
R19907 VBIAS.n1586 VBIAS.n1585 0.007
R19908 VBIAS.n1144 VBIAS.n1143 0.007
R19909 VBIAS.n1119 VBIAS.n1117 0.007
R19910 VBIAS.n1691 VBIAS.n1690 0.007
R19911 VBIAS.n1683 VBIAS.n1682 0.007
R19912 VBIAS.n1244 VBIAS.n1243 0.007
R19913 VBIAS.n1219 VBIAS.n1217 0.007
R19914 VBIAS.n1817 VBIAS.n1816 0.007
R19915 VBIAS.n1788 VBIAS.n1439 0.007
R19916 VBIAS.n1821 VBIAS.n1819 0.007
R19917 VBIAS.n1344 VBIAS.n1343 0.007
R19918 VBIAS.n1319 VBIAS.n1317 0.007
R19919 VBIAS.n1884 VBIAS.n1883 0.007
R19920 VBIAS.n1855 VBIAS.n1405 0.007
R19921 VBIAS.n1888 VBIAS.n1886 0.007
R19922 VBIAS.n1491 VBIAS.n1490 0.007
R19923 VBIAS.n1499 VBIAS.n1498 0.007
R19924 VBIAS.n921 VBIAS.n919 0.007
R19925 VBIAS.n946 VBIAS.n945 0.007
R19926 VBIAS.n218 VBIAS.n217 0.007
R19927 VBIAS.n250 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE 0.007
R19928 VBIAS.n241 VBIAS.n240 0.007
R19929 VBIAS.n619 VBIAS.n617 0.007
R19930 VBIAS.n644 VBIAS.n643 0.007
R19931 VBIAS.n314 VBIAS.n313 0.007
R19932 VBIAS.n346 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE 0.007
R19933 VBIAS.n337 VBIAS.n336 0.007
R19934 VBIAS.n720 VBIAS.n718 0.007
R19935 VBIAS.n745 VBIAS.n744 0.007
R19936 VBIAS.n410 VBIAS.n409 0.007
R19937 VBIAS.n442 VBIAS 0.007
R19938 VBIAS.n433 VBIAS.n432 0.007
R19939 VBIAS.n821 VBIAS.n819 0.007
R19940 VBIAS.n846 VBIAS.n845 0.007
R19941 VBIAS.n531 VBIAS.n530 0.007
R19942 VBIAS.n513 VBIAS.n511 0.007
R19943 VBIAS.n157 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE 0.007
R19944 VBIAS.n148 VBIAS.n147 0.007
R19945 VBIAS.n125 VBIAS.n124 0.007
R19946 VBIAS.n1918 VBIAS.n1917 0.007
R19947 VBIAS.n64 VBIAS.n63 0.007
R19948 VBIAS.n68 VBIAS.n66 0.006
R19949 VBIAS.n1922 VBIAS.n1920 0.006
R19950 VBIAS.n1830 VBIAS.n1829 0.006
R19951 VBIAS.n1763 VBIAS.n1762 0.006
R19952 VBIAS.n1036 VBIAS.n1035 0.005
R19953 VBIAS.n1052 VBIAS.n1041 0.005
R19954 VBIAS.n1051 VBIAS.n1050 0.005
R19955 VBIAS.n1045 VBIAS.n1044 0.005
R19956 VBIAS.n1043 VBIAS.n1042 0.005
R19957 VBIAS.n1079 VBIAS.n1077 0.005
R19958 VBIAS.n1053 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE 0.005
R19959 VBIAS.n1011 VBIAS.n1010 0.005
R19960 VBIAS.n1604 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE 0.005
R19961 VBIAS.n1618 VBIAS.n1617 0.005
R19962 VBIAS.n1602 VBIAS.n1583 0.005
R19963 VBIAS.n1601 VBIAS.n1600 0.005
R19964 VBIAS.n1595 VBIAS.n1586 0.005
R19965 VBIAS.n1585 VBIAS.n1584 0.005
R19966 VBIAS.n1136 VBIAS.n1135 0.005
R19967 VBIAS.n1152 VBIAS.n1141 0.005
R19968 VBIAS.n1151 VBIAS.n1150 0.005
R19969 VBIAS.n1145 VBIAS.n1144 0.005
R19970 VBIAS.n1143 VBIAS.n1142 0.005
R19971 VBIAS.n1179 VBIAS.n1177 0.005
R19972 VBIAS.n1153 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE
+ 0.005
R19973 VBIAS.n1111 VBIAS.n1110 0.005
R19974 VBIAS.n1701 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE
+ 0.005
R19975 VBIAS.n1715 VBIAS.n1714 0.005
R19976 VBIAS.n1699 VBIAS.n1680 0.005
R19977 VBIAS.n1698 VBIAS.n1697 0.005
R19978 VBIAS.n1692 VBIAS.n1683 0.005
R19979 VBIAS.n1682 VBIAS.n1681 0.005
R19980 VBIAS.n1236 VBIAS.n1235 0.005
R19981 VBIAS.n1252 VBIAS.n1241 0.005
R19982 VBIAS.n1251 VBIAS.n1250 0.005
R19983 VBIAS.n1245 VBIAS.n1244 0.005
R19984 VBIAS.n1243 VBIAS.n1242 0.005
R19985 VBIAS.n1279 VBIAS.n1277 0.005
R19986 VBIAS.n1253 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE 0.005
R19987 VBIAS.n1211 VBIAS.n1210 0.005
R19988 VBIAS.n1778 VBIAS.n1776 0.005
R19989 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE VBIAS.n1782 0.005
R19990 VBIAS.n1787 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE 0.005
R19991 VBIAS.n1768 VBIAS.n1767 0.005
R19992 VBIAS.n1791 VBIAS.n1789 0.005
R19993 VBIAS.n1819 VBIAS.n1818 0.005
R19994 VBIAS.n1336 VBIAS.n1335 0.005
R19995 VBIAS.n1352 VBIAS.n1341 0.005
R19996 VBIAS.n1351 VBIAS.n1350 0.005
R19997 VBIAS.n1345 VBIAS.n1344 0.005
R19998 VBIAS.n1343 VBIAS.n1342 0.005
R19999 VBIAS.n1379 VBIAS.n1377 0.005
R20000 VBIAS.n1353 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE 0.005
R20001 VBIAS.n1311 VBIAS.n1310 0.005
R20002 VBIAS.n1845 VBIAS.n1843 0.005
R20003 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE VBIAS.n1849 0.005
R20004 VBIAS.n1854 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE 0.005
R20005 VBIAS.n1835 VBIAS.n1834 0.005
R20006 VBIAS.n1858 VBIAS.n1856 0.005
R20007 VBIAS.n1886 VBIAS.n1885 0.005
R20008 VBIAS.n1523 VBIAS.n1522 0.005
R20009 VBIAS.n1507 VBIAS.n1488 0.005
R20010 VBIAS.n1506 VBIAS.n1505 0.005
R20011 VBIAS.n1500 VBIAS.n1491 0.005
R20012 VBIAS.n1490 VBIAS.n1489 0.005
R20013 VBIAS.n1509 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE 0.005
R20014 VBIAS.n981 VBIAS.n979 0.005
R20015 VBIAS.n955 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE 0.005
R20016 VBIAS.n913 VBIAS.n912 0.005
R20017 VBIAS.n938 VBIAS.n937 0.005
R20018 VBIAS.n954 VBIAS.n943 0.005
R20019 VBIAS.n953 VBIAS.n952 0.005
R20020 VBIAS.n947 VBIAS.n946 0.005
R20021 VBIAS.n945 VBIAS.n944 0.005
R20022 VBIAS.n264 VBIAS.n263 0.005
R20023 VBIAS.n249 VBIAS.n215 0.005
R20024 VBIAS.n248 VBIAS.n247 0.005
R20025 VBIAS.n242 VBIAS.n218 0.005
R20026 VBIAS.n217 VBIAS.n216 0.005
R20027 VBIAS.n678 VBIAS.n676 0.005
R20028 VBIAS.n611 VBIAS.n610 0.005
R20029 VBIAS.n635 VBIAS.n634 0.005
R20030 VBIAS.n641 VBIAS.n640 0.005
R20031 VBIAS.n651 VBIAS.n650 0.005
R20032 VBIAS.n645 VBIAS.n644 0.005
R20033 VBIAS.n643 VBIAS.n642 0.005
R20034 VBIAS.n360 VBIAS.n359 0.005
R20035 VBIAS.n345 VBIAS.n311 0.005
R20036 VBIAS.n344 VBIAS.n343 0.005
R20037 VBIAS.n338 VBIAS.n314 0.005
R20038 VBIAS.n313 VBIAS.n312 0.005
R20039 VBIAS.n779 VBIAS.n777 0.005
R20040 VBIAS.n712 VBIAS.n711 0.005
R20041 VBIAS.n736 VBIAS.n735 0.005
R20042 VBIAS.n742 VBIAS.n741 0.005
R20043 VBIAS.n752 VBIAS.n751 0.005
R20044 VBIAS.n746 VBIAS.n745 0.005
R20045 VBIAS.n744 VBIAS.n743 0.005
R20046 VBIAS.n456 VBIAS.n455 0.005
R20047 VBIAS.n441 VBIAS.n407 0.005
R20048 VBIAS.n440 VBIAS.n439 0.005
R20049 VBIAS.n434 VBIAS.n410 0.005
R20050 VBIAS.n409 VBIAS.n408 0.005
R20051 VBIAS.n880 VBIAS.n878 0.005
R20052 VBIAS.n813 VBIAS.n812 0.005
R20053 VBIAS.n837 VBIAS.n836 0.005
R20054 VBIAS.n843 VBIAS.n842 0.005
R20055 VBIAS.n853 VBIAS.n852 0.005
R20056 VBIAS.n847 VBIAS.n846 0.005
R20057 VBIAS.n845 VBIAS.n844 0.005
R20058 VBIAS.n555 VBIAS.n554 0.005
R20059 VBIAS.n528 VBIAS.n527 0.005
R20060 VBIAS.n538 VBIAS.n537 0.005
R20061 VBIAS.n532 VBIAS.n531 0.005
R20062 VBIAS.n530 VBIAS.n529 0.005
R20063 VBIAS.n579 VBIAS.n577 0.005
R20064 VBIAS.n505 VBIAS.n504 0.005
R20065 VBIAS.n170 VBIAS.n169 0.005
R20066 VBIAS.n156 VBIAS.n122 0.005
R20067 VBIAS.n155 VBIAS.n154 0.005
R20068 VBIAS.n149 VBIAS.n125 0.005
R20069 VBIAS.n124 VBIAS.n123 0.005
R20070 VBIAS.n1957 VBIAS.n1956 0.005
R20071 VBIAS.n39 VBIAS.n38 0.005
R20072 VBIAS.n1889 VBIAS.n1861 0.004
R20073 VBIAS.n1822 VBIAS.n1794 0.004
R20074 VBIAS.n1755 VBIAS.n1754 0.004
R20075 VBIAS.n1658 VBIAS.n1657 0.004
R20076 VBIAS.n1561 VBIAS.n1560 0.004
R20077 VBIAS.n997 VBIAS.n996 0.004
R20078 VBIAS.n1097 VBIAS.n1096 0.004
R20079 VBIAS.n1197 VBIAS.n1196 0.004
R20080 VBIAS.n1297 VBIAS.n1296 0.004
R20081 VBIAS.n1397 VBIAS.n1396 0.004
R20082 VBIAS.n898 VBIAS.n897 0.004
R20083 VBIAS.n797 VBIAS.n796 0.004
R20084 VBIAS.n696 VBIAS.n695 0.004
R20085 VBIAS.n595 VBIAS.n594 0.004
R20086 VBIAS.n208 VBIAS.n207 0.004
R20087 VBIAS.n304 VBIAS.n303 0.004
R20088 VBIAS.n400 VBIAS.n399 0.004
R20089 VBIAS.n496 VBIAS.n495 0.004
R20090 VBIAS.n1968 VBIAS.n1966 0.004
R20091 VBIAS.n1972 VBIAS.n1970 0.004
R20092 VBIAS.n50 VBIAS.n48 0.004
R20093 VBIAS.n54 VBIAS.n52 0.004
R20094 VBIAS.n58 VBIAS.n14 0.004
R20095 VBIAS.n1977 VBIAS.n1976 0.004
R20096 VBIAS.n72 VBIAS.n71 0.004
R20097 VBIAS.n1930 VBIAS.n1929 0.004
R20098 VBIAS.n60 VBIAS.n59 0.003
R20099 VBIAS.n101 VBIAS.n100 0.003
R20100 VBIAS.n1898 VBIAS.n115 0.003
R20101 VBIAS.n108 VBIAS.n103 0.003
R20102 VBIAS.n92 VBIAS.n91 0.003
R20103 VBIAS.n1615 VBIAS.n1564 0.003
R20104 VBIAS.n1615 VBIAS.n1614 0.003
R20105 VBIAS.n1603 VBIAS.n1580 0.003
R20106 VBIAS.n1712 VBIAS.n1661 0.003
R20107 VBIAS.n1712 VBIAS.n1711 0.003
R20108 VBIAS.n1700 VBIAS.n1677 0.003
R20109 VBIAS.n1770 VBIAS.n1463 0.003
R20110 VBIAS.n1787 VBIAS.n1786 0.003
R20111 VBIAS.n1821 VBIAS.n1820 0.003
R20112 VBIAS.n1837 VBIAS.n1429 0.003
R20113 VBIAS.n1854 VBIAS.n1853 0.003
R20114 VBIAS.n1888 VBIAS.n1887 0.003
R20115 VBIAS.n1520 VBIAS.n1469 0.003
R20116 VBIAS.n1520 VBIAS.n1519 0.003
R20117 VBIAS.n1508 VBIAS.n1485 0.003
R20118 VBIAS.n261 VBIAS.n211 0.003
R20119 VBIAS.n261 VBIAS.n260 0.003
R20120 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE VBIAS.n212 0.003
R20121 VBIAS.n654 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE 0.003
R20122 VBIAS.n357 VBIAS.n307 0.003
R20123 VBIAS.n357 VBIAS.n356 0.003
R20124 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE VBIAS.n308 0.003
R20125 VBIAS.n755 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE 0.003
R20126 VBIAS.n453 VBIAS.n403 0.003
R20127 VBIAS.n453 VBIAS.n452 0.003
R20128 VBIAS VBIAS.n404 0.003
R20129 VBIAS.n856 VBIAS 0.003
R20130 VBIAS.n541 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE 0.003
R20131 VBIAS.n167 VBIAS.n117 0.003
R20132 VBIAS.n167 VBIAS.n166 0.003
R20133 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE VBIAS.n119 0.003
R20134 VBIAS.n1979 VBIAS.n1978 0.003
R20135 VBIAS.n1938 VBIAS.n1937 0.003
R20136 VBIAS.n1904 VBIAS.n1903 0.002
R20137 VBIAS.n1912 VBIAS.n1909 0.002
R20138 VBIAS.n1896 VBIAS.n1895 0.002
R20139 VBIAS.n1906 VBIAS.n1901 0.002
R20140 VBIAS.n98 VBIAS.n97 0.002
R20141 VBIAS.n1037 VBIAS.n1036 0.002
R20142 VBIAS.n1038 VBIAS.n1037 0.002
R20143 VBIAS.n1052 VBIAS.n1051 0.002
R20144 VBIAS.n1077 VBIAS.n1075 0.002
R20145 VBIAS.n1065 VBIAS.n1064 0.002
R20146 VBIAS.n1064 VBIAS.n1063 0.002
R20147 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE VBIAS.n1030 0.002
R20148 VBIAS.n1026 VBIAS.n1019 0.002
R20149 VBIAS.n1617 VBIAS.n1616 0.002
R20150 VBIAS.n1616 VBIAS.n1563 0.002
R20151 VBIAS.n1602 VBIAS.n1601 0.002
R20152 VBIAS.n1137 VBIAS.n1136 0.002
R20153 VBIAS.n1138 VBIAS.n1137 0.002
R20154 VBIAS.n1152 VBIAS.n1151 0.002
R20155 VBIAS.n1177 VBIAS.n1175 0.002
R20156 VBIAS.n1165 VBIAS.n1164 0.002
R20157 VBIAS.n1164 VBIAS.n1163 0.002
R20158 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE VBIAS.n1130
+ 0.002
R20159 VBIAS.n1126 VBIAS.n1119 0.002
R20160 VBIAS.n1714 VBIAS.n1713 0.002
R20161 VBIAS.n1713 VBIAS.n1660 0.002
R20162 VBIAS.n1699 VBIAS.n1698 0.002
R20163 VBIAS.n1237 VBIAS.n1236 0.002
R20164 VBIAS.n1238 VBIAS.n1237 0.002
R20165 VBIAS.n1252 VBIAS.n1251 0.002
R20166 VBIAS.n1277 VBIAS.n1275 0.002
R20167 VBIAS.n1265 VBIAS.n1264 0.002
R20168 VBIAS.n1264 VBIAS.n1263 0.002
R20169 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE VBIAS.n1230 0.002
R20170 VBIAS.n1226 VBIAS.n1219 0.002
R20171 VBIAS.n1769 VBIAS.n1768 0.002
R20172 VBIAS.n1789 VBIAS.n1788 0.002
R20173 VBIAS.n1337 VBIAS.n1336 0.002
R20174 VBIAS.n1338 VBIAS.n1337 0.002
R20175 VBIAS.n1352 VBIAS.n1351 0.002
R20176 VBIAS.n1377 VBIAS.n1375 0.002
R20177 VBIAS.n1365 VBIAS.n1364 0.002
R20178 VBIAS.n1364 VBIAS.n1363 0.002
R20179 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE VBIAS.n1330 0.002
R20180 VBIAS.n1326 VBIAS.n1319 0.002
R20181 VBIAS.n1836 VBIAS.n1835 0.002
R20182 VBIAS.n1856 VBIAS.n1855 0.002
R20183 VBIAS.n1833 VBIAS.n1832 0.002
R20184 VBIAS.n1859 VBIAS.n1400 0.002
R20185 VBIAS.n1766 VBIAS.n1765 0.002
R20186 VBIAS.n1792 VBIAS.n1434 0.002
R20187 VBIAS.n1750 VBIAS.n1749 0.002
R20188 VBIAS.n1752 VBIAS.n1751 0.002
R20189 VBIAS.n1653 VBIAS.n1652 0.002
R20190 VBIAS.n1655 VBIAS.n1654 0.002
R20191 VBIAS.n1556 VBIAS.n1555 0.002
R20192 VBIAS.n1558 VBIAS.n1557 0.002
R20193 VBIAS.n1522 VBIAS.n1521 0.002
R20194 VBIAS.n1521 VBIAS.n1468 0.002
R20195 VBIAS.n1507 VBIAS.n1506 0.002
R20196 VBIAS.n979 VBIAS.n977 0.002
R20197 VBIAS.n967 VBIAS.n966 0.002
R20198 VBIAS.n966 VBIAS.n965 0.002
R20199 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE VBIAS.n932 0.002
R20200 VBIAS.n928 VBIAS.n921 0.002
R20201 VBIAS.n939 VBIAS.n938 0.002
R20202 VBIAS.n940 VBIAS.n939 0.002
R20203 VBIAS.n954 VBIAS.n953 0.002
R20204 VBIAS.n992 VBIAS.n991 0.002
R20205 VBIAS.n994 VBIAS.n993 0.002
R20206 VBIAS.n1092 VBIAS.n1091 0.002
R20207 VBIAS.n1094 VBIAS.n1093 0.002
R20208 VBIAS.n1192 VBIAS.n1191 0.002
R20209 VBIAS.n1194 VBIAS.n1193 0.002
R20210 VBIAS.n1292 VBIAS.n1291 0.002
R20211 VBIAS.n1294 VBIAS.n1293 0.002
R20212 VBIAS.n1392 VBIAS.n1391 0.002
R20213 VBIAS.n1394 VBIAS.n1393 0.002
R20214 VBIAS.n263 VBIAS.n262 0.002
R20215 VBIAS.n262 VBIAS.n210 0.002
R20216 VBIAS.n249 VBIAS.n248 0.002
R20217 VBIAS.n676 VBIAS.n674 0.002
R20218 VBIAS.n664 VBIAS.n663 0.002
R20219 VBIAS.n663 VBIAS.n662 0.002
R20220 VBIAS.n653 VBIAS.n652 0.002
R20221 VBIAS.n626 VBIAS.n619 0.002
R20222 VBIAS.n636 VBIAS.n635 0.002
R20223 VBIAS.n637 VBIAS.n636 0.002
R20224 VBIAS.n651 VBIAS.n641 0.002
R20225 VBIAS.n359 VBIAS.n358 0.002
R20226 VBIAS.n358 VBIAS.n306 0.002
R20227 VBIAS.n345 VBIAS.n344 0.002
R20228 VBIAS.n777 VBIAS.n775 0.002
R20229 VBIAS.n765 VBIAS.n764 0.002
R20230 VBIAS.n764 VBIAS.n763 0.002
R20231 VBIAS.n754 VBIAS.n753 0.002
R20232 VBIAS.n727 VBIAS.n720 0.002
R20233 VBIAS.n737 VBIAS.n736 0.002
R20234 VBIAS.n738 VBIAS.n737 0.002
R20235 VBIAS.n752 VBIAS.n742 0.002
R20236 VBIAS.n455 VBIAS.n454 0.002
R20237 VBIAS.n454 VBIAS.n402 0.002
R20238 VBIAS.n441 VBIAS.n440 0.002
R20239 VBIAS.n878 VBIAS.n876 0.002
R20240 VBIAS.n866 VBIAS.n865 0.002
R20241 VBIAS.n865 VBIAS.n864 0.002
R20242 VBIAS.n855 VBIAS.n854 0.002
R20243 VBIAS.n828 VBIAS.n821 0.002
R20244 VBIAS.n838 VBIAS.n837 0.002
R20245 VBIAS.n839 VBIAS.n838 0.002
R20246 VBIAS.n853 VBIAS.n843 0.002
R20247 VBIAS.n893 VBIAS.n892 0.002
R20248 VBIAS.n895 VBIAS.n894 0.002
R20249 VBIAS.n792 VBIAS.n791 0.002
R20250 VBIAS.n794 VBIAS.n793 0.002
R20251 VBIAS.n691 VBIAS.n690 0.002
R20252 VBIAS.n693 VBIAS.n692 0.002
R20253 VBIAS.n590 VBIAS.n589 0.002
R20254 VBIAS.n592 VBIAS.n591 0.002
R20255 VBIAS.n554 VBIAS.n498 0.002
R20256 VBIAS.n524 VBIAS.n498 0.002
R20257 VBIAS.n538 VBIAS.n528 0.002
R20258 VBIAS.n577 VBIAS.n575 0.002
R20259 VBIAS.n553 VBIAS.n552 0.002
R20260 VBIAS.n552 VBIAS.n551 0.002
R20261 VBIAS.n540 VBIAS.n539 0.002
R20262 VBIAS.n520 VBIAS.n513 0.002
R20263 VBIAS.n169 VBIAS.n168 0.002
R20264 VBIAS.n168 VBIAS.n116 0.002
R20265 VBIAS.n156 VBIAS.n155 0.002
R20266 VBIAS.n203 VBIAS.n202 0.002
R20267 VBIAS.n205 VBIAS.n204 0.002
R20268 VBIAS.n299 VBIAS.n298 0.002
R20269 VBIAS.n301 VBIAS.n300 0.002
R20270 VBIAS.n395 VBIAS.n394 0.002
R20271 VBIAS.n397 VBIAS.n396 0.002
R20272 VBIAS.n491 VBIAS.n490 0.002
R20273 VBIAS.n493 VBIAS.n492 0.002
R20274 VBIAS.n4 VBIAS.n3 0.002
R20275 VBIAS.n1936 VBIAS.n1932 0.002
R20276 VBIAS.n80 VBIAS.n79 0.002
R20277 VBIAS.n29 VBIAS.n28 0.002
R20278 VBIAS.n1980 VBIAS.n1979 0.002
R20279 VBIAS.n94 VBIAS.n93 0.002
R20280 VBIAS.n112 VBIAS.n111 0.002
R20281 VBIAS.n110 VBIAS.n109 0.002
R20282 VBIAS.n1894 VBIAS.n1893 0.002
R20283 VBIAS.n106 VBIAS.n105 0.002
R20284 VBIAS.n1913 VBIAS.n108 0.002
R20285 VBIAS.n1913 VBIAS.n1898 0.002
R20286 VBIAS.n100 VBIAS.n99 0.002
R20287 VBIAS.n89 VBIAS.n60 0.002
R20288 VBIAS.n97 VBIAS.n96 0.001
R20289 VBIAS.n103 VBIAS.n102 0.001
R20290 VBIAS.n114 VBIAS.n113 0.001
R20291 VBIAS.n115 VBIAS.n114 0.001
R20292 VBIAS.n96 VBIAS.n95 0.001
R20293 VBIAS.n102 VBIAS.n101 0.001
R20294 VBIAS.n1905 VBIAS.n1904 0.001
R20295 VBIAS.n1897 VBIAS.n1896 0.001
R20296 VBIAS.n1912 VBIAS.n1911 0.001
R20297 VBIAS.n107 VBIAS.n104 0.001
R20298 VBIAS.n1906 VBIAS.n1905 0.001
R20299 VBIAS.n99 VBIAS.n98 0.001
R20300 VBIAS.n1937 VBIAS.n1924 0.001
R20301 VBIAS.n1911 VBIAS.n1910 0.001
R20302 VBIAS.n1897 VBIAS.n1894 0.001
R20303 VBIAS.n107 VBIAS.n106 0.001
R20304 VBIAS.n1060 VBIAS.n1056 0.001
R20305 VBIAS.n1611 VBIAS.n1608 0.001
R20306 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE VBIAS.n1603 0.001
R20307 VBIAS.n1160 VBIAS.n1156 0.001
R20308 VBIAS.n1708 VBIAS.n1705 0.001
R20309 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE VBIAS.n1700
+ 0.001
R20310 VBIAS.n1260 VBIAS.n1256 0.001
R20311 VBIAS.n1773 VBIAS.n1772 0.001
R20312 VBIAS.n1781 VBIAS.n1780 0.001
R20313 VBIAS.n1761 VBIAS.n1758 0.001
R20314 VBIAS.n1436 VBIAS.n1435 0.001
R20315 VBIAS.n1438 VBIAS.n1437 0.001
R20316 VBIAS.n1360 VBIAS.n1356 0.001
R20317 VBIAS.n1840 VBIAS.n1839 0.001
R20318 VBIAS.n1848 VBIAS.n1847 0.001
R20319 VBIAS.n1828 VBIAS.n1825 0.001
R20320 VBIAS.n1402 VBIAS.n1401 0.001
R20321 VBIAS.n1404 VBIAS.n1403 0.001
R20322 VBIAS.n1516 VBIAS.n1513 0.001
R20323 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE VBIAS.n1508 0.001
R20324 VBIAS.n962 VBIAS.n958 0.001
R20325 VBIAS.n257 VBIAS.n254 0.001
R20326 VBIAS.n660 VBIAS.n656 0.001
R20327 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE VBIAS.n653 0.001
R20328 VBIAS.n353 VBIAS.n350 0.001
R20329 VBIAS.n761 VBIAS.n757 0.001
R20330 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE VBIAS.n754 0.001
R20331 VBIAS.n449 VBIAS.n446 0.001
R20332 VBIAS.n862 VBIAS.n858 0.001
R20333 VBIAS VBIAS.n855 0.001
R20334 VBIAS.n548 VBIAS.n544 0.001
R20335 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE VBIAS.n540 0.001
R20336 VBIAS.n164 VBIAS.n161 0.001
R20337 VBIAS.n14 VBIAS.n13 0.001
R20338 VBIAS.n59 VBIAS.n58 0.001
R20339 VBIAS.n1976 VBIAS.n1938 0.001
R20340 VBIAS.n1978 VBIAS.n1977 0.001
R20341 VBIAS.n95 VBIAS.n94 0.001
R20342 VBIAS.n113 VBIAS.n112 0.001
R20343 VBIAS.n111 VBIAS.n110 0.001
R20344 VBIAS.n1903 VBIAS.n1902 0.001
R20345 VBIAS.n1900 VBIAS.n1899 0.001
R20346 VBIAS.n1908 VBIAS.n1907 0.001
R20347 VBIAS.n1909 VBIAS.n1908 0.001
R20348 VBIAS.n1901 VBIAS.n1900 0.001
R20349 VBIAS.n93 VBIAS.n92 0.001
R20350 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n43
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n686 9.305
R20351 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n44
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1257 9.305
R20352 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n45
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1184 9.305
R20353 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n46
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1123 9.305
R20354 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n47
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1071 9.305
R20355 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n48
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n996 9.305
R20356 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n49
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n935 9.305
R20357 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n320
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n319 9.304
R20358 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n290
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n289 9.304
R20359 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n666
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n665 9.304
R20360 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n616
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n615 9.304
R20361 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n562
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n561 9.304
R20362 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n512
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n511 9.304
R20363 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n458
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n457 9.304
R20364 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n408
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n407 9.304
R20365 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1707
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1706 9.304
R20366 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1657
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1656 9.304
R20367 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1603
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1602 9.304
R20368 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1553
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1552 9.304
R20369 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1499
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1498 9.304
R20370 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1449
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1448 9.304
R20371 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1395
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1394 9.304
R20372 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1345
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1344 9.304
R20373 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n325
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n324 9.3
R20374 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n51
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n353 9.3
R20375 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n39
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n342 9.3
R20376 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n359
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n358 9.3
R20377 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n313
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n312 9.3
R20378 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n316
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n318 9.3
R20379 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n364
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n363 9.3
R20380 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n206
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n360 9.3
R20381 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n347
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n346 9.3
R20382 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n345
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n344 9.3
R20383 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n50
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n351 9.3
R20384 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n336
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n335 9.3
R20385 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n51
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n354 9.3
R20386 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n661
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n664 9.3
R20387 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n55
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n656 9.3
R20388 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n13
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n645 9.3
R20389 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n629
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n628 9.3
R20390 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n678
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n677 9.3
R20391 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n669
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n673 9.3
R20392 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n625
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n624 9.3
R20393 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n208
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n627 9.3
R20394 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n650
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n649 9.3
R20395 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n648
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n647 9.3
R20396 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n54
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n654 9.3
R20397 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n641
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n640 9.3
R20398 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n55
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n657 9.3
R20399 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n595
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n594 9.3
R20400 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n57
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n601 9.3
R20401 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n587
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n586 9.3
R20402 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n610
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n609 9.3
R20403 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n593
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n592 9.3
R20404 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n57
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n602 9.3
R20405 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n56
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n599 9.3
R20406 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n619
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n622 9.3
R20407 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n557
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n560 9.3
R20408 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n59
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n552 9.3
R20409 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n17
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n541 9.3
R20410 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n525
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n524 9.3
R20411 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n574
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n573 9.3
R20412 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n565
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n569 9.3
R20413 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n521
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n520 9.3
R20414 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n209
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n523 9.3
R20415 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n546
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n545 9.3
R20416 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n544
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n543 9.3
R20417 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n58
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n550 9.3
R20418 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n537
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n536 9.3
R20419 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n59
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n553 9.3
R20420 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n491
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n490 9.3
R20421 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n61
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n497 9.3
R20422 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n483
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n482 9.3
R20423 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n506
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n505 9.3
R20424 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n489
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n488 9.3
R20425 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n61
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n498 9.3
R20426 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n60
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n495 9.3
R20427 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n515
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n518 9.3
R20428 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n453
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n456 9.3
R20429 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n63
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n448 9.3
R20430 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n21
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n437 9.3
R20431 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n421
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n420 9.3
R20432 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n470
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n469 9.3
R20433 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n461
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n465 9.3
R20434 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n417
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n416 9.3
R20435 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n210
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n419 9.3
R20436 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n442
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n441 9.3
R20437 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n440
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n439 9.3
R20438 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n62
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n446 9.3
R20439 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n433
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n432 9.3
R20440 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n63
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n449 9.3
R20441 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n387
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n386 9.3
R20442 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n65
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n393 9.3
R20443 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n379
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n378 9.3
R20444 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n402
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n401 9.3
R20445 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n385
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n384 9.3
R20446 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n65
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n394 9.3
R20447 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n64
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n391 9.3
R20448 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n411
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n414 9.3
R20449 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n66
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n912 9.3
R20450 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n907
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n906 9.3
R20451 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n922
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n921 9.3
R20452 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n66
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n913 9.3
R20453 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n67
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n911 9.3
R20454 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n905
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n904 9.3
R20455 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n901
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n900 9.3
R20456 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n880
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n879 9.3
R20457 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n877
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n876 9.3
R20458 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n873
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n872 9.3
R20459 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n109
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n871 9.3
R20460 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n890
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n889 9.3
R20461 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n894
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n893 9.3
R20462 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n896
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n895 9.3
R20463 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n697
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n696 9.3
R20464 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n690
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n689 9.3
R20465 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n721
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n720 9.3
R20466 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n710
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n709 9.3
R20467 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n736
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n735 9.3
R20468 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n719
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n718 9.3
R20469 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n715
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n714 9.3
R20470 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n708
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n707 9.3
R20471 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n703
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n702 9.3
R20472 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n69
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n725 9.3
R20473 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n68
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n727 9.3
R20474 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n68
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n726 9.3
R20475 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n694
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n693 9.3
R20476 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n830
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n829 9.3
R20477 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n861
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n860 9.3
R20478 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n846
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n845 9.3
R20479 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n813
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n812 9.3
R20480 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n70
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n835 9.3
R20481 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n70
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n836 9.3
R20482 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n71
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n834 9.3
R20483 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n828
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n827 9.3
R20484 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n824
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n823 9.3
R20485 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n848
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n847 9.3
R20486 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n865
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n864 9.3
R20487 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n868
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n867 9.3
R20488 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n854
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n853 9.3
R20489 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n111
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n859 9.3
R20490 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n72
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n265 9.3
R20491 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n229
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n228 9.3
R20492 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n253
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n252 9.3
R20493 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n259
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n258 9.3
R20494 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n248
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n247 9.3
R20495 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n246
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n245 9.3
R20496 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n233
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n232 9.3
R20497 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n236
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n235 9.3
R20498 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n242
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n241 9.3
R20499 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n257
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n256 9.3
R20500 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n73
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n263 9.3
R20501 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n72
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n266 9.3
R20502 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n274
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n273 9.3
R20503 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n113
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n227 9.3
R20504 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n74
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n176 9.3
R20505 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n74
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n175 9.3
R20506 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n169
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n168 9.3
R20507 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n75
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n173 9.3
R20508 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n164
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n163 9.3
R20509 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n167
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n166 9.3
R20510 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n202
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n201 9.3
R20511 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n199
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n198 9.3
R20512 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n195
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n194 9.3
R20513 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n115
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n193 9.3
R20514 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n153
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n152 9.3
R20515 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n157
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n156 9.3
R20516 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n159
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n158 9.3
R20517 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n184
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n183 9.3
R20518 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n774
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n773 9.3
R20519 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n77
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n788 9.3
R20520 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n76
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n790 9.3
R20521 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n76
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n789 9.3
R20522 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n799
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n798 9.3
R20523 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n772
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n771 9.3
R20524 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n767
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n766 9.3
R20525 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n761
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n760 9.3
R20526 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n757
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n756 9.3
R20527 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n753
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n752 9.3
R20528 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n117
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n751 9.3
R20529 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n779
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n778 9.3
R20530 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n782
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n781 9.3
R20531 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n784
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n783 9.3
R20532 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1261
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1260 9.3
R20533 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n79
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1299 9.3
R20534 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1282
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1281 9.3
R20535 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1265
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1264 9.3
R20536 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1269
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1268 9.3
R20537 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1275
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1274 9.3
R20538 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1291
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1290 9.3
R20539 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1293
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1292 9.3
R20540 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1287
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1286 9.3
R20541 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1280
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1279 9.3
R20542 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n78
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1297 9.3
R20543 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1251
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1250 9.3
R20544 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n79
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1300 9.3
R20545 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n81
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1238 9.3
R20546 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n80
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1236 9.3
R20547 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1219
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1218 9.3
R20548 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1221
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1220 9.3
R20549 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1226
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1225 9.3
R20550 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1230
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1229 9.3
R20551 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1232
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1231 9.3
R20552 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1214
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1213 9.3
R20553 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1196
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1195 9.3
R20554 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1192
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1191 9.3
R20555 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1188
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1187 9.3
R20556 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1208
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1207 9.3
R20557 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n81
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1239 9.3
R20558 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1148
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1147 9.3
R20559 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1141
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1140 9.3
R20560 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1153
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1152 9.3
R20561 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n82
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1163 9.3
R20562 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n83
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1165 9.3
R20563 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1159
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1158 9.3
R20564 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1157
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1156 9.3
R20565 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n83
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1166 9.3
R20566 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1176
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1175 9.3
R20567 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1131
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1130 9.3
R20568 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1127
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1126 9.3
R20569 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1135
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1134 9.3
R20570 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1146
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1145 9.3
R20571 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1075
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1074 9.3
R20572 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n85
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1113 9.3
R20573 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1096
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1095 9.3
R20574 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1079
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1078 9.3
R20575 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1083
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1082 9.3
R20576 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1089
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1088 9.3
R20577 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1105
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1104 9.3
R20578 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1107
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1106 9.3
R20579 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1101
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1100 9.3
R20580 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1094
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1093 9.3
R20581 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n84
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1111 9.3
R20582 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1065
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1064 9.3
R20583 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n85
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1114 9.3
R20584 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n87
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1050 9.3
R20585 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n86
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1048 9.3
R20586 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1031
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1030 9.3
R20587 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1033
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1032 9.3
R20588 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1038
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1037 9.3
R20589 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1042
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1041 9.3
R20590 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1044
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1043 9.3
R20591 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1026
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1025 9.3
R20592 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1008
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1007 9.3
R20593 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1004
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1003 9.3
R20594 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1000
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n999 9.3
R20595 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1020
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1019 9.3
R20596 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n87
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1051 9.3
R20597 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n960
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n959 9.3
R20598 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n953
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n952 9.3
R20599 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n965
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n964 9.3
R20600 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n88
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n975 9.3
R20601 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n89
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n977 9.3
R20602 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n971
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n970 9.3
R20603 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n969
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n968 9.3
R20604 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n89
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n978 9.3
R20605 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n988
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n987 9.3
R20606 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n943
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n942 9.3
R20607 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n939
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n938 9.3
R20608 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n947
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n946 9.3
R20609 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n958
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n957 9.3
R20610 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1702
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1705 9.3
R20611 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n91
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1697 9.3
R20612 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n25
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1686 9.3
R20613 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1670
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1669 9.3
R20614 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1719
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1718 9.3
R20615 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1710
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1714 9.3
R20616 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1666
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1665 9.3
R20617 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n211
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1668 9.3
R20618 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1691
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1690 9.3
R20619 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1689
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1688 9.3
R20620 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n90
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1695 9.3
R20621 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1682
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1681 9.3
R20622 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n91
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1698 9.3
R20623 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1636
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1635 9.3
R20624 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n93
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1642 9.3
R20625 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1628
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1627 9.3
R20626 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1651
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1650 9.3
R20627 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1634
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1633 9.3
R20628 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n93
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1643 9.3
R20629 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n92
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1640 9.3
R20630 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1660
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1663 9.3
R20631 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1598
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1601 9.3
R20632 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n95
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1593 9.3
R20633 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n29
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1582 9.3
R20634 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1566
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1565 9.3
R20635 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1615
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1614 9.3
R20636 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1606
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1610 9.3
R20637 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1562
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1561 9.3
R20638 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n212
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1564 9.3
R20639 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1587
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1586 9.3
R20640 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1585
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1584 9.3
R20641 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n94
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1591 9.3
R20642 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1578
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1577 9.3
R20643 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n95
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1594 9.3
R20644 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1532
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1531 9.3
R20645 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n97
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1538 9.3
R20646 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1524
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1523 9.3
R20647 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1547
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1546 9.3
R20648 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1530
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1529 9.3
R20649 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n97
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1539 9.3
R20650 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n96
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1536 9.3
R20651 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1556
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1559 9.3
R20652 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1494
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1497 9.3
R20653 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n99
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1489 9.3
R20654 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n33
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1478 9.3
R20655 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1462
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1461 9.3
R20656 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1511
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1510 9.3
R20657 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1502
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1506 9.3
R20658 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1458
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1457 9.3
R20659 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n213
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1460 9.3
R20660 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1483
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1482 9.3
R20661 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1481
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1480 9.3
R20662 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n98
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1487 9.3
R20663 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1474
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1473 9.3
R20664 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n99
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1490 9.3
R20665 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1428
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1427 9.3
R20666 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n101
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1434 9.3
R20667 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1420
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1419 9.3
R20668 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1443
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1442 9.3
R20669 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1426
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1425 9.3
R20670 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n101
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1435 9.3
R20671 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n100
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1432 9.3
R20672 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1452
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1455 9.3
R20673 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1390
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1393 9.3
R20674 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n103
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1385 9.3
R20675 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n37
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1374 9.3
R20676 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1358
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1357 9.3
R20677 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1407
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1406 9.3
R20678 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1398
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1402 9.3
R20679 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1354
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1353 9.3
R20680 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n214
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1356 9.3
R20681 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1379
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1378 9.3
R20682 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1377
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1376 9.3
R20683 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n102
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1383 9.3
R20684 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1370
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1369 9.3
R20685 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n103
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1386 9.3
R20686 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1324
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1323 9.3
R20687 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n105
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1330 9.3
R20688 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1316
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1315 9.3
R20689 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1339
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1338 9.3
R20690 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1322
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1321 9.3
R20691 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n105
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1331 9.3
R20692 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n104
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1328 9.3
R20693 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1348
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1351 9.3
R20694 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1743
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1742 9.3
R20695 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n53
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1749 9.3
R20696 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1730
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1729 9.3
R20697 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n288
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n287 9.3
R20698 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n307
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n306 9.3
R20699 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n207
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n285 9.3
R20700 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1741
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1740 9.3
R20701 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n53
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1750 9.3
R20702 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n293
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n296 9.3
R20703 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n301
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n300 9.3
R20704 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n283
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n282 9.3
R20705 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n41
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1738 9.3
R20706 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n52
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1747 9.3
R20707 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n12
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n591 9
R20708 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n56
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n600 9
R20709 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n604
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n603 9
R20710 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n585
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n581 9
R20711 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n639
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n635 9
R20712 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n680
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n679 9
R20713 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n14
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n646 9
R20714 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n612
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n611 9
R20715 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n618
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n617 9
R20716 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n106
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n626 9
R20717 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n659
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n658 9
R20718 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n54
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n655 9
R20719 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n668
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n667 9
R20720 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n16
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n487 9
R20721 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n60
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n496 9
R20722 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n500
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n499 9
R20723 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n481
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n477 9
R20724 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n535
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n531 9
R20725 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n576
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n575 9
R20726 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n18
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n542 9
R20727 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n508
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n507 9
R20728 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n514
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n513 9
R20729 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n107
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n522 9
R20730 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n555
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n554 9
R20731 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n58
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n551 9
R20732 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n564
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n563 9
R20733 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n20
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n383 9
R20734 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n64
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n392 9
R20735 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n396
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n395 9
R20736 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n377
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n373 9
R20737 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n431
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n427 9
R20738 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n472
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n471 9
R20739 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n22
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n438 9
R20740 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n404
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n403 9
R20741 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n410
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n409 9
R20742 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n108
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n418 9
R20743 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n451
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n450 9
R20744 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n62
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n447 9
R20745 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n460
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n459 9
R20746 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n71
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n820 9
R20747 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n826
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n825 9
R20748 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n110
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n870 9
R20749 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n878
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n869 9
R20750 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n866
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n857 9
R20751 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n811
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n810 9
R20752 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n69
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n684 9
R20753 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n717
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n716 9
R20754 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n705
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n704 9
R20755 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n838
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n837 9
R20756 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n851
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n850 9
R20757 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n891
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n886 9
R20758 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n920
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n919 9
R20759 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n915
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n914 9
R20760 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n729
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n728 9
R20761 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n734
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n733 9
R20762 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n67
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n885 9
R20763 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n903
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n902 9
R20764 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n112
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n858 9
R20765 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n43
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n687 9
R20766 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n695
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n685 9
R20767 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n797
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n796 9
R20768 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n267
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n223 9
R20769 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n73
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n264 9
R20770 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n165
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n148 9
R20771 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n780
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n749 9
R20772 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n769
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n768 9
R20773 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n759
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n758 9
R20774 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n118
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n750 9
R20775 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n116
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n192 9
R20776 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n200
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n191 9
R20777 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n234
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n225 9
R20778 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n272
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n271 9
R20779 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n243
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n224 9
R20780 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n154
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n149 9
R20781 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n177
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n147 9
R20782 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n77
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n748 9
R20783 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n792
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n791 9
R20784 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n75
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n174 9
R20785 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n255
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n254 9
R20786 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n114
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n226 9
R20787 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n182
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n181 9
R20788 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1174
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1170 9
R20789 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1249
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1245 9
R20790 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n45
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1185 9
R20791 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1194
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1193 9
R20792 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1155
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1154 9
R20793 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n82
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1164 9
R20794 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1267
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1266 9
R20795 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1289
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1288 9
R20796 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1277
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1276 9
R20797 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1228
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1227 9
R20798 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n80
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1237 9
R20799 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1216
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1215 9
R20800 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1206
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1202 9
R20801 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1241
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1240 9
R20802 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n78
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1298 9
R20803 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1302
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1301 9
R20804 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1181
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1180 9
R20805 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n46
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1124 9
R20806 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1133
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1132 9
R20807 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n44
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1258 9
R20808 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1143
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1142 9
R20809 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n986
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n982 9
R20810 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1063
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1059 9
R20811 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n48
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n997 9
R20812 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1006
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1005 9
R20813 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n967
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n966 9
R20814 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n88
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n976 9
R20815 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1081
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1080 9
R20816 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1103
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1102 9
R20817 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1091
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1090 9
R20818 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1040
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1039 9
R20819 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n86
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1049 9
R20820 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1028
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1027 9
R20821 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1018
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1014 9
R20822 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1053
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1052 9
R20823 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n84
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1112 9
R20824 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1116
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1115 9
R20825 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n993
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n992 9
R20826 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n49
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n936 9
R20827 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n945
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n944 9
R20828 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n47
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1072 9
R20829 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n955
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n954 9
R20830 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n24
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1632 9
R20831 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n92
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1641 9
R20832 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1645
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1644 9
R20833 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1626
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1622 9
R20834 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1680
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1676 9
R20835 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1721
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1720 9
R20836 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n26
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1687 9
R20837 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1653
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1652 9
R20838 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1659
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1658 9
R20839 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n119
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1667 9
R20840 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1700
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1699 9
R20841 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n90
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1696 9
R20842 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1709
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1708 9
R20843 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n28
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1528 9
R20844 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n96
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1537 9
R20845 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1541
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1540 9
R20846 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1522
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1518 9
R20847 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1576
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1572 9
R20848 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1617
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1616 9
R20849 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n30
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1583 9
R20850 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1549
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1548 9
R20851 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1555
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1554 9
R20852 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n120
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1563 9
R20853 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1596
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1595 9
R20854 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n94
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1592 9
R20855 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1605
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1604 9
R20856 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n32
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1424 9
R20857 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n100
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1433 9
R20858 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1437
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1436 9
R20859 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1418
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1414 9
R20860 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1472
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1468 9
R20861 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1513
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1512 9
R20862 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n34
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1479 9
R20863 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1445
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1444 9
R20864 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1451
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1450 9
R20865 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n121
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1459 9
R20866 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1492
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1491 9
R20867 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n98
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1488 9
R20868 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1501
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1500 9
R20869 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n36
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1320 9
R20870 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n104
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1329 9
R20871 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1333
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1332 9
R20872 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1314
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1310 9
R20873 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1368
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1364 9
R20874 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1409
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1408 9
R20875 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n38
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1375 9
R20876 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1341
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1340 9
R20877 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1347
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1346 9
R20878 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n122
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1355 9
R20879 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1388
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1387 9
R20880 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n102
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1384 9
R20881 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1397
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1396 9
R20882 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n334
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n330 9
R20883 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n315
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n314 9
R20884 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n40
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n343 9
R20885 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n123
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n361 9
R20886 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n356
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n355 9
R20887 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n50
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n352 9
R20888 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n322
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n321 9
R20889 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n42
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1739 9
R20890 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n52
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1748 9
R20891 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1752
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1751 9
R20892 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1728
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1727 9
R20893 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n124
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n284 9
R20894 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n303
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n302 9
R20895 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n292
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n291 9
R20896 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n643
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n634 4.574
R20897 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n589
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n580 4.574
R20898 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n539
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n530 4.574
R20899 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n485
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n476 4.574
R20900 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n435
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n426 4.574
R20901 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n381
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n372 4.574
R20902 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n818
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n817 4.574
R20903 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n927
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n926 4.574
R20904 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n741
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n740 4.574
R20905 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n279
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n278 4.574
R20906 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n804
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n803 4.574
R20907 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n189
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n188 4.574
R20908 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1210
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1201 4.574
R20909 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1256
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1255 4.574
R20910 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1178
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1169 4.574
R20911 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1022
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1013 4.574
R20912 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1070
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1069 4.574
R20913 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n990
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n981 4.574
R20914 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1684
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1675 4.574
R20915 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1630
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1621 4.574
R20916 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1580
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1571 4.574
R20917 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1526
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1517 4.574
R20918 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1476
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1467 4.574
R20919 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1422
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1413 4.574
R20920 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1372
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1363 4.574
R20921 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1318
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1309 4.574
R20922 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n338
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n329 4.574
R20923 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1735
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1734 4.574
R20924 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n329
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n328 3.388
R20925 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n634
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n633 3.388
R20926 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n580
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n579 3.388
R20927 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n530
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n529 3.388
R20928 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n476
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n475 3.388
R20929 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n426
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n425 3.388
R20930 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n372
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n371 3.388
R20931 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n926
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n924 3.388
R20932 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n740
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n738 3.388
R20933 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n817
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n815 3.388
R20934 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n278
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n276 3.388
R20935 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n188
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n186 3.388
R20936 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n803
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n801 3.388
R20937 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1255
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1254 3.388
R20938 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1201
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1200 3.388
R20939 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1169
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1168 3.388
R20940 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1069
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1068 3.388
R20941 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1013
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1012 3.388
R20942 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n981
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n980 3.388
R20943 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1675
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1674 3.388
R20944 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1621
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1620 3.388
R20945 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1571
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1570 3.388
R20946 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1517
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1516 3.388
R20947 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1467
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1466 3.388
R20948 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1413
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1412 3.388
R20949 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1363
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1362 3.388
R20950 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1309
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1308 3.388
R20951 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1734
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1733 3.388
R20952 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n331
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t38 3.326
R20953 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n331
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t23 3.326
R20954 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n636
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t47 3.326
R20955 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n636
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t22 3.326
R20956 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n582
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t34 3.326
R20957 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n582
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t35 3.326
R20958 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n532
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t40 3.326
R20959 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n532
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t25 3.326
R20960 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n478
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t36 3.326
R20961 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n478
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t37 3.326
R20962 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n428
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t45 3.326
R20963 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n428
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t20 3.326
R20964 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n374
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t27 3.326
R20965 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n374
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t44 3.326
R20966 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n916
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t8 3.326
R20967 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n916
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t1 3.326
R20968 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n730
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t5 3.326
R20969 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n807
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t13 3.326
R20970 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n268
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t2 3.326
R20971 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n178
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t10 3.326
R20972 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n178
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t6 3.326
R20973 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n793
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t11 3.326
R20974 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1246
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t15 3.326
R20975 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1203
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t14 3.326
R20976 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1203
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t12 3.326
R20977 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1171
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t0 3.326
R20978 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1060
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t4 3.326
R20979 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1015
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t9 3.326
R20980 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1015
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t3 3.326
R20981 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n983
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t7 3.326
R20982 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1677
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t42 3.326
R20983 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1677
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t17 3.326
R20984 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1623
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t29 3.326
R20985 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1623
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t30 3.326
R20986 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1573
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t33 3.326
R20987 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1573
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t21 3.326
R20988 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1519
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t28 3.326
R20989 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1519
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t32 3.326
R20990 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1469
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t41 3.326
R20991 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1469
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t16 3.326
R20992 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1415
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t26 3.326
R20993 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1415
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t39 3.326
R20994 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1365
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t31 3.326
R20995 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1365
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t18 3.326
R20996 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1311
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t19 3.326
R20997 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1311
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t43 3.326
R20998 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1724
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t24 3.326
R20999 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1724
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t46 3.326
R21000 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n843
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n842 2.481
R21001 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n607 2.473
R21002 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n503 2.473
R21003 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n399 2.473
R21004 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1648 2.473
R21005 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1544 2.473
R21006 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1440 2.473
R21007 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1336 2.473
R21008 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n207 2.473
R21009 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n215
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n631 2.473
R21010 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n216
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n527 2.473
R21011 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n217
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n423 2.473
R21012 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n218
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1672 2.473
R21013 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n219
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1568 2.473
R21014 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n220
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1464 2.473
R21015 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n221
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1360 2.473
R21016 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n222
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n366 2.473
R21017 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n215
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n662 2.469
R21018 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n215
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n670 2.469
R21019 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n620 2.469
R21020 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n613 2.469
R21021 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n216
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n558 2.469
R21022 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n216
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n566 2.469
R21023 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n516 2.469
R21024 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n509 2.469
R21025 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n217
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n454 2.469
R21026 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n217
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n462 2.469
R21027 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n412 2.469
R21028 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n405 2.469
R21029 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n218
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1703 2.469
R21030 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n218
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1711 2.469
R21031 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1661 2.469
R21032 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1654 2.469
R21033 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n219
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1599 2.469
R21034 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n219
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1607 2.469
R21035 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1557 2.469
R21036 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1550 2.469
R21037 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n220
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1495 2.469
R21038 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n220
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1503 2.469
R21039 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1453 2.469
R21040 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1446 2.469
R21041 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n221
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1391 2.469
R21042 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n221
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1399 2.469
R21043 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1349 2.469
R21044 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1342 2.469
R21045 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n222
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n326 2.469
R21046 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n308 2.469
R21047 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n294 2.469
R21048 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n222
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n317 2.469
R21049 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n215
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n660 2.235
R21050 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n216
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n556 2.235
R21051 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n217
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n452 2.235
R21052 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n218
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1701 2.235
R21053 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n219
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1597 2.235
R21054 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n220
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1493 2.235
R21055 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n221
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1389 2.235
R21056 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n222
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n357 2.235
R21057 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1183
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1198 2.232
R21058 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n995
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1010 2.232
R21059 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n884
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n882 2.232
R21060 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n205
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n204 2.232
R21061 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n605 2.231
R21062 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n501 2.231
R21063 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n397 2.231
R21064 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1646 2.231
R21065 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1542 2.231
R21066 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1438 2.231
R21067 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1334 2.231
R21068 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1753 2.231
R21069 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n125
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n742 2.23
R21070 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n126
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n805 2.23
R21071 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n128
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1303 2.23
R21072 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n129
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1117 2.23
R21073 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1121
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1181 1.94
R21074 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n933
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n993 1.94
R21075 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n884
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n928 1.779
R21076 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n205
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n190 1.779
R21077 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1183
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1242 1.779
R21078 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n995
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1054 1.779
R21079 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n917
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n916 1.155
R21080 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n179
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n178 1.155
R21081 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1247
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1246 1.155
R21082 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1061
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1060 1.155
R21083 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1725
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1724 1.155
R21084 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n332
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n331 1.155
R21085 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n637
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n636 1.155
R21086 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n533
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n532 1.155
R21087 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n429
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n428 1.155
R21088 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1678
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1677 1.155
R21089 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1574
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1573 1.155
R21090 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1470
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1469 1.155
R21091 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1366
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1365 1.155
R21092 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n583
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n582 1.155
R21093 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n479
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n478 1.155
R21094 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n375
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n374 1.155
R21095 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1204
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1203 1.155
R21096 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1016
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1015 1.155
R21097 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1624
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1623 1.155
R21098 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1520
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1519 1.155
R21099 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1416
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1415 1.155
R21100 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1312
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1311 1.155
R21101 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n794
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n793 1.155
R21102 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1172
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1171 1.155
R21103 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n984
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n983 1.155
R21104 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n731
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n730 1.155
R21105 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n808
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n807 1.155
R21106 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n269
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n268 1.155
R21107 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n918
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n917 0.921
R21108 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n732
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n731 0.921
R21109 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n333
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n332 0.921
R21110 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n638
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n637 0.921
R21111 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n534
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n533 0.921
R21112 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n430
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n429 0.921
R21113 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1679
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1678 0.921
R21114 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1575
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1574 0.921
R21115 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1471
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1470 0.921
R21116 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1367
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1366 0.921
R21117 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n584
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n583 0.921
R21118 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n480
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n479 0.921
R21119 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n376
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n375 0.921
R21120 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1205
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1204 0.921
R21121 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1017
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1016 0.921
R21122 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1625
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1624 0.921
R21123 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1521
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1520 0.921
R21124 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1417
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1416 0.921
R21125 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1313
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1312 0.921
R21126 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n795
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n794 0.921
R21127 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1248
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1247 0.921
R21128 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1062
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1061 0.921
R21129 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1726
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1725 0.921
R21130 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n809
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n808 0.921
R21131 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n270
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n269 0.921
R21132 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1173
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1172 0.921
R21133 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n985
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n984 0.921
R21134 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n180
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n179 0.903
R21135 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n329
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n327 0.506
R21136 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n634
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n632 0.506
R21137 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n580
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n578 0.506
R21138 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n530
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n528 0.506
R21139 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n476
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n474 0.506
R21140 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n426
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n424 0.506
R21141 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n372
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n370 0.506
R21142 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n926
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n925 0.506
R21143 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n740
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n739 0.506
R21144 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n817
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n816 0.506
R21145 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n278
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n277 0.506
R21146 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n188
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n187 0.506
R21147 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1201
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1199 0.506
R21148 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1169
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1167 0.506
R21149 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1013
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1011 0.506
R21150 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n981
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n979 0.506
R21151 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1675
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1673 0.506
R21152 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1621
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1619 0.506
R21153 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1571
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1569 0.506
R21154 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1517
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1515 0.506
R21155 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1467
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1465 0.506
R21156 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1413
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1411 0.506
R21157 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1363
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1361 0.506
R21158 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1309
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1307 0.506
R21159 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n803
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n802 0.506
R21160 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1255
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1253 0.506
R21161 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1069
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1067 0.506
R21162 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1734
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1732 0.506
R21163 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n682
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n126 0.494
R21164 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1058
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n128 0.494
R21165 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1722
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1305 0.49
R21166 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n351
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n350 0.476
R21167 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n654
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n653 0.476
R21168 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n599
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n598 0.476
R21169 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n550
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n549 0.476
R21170 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n495
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n494 0.476
R21171 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n446
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n445 0.476
R21172 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n391
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n390 0.476
R21173 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n911
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n910 0.476
R21174 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n725
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n724 0.476
R21175 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n834
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n833 0.476
R21176 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n263
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n262 0.476
R21177 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n173
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n172 0.476
R21178 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n788
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n787 0.476
R21179 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1236
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1235 0.476
R21180 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1048
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1047 0.476
R21181 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1695
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1694 0.476
R21182 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1640
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1639 0.476
R21183 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1591
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1590 0.476
R21184 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1536
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1535 0.476
R21185 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1487
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1486 0.476
R21186 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1432
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1431 0.476
R21187 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1383
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1382 0.476
R21188 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1328
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1327 0.476
R21189 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1297
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1296 0.475
R21190 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1163
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1162 0.475
R21191 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1111
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1110 0.475
R21192 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n975
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n974 0.475
R21193 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1747
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1746 0.475
R21194 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n127
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n125 0.468
R21195 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n130
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n129 0.468
R21196 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n342
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n341 0.445
R21197 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n645
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n644 0.445
R21198 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n11
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n590 0.445
R21199 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n541
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n540 0.445
R21200 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n15
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n486 0.445
R21201 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n437
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n436 0.445
R21202 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n19
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n382 0.445
R21203 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n900
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n899 0.445
R21204 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n714
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n713 0.445
R21205 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n823
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n822 0.445
R21206 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n252
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n251 0.445
R21207 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n163
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n162 0.445
R21208 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1225
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1224 0.445
R21209 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1037
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1036 0.445
R21210 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1686
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1685 0.445
R21211 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n23
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1631 0.445
R21212 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1582
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1581 0.445
R21213 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n27
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1527 0.445
R21214 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1478
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1477 0.445
R21215 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n31
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1423 0.445
R21216 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1374
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1373 0.445
R21217 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n35
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1319 0.445
R21218 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n778
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n777 0.445
R21219 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1286
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1285 0.445
R21220 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1152
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1151 0.445
R21221 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1100
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1099 0.445
R21222 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n964
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n963 0.445
R21223 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1738
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1737 0.445
R21224 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1305
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n681 0.432
R21225 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1722 0.427
R21226 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n363
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n362 0.414
R21227 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n624
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n623 0.414
R21228 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n520
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n519 0.414
R21229 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n416
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n415 0.414
R21230 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n889
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n888 0.414
R21231 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n702
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n701 0.414
R21232 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n853
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n852 0.414
R21233 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n241
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n240 0.414
R21234 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n152
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n151 0.414
R21235 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n766
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n765 0.414
R21236 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1213
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1212 0.414
R21237 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1025
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1024 0.414
R21238 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1665
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1664 0.414
R21239 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1561
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1560 0.414
R21240 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1457
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1456 0.414
R21241 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1353
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1352 0.414
R21242 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1140
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1139 0.413
R21243 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n952
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n951 0.413
R21244 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1274
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1273 0.413
R21245 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1088
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1087 0.413
R21246 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n282
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n281 0.413
R21247 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n312
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n311 0.382
R21248 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n677
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n676 0.382
R21249 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n609
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n608 0.382
R21250 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n573
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n572 0.382
R21251 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n505
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n504 0.382
R21252 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n469
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n468 0.382
R21253 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n401
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n400 0.382
R21254 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n876
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n875 0.382
R21255 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n693
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n692 0.382
R21256 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n864
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n863 0.382
R21257 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n232
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n231 0.382
R21258 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n198
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n197 0.382
R21259 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1191
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1190 0.382
R21260 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1003
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1002 0.382
R21261 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1718
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1717 0.382
R21262 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1650
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1649 0.382
R21263 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1614
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1613 0.382
R21264 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1546
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1545 0.382
R21265 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1510
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1509 0.382
R21266 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1442
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1441 0.382
R21267 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1406
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1405 0.382
R21268 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1338
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1337 0.382
R21269 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n300
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n299 0.382
R21270 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n756
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n755 0.382
R21271 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1264
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1263 0.382
R21272 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1130
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1129 0.382
R21273 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1078
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1077 0.382
R21274 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n942
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n941 0.382
R21275 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n747
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n205 0.341
R21276 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1305
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1057 0.33
R21277 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n744
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n280 2.648
R21278 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n840
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n838 2.887
R21279 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n930
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n843 0.31
R21280 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1244
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1122 0.31
R21281 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1056
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n934 0.31
R21282 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n144
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1755 0.299
R21283 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n142
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1756 0.299
R21284 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n140
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1757 0.299
R21285 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n137
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1758 0.299
R21286 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n135
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1759 0.299
R21287 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n133
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1760 0.299
R21288 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n131
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1761 0.299
R21289 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n131
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n221 0.295
R21290 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n133
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n220 0.295
R21291 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n135
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n219 0.295
R21292 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n137
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n218 0.295
R21293 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n140
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n217 0.295
R21294 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n142
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n216 0.295
R21295 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n144
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n215 0.295
R21296 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n141
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8 0.294
R21297 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n143
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9 0.294
R21298 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n146
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10 0.294
R21299 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n132
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4 0.294
R21300 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n134
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5 0.294
R21301 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n136
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6 0.294
R21302 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n139
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7 0.294
R21303 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n2
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n368 0.213
R21304 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n141
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n143 0.116
R21305 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n134
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n136 0.116
R21306 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n839
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n930 0.095
R21307 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n743
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n747 0.095
R21308 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n931
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1056 0.095
R21309 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1119
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1244 0.095
R21310 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1722
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n132 0.078
R21311 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n862
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n861 0.077
R21312 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n230
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n229 0.077
R21313 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1128
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1127 0.077
R21314 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1262
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1261 0.077
R21315 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n940
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n939 0.077
R21316 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1076
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1075 0.077
R21317 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n874
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n873 0.077
R21318 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n691
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n690 0.077
R21319 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n196
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n195 0.077
R21320 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n754
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n753 0.077
R21321 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1189
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1188 0.077
R21322 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1001
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1000 0.077
R21323 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n838
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n819 0.075
R21324 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n897
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n896 0.073
R21325 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n160
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n159 0.073
R21326 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1222
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1221 0.073
R21327 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1034
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1033 0.073
R21328 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n368
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1 0.068
R21329 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n928
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n927 0.064
R21330 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n190
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n189 0.064
R21331 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1242
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1210 0.063
R21332 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1054
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1022 0.063
R21333 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n908
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n907 0.063
R21334 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n170
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n169 0.063
R21335 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n348
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n347 0.06
R21336 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n288
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n286 0.06
R21337 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1744
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1743 0.06
R21338 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n630
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n629 0.06
R21339 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n651
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n650 0.06
R21340 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n596
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n595 0.06
R21341 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n526
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n525 0.06
R21342 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n547
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n546 0.06
R21343 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n492
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n491 0.06
R21344 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n422
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n421 0.06
R21345 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n443
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n442 0.06
R21346 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n388
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n387 0.06
R21347 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n711
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n710 0.06
R21348 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n846
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n844 0.06
R21349 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n249
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n248 0.06
R21350 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n775
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n774 0.06
R21351 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1283
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1282 0.06
R21352 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1149
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1148 0.06
R21353 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1097
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1096 0.06
R21354 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n961
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n960 0.06
R21355 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1671
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1670 0.06
R21356 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1692
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1691 0.06
R21357 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1637
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1636 0.06
R21358 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1567
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1566 0.06
R21359 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1588
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1587 0.06
R21360 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1533
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1532 0.06
R21361 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1463
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1462 0.06
R21362 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1484
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1483 0.06
R21363 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1429
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1428 0.06
R21364 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1359
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1358 0.06
R21365 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1380
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1379 0.06
R21366 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1325
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1324 0.06
R21367 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1181
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1179 0.058
R21368 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n993
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n991 0.058
R21369 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n805
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n792 0.057
R21370 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n280
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n267 0.057
R21371 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1303
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1302 0.057
R21372 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1117
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1116 0.057
R21373 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n742
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n729 0.057
R21374 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n143
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n146 0.055
R21375 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n141 0.055
R21376 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n136
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n139 0.055
R21377 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n132
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n134 0.055
R21378 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1753
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1735 0.054
R21379 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n660
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n643 0.054
R21380 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n605
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n589 0.054
R21381 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n556
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n539 0.054
R21382 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n501
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n485 0.054
R21383 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n452
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n435 0.054
R21384 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n397
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n381 0.054
R21385 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1701
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1684 0.054
R21386 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1646
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1630 0.054
R21387 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1597
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1580 0.054
R21388 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1542
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1526 0.054
R21389 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1493
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1476 0.054
R21390 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1438
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1422 0.054
R21391 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1389
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1372 0.054
R21392 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1334
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1318 0.054
R21393 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n357
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n338 0.054
R21394 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n357
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n356 0.054
R21395 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n660
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n659 0.054
R21396 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n605
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n604 0.054
R21397 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n556
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n555 0.054
R21398 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n501
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n500 0.054
R21399 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n452
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n451 0.054
R21400 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n397
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n396 0.054
R21401 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1701
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1700 0.054
R21402 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1646
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1645 0.054
R21403 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1597
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1596 0.054
R21404 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1542
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1541 0.054
R21405 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1493
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1492 0.054
R21406 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1438
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1437 0.054
R21407 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1389
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1388 0.054
R21408 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1334
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1333 0.054
R21409 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1753
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1752 0.054
R21410 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n577
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN 0.054
R21411 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n473
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/DRAIN 0.054
R21412 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n369
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN 0.054
R21413 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1618
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN 0.054
R21414 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1514
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN 0.054
R21415 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1410
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN 0.054
R21416 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1306
+ buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN 0.054
R21417 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1754 0.054
R21418 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n182
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n180 0.053
R21419 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n742
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n741 0.053
R21420 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1303
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1256 0.052
R21421 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1117
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1070 0.052
R21422 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n280
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n279 0.052
R21423 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n805
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n804 0.052
R21424 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n694
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n691 0.052
R21425 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n877
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n874 0.052
R21426 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n757
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n754 0.052
R21427 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n199
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n196 0.052
R21428 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1192
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1189 0.052
R21429 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1004
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1001 0.052
R21430 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1179
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1178 0.052
R21431 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n991
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n990 0.052
R21432 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n865
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n862 0.052
R21433 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n233
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n230 0.052
R21434 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1265
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1262 0.052
R21435 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1131
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1128 0.052
R21436 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1079
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1076 0.052
R21437 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n943
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n940 0.052
R21438 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n723
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n722 0.049
R21439 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n832
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n831 0.049
R21440 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n261
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n260 0.049
R21441 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n786
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n785 0.049
R21442 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1295
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1294 0.049
R21443 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1234
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1233 0.049
R21444 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1161
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1160 0.049
R21445 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1109
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1108 0.049
R21446 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1046
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1045 0.049
R21447 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n973
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n972 0.049
R21448 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n307
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n305 0.049
R21449 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n669
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n672 0.049
R21450 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n565
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n568 0.049
R21451 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n461
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n464 0.049
R21452 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1710
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1713 0.049
R21453 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1606
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1609 0.049
R21454 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1502
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1505 0.049
R21455 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1398
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1401 0.049
R21456 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n366
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n364 0.048
R21457 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n682
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n744 0.048
R21458 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n681
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n840 0.048
R21459 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n722
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n721 0.046
R21460 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n831
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n830 0.046
R21461 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n260
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n259 0.046
R21462 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n785
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n784 0.046
R21463 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1294
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1293 0.046
R21464 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1233
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1232 0.046
R21465 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1160
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1159 0.046
R21466 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1108
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1107 0.046
R21467 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1045
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1044 0.046
R21468 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n972
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n971 0.046
R21469 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n700
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n699 0.046
R21470 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n856
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n855 0.046
R21471 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n239
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n238 0.046
R21472 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n764
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n763 0.046
R21473 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1272
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1271 0.046
R21474 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1138
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1137 0.046
R21475 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1086
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1085 0.046
R21476 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n950
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n949 0.046
R21477 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n190
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n177 0.046
R21478 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n928
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n915 0.046
R21479 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1242
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1241 0.046
R21480 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1054
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1053 0.046
R21481 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n39
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n339 0.043
R21482 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n41
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1736 0.043
R21483 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n50
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n349 0.04
R21484 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n52
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1745 0.04
R21485 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n54
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n652 0.04
R21486 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n56
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n597 0.04
R21487 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n58
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n548 0.04
R21488 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n60
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n493 0.04
R21489 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n62
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n444 0.04
R21490 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n64
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n389 0.04
R21491 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n90
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1693 0.04
R21492 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n92
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1638 0.04
R21493 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n94
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1589 0.04
R21494 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n96
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1534 0.04
R21495 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n98
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1485 0.04
R21496 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n100
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1430 0.04
R21497 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n102
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1381 0.04
R21498 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n104
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1326 0.04
R21499 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1198
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1197 0.039
R21500 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1010
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1009 0.039
R21501 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n882
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n881 0.038
R21502 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n204
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n203 0.038
R21503 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n639
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n638 0.036
R21504 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n585
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n584 0.036
R21505 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n535
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n534 0.036
R21506 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n481
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n480 0.036
R21507 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n431
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n430 0.036
R21508 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n377
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n376 0.036
R21509 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n811
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n809 0.036
R21510 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n797
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n795 0.036
R21511 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n272
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n270 0.036
R21512 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1206
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1205 0.036
R21513 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1249
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1248 0.036
R21514 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1174
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1173 0.036
R21515 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1018
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1017 0.036
R21516 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1063
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1062 0.036
R21517 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n986
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n985 0.036
R21518 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1680
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1679 0.036
R21519 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1626
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1625 0.036
R21520 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1576
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1575 0.036
R21521 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1522
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1521 0.036
R21522 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1472
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1471 0.036
R21523 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1418
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1417 0.036
R21524 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1368
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1367 0.036
R21525 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1314
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1313 0.036
R21526 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n334
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n333 0.036
R21527 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1728
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1726 0.036
R21528 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n920
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n918 0.036
R21529 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n734
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n732 0.036
R21530 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n699
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n698 0.034
R21531 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n842
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n856 0.034
R21532 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n238
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n237 0.034
R21533 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n763
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n762 0.034
R21534 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1271
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1270 0.034
R21535 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1137
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1136 0.034
R21536 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1085
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1084 0.034
R21537 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n949
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n948 0.034
R21538 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n819
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n818 0.033
R21539 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n909
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n908 0.033
R21540 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n171
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n170 0.033
R21541 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n683
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE 0.032
R21542 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n806
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE 0.032
R21543 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1304
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE 0.032
R21544 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1118
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE 0.032
R21545 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n127
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n682 0.031
R21546 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n130
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1058 0.031
R21547 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n66
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n67 0.031
R21548 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n905
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n903 0.031
R21549 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n890
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n887 0.031
R21550 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n68
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n69 0.031
R21551 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n719
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n717 0.031
R21552 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n703
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n700 0.031
R21553 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n70
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n71 0.031
R21554 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n828
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n826 0.031
R21555 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n855
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n854 0.031
R21556 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n72
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n73 0.031
R21557 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n257
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n255 0.031
R21558 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n242
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n239 0.031
R21559 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n74
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n75 0.031
R21560 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n167
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n165 0.031
R21561 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n153
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n150 0.031
R21562 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n76
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n77 0.031
R21563 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n782
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n780 0.031
R21564 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n767
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n764 0.031
R21565 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1275
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1272 0.031
R21566 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1291
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1289 0.031
R21567 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n79
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n78 0.031
R21568 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1214
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1211 0.031
R21569 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1230
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1228 0.031
R21570 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n81
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n80 0.031
R21571 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1141
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1138 0.031
R21572 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1157
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1155 0.031
R21573 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n83
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n82 0.031
R21574 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1089
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1086 0.031
R21575 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1105
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1103 0.031
R21576 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n85
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n84 0.031
R21577 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1026
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1023 0.031
R21578 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1042
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1040 0.031
R21579 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n87
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n86 0.031
R21580 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n953
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n950 0.031
R21581 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n969
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n967 0.031
R21582 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n89
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n88 0.031
R21583 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n843
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n884 0.031
R21584 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1122
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1183 0.031
R21585 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n934
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n995 0.031
R21586 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n672
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n671 0.03
R21587 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n568
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n567 0.03
R21588 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n464
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n463 0.03
R21589 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1713
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1712 0.03
R21590 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1609
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1608 0.03
R21591 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1505
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1504 0.03
R21592 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1401
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1400 0.03
R21593 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n366
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n365 0.03
R21594 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n305
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n304 0.03
R21595 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n313
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n310 0.029
R21596 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n301
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n298 0.029
R21597 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n678
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n675 0.029
R21598 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n574
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n571 0.029
R21599 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n470
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n467 0.029
R21600 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1719
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1716 0.029
R21601 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1615
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1612 0.029
R21602 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1511
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1508 0.029
R21603 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1407
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1404 0.029
R21604 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n873
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n110 0.028
R21605 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n861
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n112 0.028
R21606 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n229
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n114 0.028
R21607 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n195
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n116 0.028
R21608 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n753
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n118 0.028
R21609 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n2
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n367 0.027
R21610 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n123
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n206 0.026
R21611 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n207
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n124 0.026
R21612 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n208
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n106 0.026
R21613 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n209
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n107 0.026
R21614 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n210
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n108 0.026
R21615 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n901
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n898 0.026
R21616 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n880
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n878 0.026
R21617 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n715
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n712 0.026
R21618 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n712
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n711 0.026
R21619 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n697
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n695 0.026
R21620 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n824
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n821 0.026
R21621 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n868
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n866 0.026
R21622 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n253
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n250 0.026
R21623 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n250
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n249 0.026
R21624 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n236
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n234 0.026
R21625 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n164
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n161 0.026
R21626 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n202
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n200 0.026
R21627 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n779
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n776 0.026
R21628 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n776
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n775 0.026
R21629 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n761
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n759 0.026
R21630 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1269
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1267 0.026
R21631 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1284
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1283 0.026
R21632 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1287
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1284 0.026
R21633 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1196
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1194 0.026
R21634 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1226
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1223 0.026
R21635 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1135
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1133 0.026
R21636 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1150
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1149 0.026
R21637 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1153
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1150 0.026
R21638 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1083
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1081 0.026
R21639 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1098
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1097 0.026
R21640 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1101
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1098 0.026
R21641 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1008
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1006 0.026
R21642 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1038
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1035 0.026
R21643 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n947
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n945 0.026
R21644 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n962
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n961 0.026
R21645 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n965
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n962 0.026
R21646 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n211
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n119 0.026
R21647 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n212
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n120 0.026
R21648 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n213
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n121 0.026
R21649 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n214
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n122 0.026
R21650 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n345
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n40 0.026
R21651 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1741
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n42 0.026
R21652 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n648
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n14 0.026
R21653 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n544
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n18 0.026
R21654 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n440
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n22 0.026
R21655 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1689
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n26 0.026
R21656 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1585
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n30 0.026
R21657 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1481
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n34 0.026
R21658 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1377
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n38 0.026
R21659 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n743
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n745 0.024
R21660 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n839
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n841 0.024
R21661 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n931
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n932 0.024
R21662 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1119
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1120 0.024
R21663 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n325
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n323 0.024
R21664 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n293
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n295 0.024
R21665 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n661
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n663 0.024
R21666 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n619
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n621 0.024
R21667 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n557
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n559 0.024
R21668 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n515
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n517 0.024
R21669 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n453
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n455 0.024
R21670 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n411
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n413 0.024
R21671 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n690
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n688 0.024
R21672 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1261
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1259 0.024
R21673 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1188
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1186 0.024
R21674 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1127
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1125 0.024
R21675 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1075
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1073 0.024
R21676 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1000
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n998 0.024
R21677 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n939
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n937 0.024
R21678 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1702
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1704 0.024
R21679 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1660
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1662 0.024
R21680 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1598
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1600 0.024
R21681 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1556
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1558 0.024
R21682 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1494
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1496 0.024
R21683 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1452
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1454 0.024
R21684 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1390
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1392 0.024
R21685 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1348
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1350 0.024
R21686 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n310
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n309 0.022
R21687 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n298
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n297 0.022
R21688 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n675
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n674 0.022
R21689 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n607
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n606 0.022
R21690 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n571
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n570 0.022
R21691 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n503
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n502 0.022
R21692 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n467
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n466 0.022
R21693 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n399
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n398 0.022
R21694 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1716
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1715 0.022
R21695 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1648
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1647 0.022
R21696 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1612
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1611 0.022
R21697 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1544
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1543 0.022
R21698 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1508
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1507 0.022
R21699 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1440
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1439 0.022
R21700 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1404
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1403 0.022
R21701 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1336
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1335 0.022
R21702 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n747
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n746 0.022
R21703 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n930
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n929 0.022
R21704 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1056
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1055 0.022
R21705 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1244
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1243 0.022
R21706 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n338
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n337 0.021
R21707 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1735
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1731 0.021
R21708 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n643
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n642 0.021
R21709 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n589
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n588 0.021
R21710 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n539
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n538 0.021
R21711 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n485
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n484 0.021
R21712 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n435
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n434 0.021
R21713 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n381
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n380 0.021
R21714 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n927
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n923 0.021
R21715 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n741
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n737 0.021
R21716 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n818
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n814 0.021
R21717 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n279
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n275 0.021
R21718 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n189
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n185 0.021
R21719 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n804
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n800 0.021
R21720 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1256
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1252 0.021
R21721 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1210
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1209 0.021
R21722 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1178
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1177 0.021
R21723 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1070
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1066 0.021
R21724 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1022
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1021 0.021
R21725 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n990
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n989 0.021
R21726 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1684
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1683 0.021
R21727 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1630
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1629 0.021
R21728 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1580
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1579 0.021
R21729 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1526
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1525 0.021
R21730 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1476
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1475 0.021
R21731 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1422
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1421 0.021
R21732 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1372
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1371 0.021
R21733 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1318
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1317 0.021
R21734 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n337
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n336 0.019
R21735 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1731
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1730 0.019
R21736 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n642
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n641 0.019
R21737 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n588
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n587 0.019
R21738 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n538
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n537 0.019
R21739 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n484
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n483 0.019
R21740 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n434
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n433 0.019
R21741 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n380
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n379 0.019
R21742 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n923
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n922 0.019
R21743 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n737
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n736 0.019
R21744 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n814
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n813 0.019
R21745 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n275
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n274 0.019
R21746 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n185
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n184 0.019
R21747 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n800
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n799 0.019
R21748 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1252
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1251 0.019
R21749 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1209
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1208 0.019
R21750 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1177
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1176 0.019
R21751 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1066
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1065 0.019
R21752 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1021
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1020 0.019
R21753 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n989
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n988 0.019
R21754 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1683
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1682 0.019
R21755 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1629
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1628 0.019
R21756 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1579
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1578 0.019
R21757 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1525
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1524 0.019
R21758 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1475
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1474 0.019
R21759 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1421
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1420 0.019
R21760 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1371
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1370 0.019
R21761 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1317
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1316 0.019
R21762 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n326
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n322 0.018
R21763 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n294
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n292 0.018
R21764 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n308
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n303 0.018
R21765 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n662
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n668 0.018
R21766 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n670
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n680 0.018
R21767 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n613
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n612 0.018
R21768 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n620
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n618 0.018
R21769 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n558
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n564 0.018
R21770 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n566
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n576 0.018
R21771 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n509
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n508 0.018
R21772 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n516
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n514 0.018
R21773 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n454
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n460 0.018
R21774 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n462
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n472 0.018
R21775 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n405
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n404 0.018
R21776 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n412
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n410 0.018
R21777 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1703
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1709 0.018
R21778 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1711
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1721 0.018
R21779 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1654
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1653 0.018
R21780 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1661
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1659 0.018
R21781 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1599
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1605 0.018
R21782 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1607
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1617 0.018
R21783 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1550
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1549 0.018
R21784 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1557
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1555 0.018
R21785 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1495
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1501 0.018
R21786 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1503
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1513 0.018
R21787 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1446
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1445 0.018
R21788 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1453
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1451 0.018
R21789 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1391
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1397 0.018
R21790 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1399
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1409 0.018
R21791 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1342
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1341 0.018
R21792 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1349
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1347 0.018
R21793 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n317
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n315 0.018
R21794 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n894
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n892 0.017
R21795 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n708
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n706 0.017
R21796 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n849
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n848 0.017
R21797 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n246
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n244 0.017
R21798 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n157
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n155 0.017
R21799 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n772
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n770 0.017
R21800 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1280
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1278 0.017
R21801 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1219
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1217 0.017
R21802 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1146
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1144 0.017
R21803 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1094
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1092 0.017
R21804 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1031
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1029 0.017
R21805 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n958
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n956 0.017
R21806 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n349
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n348 0.016
R21807 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1745
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1744 0.016
R21808 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n652
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n651 0.016
R21809 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n597
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n596 0.016
R21810 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n548
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n547 0.016
R21811 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n493
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n492 0.016
R21812 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n444
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n443 0.016
R21813 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n389
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n388 0.016
R21814 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1693
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1692 0.016
R21815 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1638
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1637 0.016
R21816 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1589
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1588 0.016
R21817 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1534
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1533 0.016
R21818 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1485
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1484 0.016
R21819 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1430
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1429 0.016
R21820 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1381
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1380 0.016
R21821 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1326
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1325 0.016
R21822 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n368
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1723 0.015
R21823 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n294
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n293 0.014
R21824 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n326
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n325 0.014
R21825 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n412
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n411 0.014
R21826 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n454
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n453 0.014
R21827 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n516
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n515 0.014
R21828 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n558
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n557 0.014
R21829 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n620
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n619 0.014
R21830 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n662
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n661 0.014
R21831 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1349
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1348 0.014
R21832 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1391
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1390 0.014
R21833 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1453
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1452 0.014
R21834 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1495
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1494 0.014
R21835 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1557
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1556 0.014
R21836 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1599
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1598 0.014
R21837 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1661
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1660 0.014
R21838 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1703
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1702 0.014
R21839 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n315
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n313 0.014
R21840 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n336
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n334 0.014
R21841 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n303
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n301 0.014
R21842 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1730
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1728 0.014
R21843 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n680
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n678 0.014
R21844 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n641
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n639 0.014
R21845 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n612
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n610 0.014
R21846 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n587
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n585 0.014
R21847 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n576
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n574 0.014
R21848 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n537
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n535 0.014
R21849 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n508
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n506 0.014
R21850 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n483
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n481 0.014
R21851 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n472
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n470 0.014
R21852 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n433
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n431 0.014
R21853 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n404
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n402 0.014
R21854 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n379
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n377 0.014
R21855 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n922
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n920 0.014
R21856 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n896
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n894 0.014
R21857 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n891
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n890 0.014
R21858 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n881
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n880 0.014
R21859 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n878
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n877 0.014
R21860 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n736
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n734 0.014
R21861 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n710
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n708 0.014
R21862 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n705
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n703 0.014
R21863 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n698
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n697 0.014
R21864 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n695
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n694 0.014
R21865 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n813
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n811 0.014
R21866 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n848
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n846 0.014
R21867 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n854
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n851 0.014
R21868 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n842
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n868 0.014
R21869 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n866
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n865 0.014
R21870 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n274
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n272 0.014
R21871 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n248
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n246 0.014
R21872 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n243
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n242 0.014
R21873 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n237
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n236 0.014
R21874 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n234
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n233 0.014
R21875 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n184
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n182 0.014
R21876 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n159
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n157 0.014
R21877 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n154
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n153 0.014
R21878 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n203
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n202 0.014
R21879 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n200
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n199 0.014
R21880 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n799
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n797 0.014
R21881 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n774
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n772 0.014
R21882 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n769
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n767 0.014
R21883 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n762
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n761 0.014
R21884 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n759
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n757 0.014
R21885 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1267
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1265 0.014
R21886 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1270
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1269 0.014
R21887 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1277
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1275 0.014
R21888 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1282
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1280 0.014
R21889 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1251
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1249 0.014
R21890 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1194
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1192 0.014
R21891 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1197
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1196 0.014
R21892 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1216
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1214 0.014
R21893 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1221
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1219 0.014
R21894 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1208
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1206 0.014
R21895 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1133
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1131 0.014
R21896 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1136
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1135 0.014
R21897 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1143
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1141 0.014
R21898 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1148
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1146 0.014
R21899 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1176
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1174 0.014
R21900 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1081
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1079 0.014
R21901 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1084
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1083 0.014
R21902 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1091
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1089 0.014
R21903 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1096
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1094 0.014
R21904 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1065
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1063 0.014
R21905 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1006
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1004 0.014
R21906 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1009
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1008 0.014
R21907 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1028
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1026 0.014
R21908 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1033
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1031 0.014
R21909 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1020
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1018 0.014
R21910 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n945
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n943 0.014
R21911 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n948
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n947 0.014
R21912 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n955
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n953 0.014
R21913 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n960
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n958 0.014
R21914 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n988
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n986 0.014
R21915 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1721
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1719 0.014
R21916 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1682
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1680 0.014
R21917 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1653
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1651 0.014
R21918 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1628
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1626 0.014
R21919 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1617
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1615 0.014
R21920 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1578
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1576 0.014
R21921 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1549
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1547 0.014
R21922 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1524
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1522 0.014
R21923 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1513
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1511 0.014
R21924 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1474
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1472 0.014
R21925 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1445
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1443 0.014
R21926 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1420
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1418 0.014
R21927 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1409
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1407 0.014
R21928 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1370
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1368 0.014
R21929 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1341
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1339 0.014
R21930 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1316
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1314 0.014
R21931 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n898
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n897 0.013
R21932 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n161
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n160 0.013
R21933 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1223
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1222 0.013
R21934 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1035
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1034 0.013
R21935 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n367
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n222 0.011
R21936 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n884
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n883 0.011
R21937 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1183
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1182 0.011
R21938 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n995
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n994 0.011
R21939 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1754
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3 0.01
R21940 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n308
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n307 0.009
R21941 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n317
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n316 0.009
R21942 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n405
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n406 9.309
R21943 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n462
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n461 0.009
R21944 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n509
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n510 9.309
R21945 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n566
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n565 0.009
R21946 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n613
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n614 9.309
R21947 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n670
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n669 0.009
R21948 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1342
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1343 9.309
R21949 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1399
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1398 0.009
R21950 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1446
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1447 9.309
R21951 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1503
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1502 0.009
R21952 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1550
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1551 9.309
R21953 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1607
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1606 0.009
R21954 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1654
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1655 9.309
R21955 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1711
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1710 0.009
R21956 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n339
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n340 0.009
R21957 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n347
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n345 0.009
R21958 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1743
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1741 0.009
R21959 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n631
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n630 0.009
R21960 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n650
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n648 0.009
R21961 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n12
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n11 9.309
R21962 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n595
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n593 0.009
R21963 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n527
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n526 0.009
R21964 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n546
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n544 0.009
R21965 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n16
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n15 9.309
R21966 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n491
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n489 0.009
R21967 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n423
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n422 0.009
R21968 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n442
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n440 0.009
R21969 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n20
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n19 9.309
R21970 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n387
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n385 0.009
R21971 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n907
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n905 0.009
R21972 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n903
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n901 0.009
R21973 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n721
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n719 0.009
R21974 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n717
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n715 0.009
R21975 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n830
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n828 0.009
R21976 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n826
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n824 0.009
R21977 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n259
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n257 0.009
R21978 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n255
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n253 0.009
R21979 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n169
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n167 0.009
R21980 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n165
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n164 0.009
R21981 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n784
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n782 0.009
R21982 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n780
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n779 0.009
R21983 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1289
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1287 0.009
R21984 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1293
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1291 0.009
R21985 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1228
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1226 0.009
R21986 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1232
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1230 0.009
R21987 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1155
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1153 0.009
R21988 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1159
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1157 0.009
R21989 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1103
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1101 0.009
R21990 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1107
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1105 0.009
R21991 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1040
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1038 0.009
R21992 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1044
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1042 0.009
R21993 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n967
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n965 0.009
R21994 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n971
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n969 0.009
R21995 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1672
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1671 0.009
R21996 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1691
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1689 0.009
R21997 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n24
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n23 9.309
R21998 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1636
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1634 0.009
R21999 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1568
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1567 0.009
R22000 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1587
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1585 0.009
R22001 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n28
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n27 9.309
R22002 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1532
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1530 0.009
R22003 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1464
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1463 0.009
R22004 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1483
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1481 0.009
R22005 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n32
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n31 9.309
R22006 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1428
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1426 0.009
R22007 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1360
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1359 0.009
R22008 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1379
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1377 0.009
R22009 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n36
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n35 9.309
R22010 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n105
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n104 0.035
R22011 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n103
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n102 0.035
R22012 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n101
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n100 0.035
R22013 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n99
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n98 0.035
R22014 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n97
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n96 0.035
R22015 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n95
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n94 0.035
R22016 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n93
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n92 0.035
R22017 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n91
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n90 0.035
R22018 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n65
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n64 0.035
R22019 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n63
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n62 0.035
R22020 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n61
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n60 0.035
R22021 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n59
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n58 0.035
R22022 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n57
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n56 0.035
R22023 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n55
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n54 0.035
R22024 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n53
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n52 0.035
R22025 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n51
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n50 0.035
R22026 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1057
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n130 0.026
R22027 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n681
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n127 0.026
R22028 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n88
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n973 0.025
R22029 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n86
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1046 0.025
R22030 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n84
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1109 0.025
R22031 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n82
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1161 0.025
R22032 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n80
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1234 0.025
R22033 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n78
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1295 0.025
R22034 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n77
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n786 0.025
R22035 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n75
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n171 0.025
R22036 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n73
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n261 0.025
R22037 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n71
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n832 0.025
R22038 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n69
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n723 0.025
R22039 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n67
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n909 0.025
R22040 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1333
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n105 0.023
R22041 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1388
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n103 0.023
R22042 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1437
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n101 0.023
R22043 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1492
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n99 0.023
R22044 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1541
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n97 0.023
R22045 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1596
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n95 0.023
R22046 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1645
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n93 0.023
R22047 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1700
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n91 0.023
R22048 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n993
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n89 0.023
R22049 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1053
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n87 0.023
R22050 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1116
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n85 0.023
R22051 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1181
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n83 0.023
R22052 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1241
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n81 0.023
R22053 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1302
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n79 0.023
R22054 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n792
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n76 0.023
R22055 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n177
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n74 0.023
R22056 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n267
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n72 0.023
R22057 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n838
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n70 0.023
R22058 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n729
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n68 0.023
R22059 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n915
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n66 0.023
R22060 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n396
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n65 0.023
R22061 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n451
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n63 0.023
R22062 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n500
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n61 0.023
R22063 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n555
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n59 0.023
R22064 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n604
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n57 0.023
R22065 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n659
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n55 0.023
R22066 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1752
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n53 0.023
R22067 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n356
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n51 0.023
R22068 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n124
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n283 0.015
R22069 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n364
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n123 0.015
R22070 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n122
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1354 0.015
R22071 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n121
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1458 0.015
R22072 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n120
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1562 0.015
R22073 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n119
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1666 0.015
R22074 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n108
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n417 0.015
R22075 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n107
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n521 0.015
R22076 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n106
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n625 0.015
R22077 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1358
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n214 0.014
R22078 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1462
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n213 0.014
R22079 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1566
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n212 0.014
R22080 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1670
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n211 0.014
R22081 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n421
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n210 0.014
R22082 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n525
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n209 0.014
R22083 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n629
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n208 0.014
R22084 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n207
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n288 0.014
R22085 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n206
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n359 0.014
R22086 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n129
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1118 0.013
R22087 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n128
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1304 0.013
R22088 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n126
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n806 0.013
R22089 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n125
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n683 0.013
R22090 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n118
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n117 0.013
R22091 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n116
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n115 0.013
R22092 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n114
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n113 0.013
R22093 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n112
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n111 0.013
R22094 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n110
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n109 0.013
R22095 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1324
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1322 0.009
R22096 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n851
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n849 0.008
R22097 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n706
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n705 0.008
R22098 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n892
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n891 0.008
R22099 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n244
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n243 0.008
R22100 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n770
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n769 0.008
R22101 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n155
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n154 0.008
R22102 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1278
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1277 0.008
R22103 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1217
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1216 0.008
R22104 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1144
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1143 0.008
R22105 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1092
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1091 0.008
R22106 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1029
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1028 0.008
R22107 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n956
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n955 0.008
R22108 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n934
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n933 0.008
R22109 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1122
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1121 0.008
R22110 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n146
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n144 0.008
R22111 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n143
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n142 0.008
R22112 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n141
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n140 0.008
R22113 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n139
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n137 0.008
R22114 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n136
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n135 0.008
R22115 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n134
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n133 0.008
R22116 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n132
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n131 0.008
R22117 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n322
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n320 0.006
R22118 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n292
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n290 0.006
R22119 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n668
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n666 0.006
R22120 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n618
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n616 0.006
R22121 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n564
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n562 0.006
R22122 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n514
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n512 0.006
R22123 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n460
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n458 0.006
R22124 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n410
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n408 0.006
R22125 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1709
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1707 0.006
R22126 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1659
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1657 0.006
R22127 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1605
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1603 0.006
R22128 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1555
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1553 0.006
R22129 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1501
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1499 0.006
R22130 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1451
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1449 0.006
R22131 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1397
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1395 0.006
R22132 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1347
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1345 0.006
R22133 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n146
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n145 0.006
R22134 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n139
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n138 0.006
R22135 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n744
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n743 0.005
R22136 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n840
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n839 0.005
R22137 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1057
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n931 0.053
R22138 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1058
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1119 0.053
R22139 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1322
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n36 0.031
R22140 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1426
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n32 0.031
R22141 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1530
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n28 0.031
R22142 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1634
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n24 0.031
R22143 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n385
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n20 0.031
R22144 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n489
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n16 0.031
R22145 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n593
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n12 0.031
R22146 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n577 0.015
R22147 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n473 0.015
R22148 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n369 0.015
R22149 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1618 0.015
R22150 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1514 0.015
R22151 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1410 0.015
R22152 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1306 0.015
R22153 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n0 0.014
R22154 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n42
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n41 0.014
R22155 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n40
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n39 0.014
R22156 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n38
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n37 0.014
R22157 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n34
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n33 0.014
R22158 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n30
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n29 0.014
R22159 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n26
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n25 0.014
R22160 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n22
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n21 0.014
R22161 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n18
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n17 0.014
R22162 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n14
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n13 0.014
R22163 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n2 0.012
R22164 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n937
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n49 0.012
R22165 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n998
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n48 0.012
R22166 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1073
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n47 0.012
R22167 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1125
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n46 0.012
R22168 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1186
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n45 0.012
R22169 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1259
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n44 0.012
R22170 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n688
+ buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n43 0.012
R22171 IN_N.n277 IN_N.t6 846.712
R22172 IN_N.n258 IN_N.t3 846.712
R22173 IN_N.n17 IN_N.t2 846.712
R22174 IN_N.n292 IN_N.t0 846.712
R22175 IN_N.n373 IN_N.t5 846.712
R22176 IN_N.n326 IN_N.t7 846.712
R22177 IN_N.n2 IN_N.t4 846.712
R22178 IN_N.n362 IN_N.t1 846.712
R22179 IN_N.n150 IN_N.n148 15.887
R22180 IN_N.n293 IN_N.n292 15.887
R22181 IN_N.n18 IN_N.n17 15.887
R22182 IN_N.n52 IN_N.n51 15.887
R22183 IN_N.n3 IN_N.n2 15.887
R22184 IN_N.n363 IN_N.n362 15.887
R22185 IN_N.n160 IN_N.n159 12.054
R22186 IN_N.n62 IN_N.n61 12.054
R22187 IN_N.n182 IN_N.n181 10.328
R22188 IN_N.n205 IN_N.n204 10.328
R22189 IN_N.n279 IN_N.n278 10.328
R22190 IN_N.n260 IN_N.n259 10.328
R22191 IN_N.n84 IN_N.n83 10.328
R22192 IN_N.n107 IN_N.n106 10.328
R22193 IN_N.n328 IN_N.n327 10.328
R22194 IN_N.n375 IN_N.n374 10.328
R22195 IN_N.n174 IN_N.n173 9.3
R22196 IN_N.n185 IN_N.n184 9.3
R22197 IN_N.n184 IN_N.n183 9.3
R22198 IN_N.n207 IN_N.n206 9.3
R22199 IN_N.n287 IN_N.n286 9.3
R22200 IN_N.n263 IN_N.n262 9.3
R22201 IN_N.n262 IN_N.n261 9.3
R22202 IN_N.n252 IN_N.n14 9.3
R22203 IN_N.n282 IN_N.n281 9.3
R22204 IN_N.n281 IN_N.n280 9.3
R22205 IN_N.n76 IN_N.n75 9.3
R22206 IN_N.n109 IN_N.n108 9.3
R22207 IN_N.n87 IN_N.n86 9.3
R22208 IN_N.n86 IN_N.n85 9.3
R22209 IN_N.n320 IN_N.n319 9.3
R22210 IN_N.n331 IN_N.n330 9.3
R22211 IN_N.n330 IN_N.n329 9.3
R22212 IN_N.n378 IN_N.n377 9.3
R22213 IN_N.n377 IN_N.n376 9.3
R22214 IN_N.n367 IN_N.n341 9.3
R22215 IN_N.n177 IN_N.n176 9
R22216 IN_N.n255 IN_N.n254 9
R22217 IN_N.n284 IN_N.n283 9
R22218 IN_N.n79 IN_N.n78 9
R22219 IN_N.n370 IN_N.n369 9
R22220 IN_N.n323 IN_N.n322 9
R22221 IN_N.n192 IN_N.n191 8.764
R22222 IN_N.n270 IN_N.n269 8.764
R22223 IN_N.n94 IN_N.n93 8.764
R22224 IN_N.n336 IN_N.n335 8.764
R22225 IN_N.n181 IN_N.n180 6.885
R22226 IN_N.n204 IN_N.n203 6.885
R22227 IN_N.n278 IN_N.n277 6.885
R22228 IN_N.n259 IN_N.n258 6.885
R22229 IN_N.n83 IN_N.n82 6.885
R22230 IN_N.n106 IN_N.n105 6.885
R22231 IN_N.n327 IN_N.n326 6.885
R22232 IN_N.n374 IN_N.n373 6.885
R22233 IN_N.n150 IN_N.n149 6.276
R22234 IN_N.n293 IN_N.n290 6.276
R22235 IN_N.n18 IN_N.n15 6.276
R22236 IN_N.n52 IN_N.n49 6.276
R22237 IN_N.n3 IN_N.n0 6.276
R22238 IN_N.n363 IN_N.n360 6.276
R22239 IN_N.n179 IN_N.n178 5.647
R22240 IN_N.n202 IN_N.n201 5.647
R22241 IN_N.n276 IN_N.n275 5.647
R22242 IN_N.n257 IN_N.n256 5.647
R22243 IN_N.n81 IN_N.n80 5.647
R22244 IN_N.n104 IN_N.n103 5.647
R22245 IN_N.n325 IN_N.n324 5.647
R22246 IN_N.n372 IN_N.n371 5.647
R22247 IN_N.n161 IN_N.n160 4.934
R22248 IN_N.n63 IN_N.n62 4.934
R22249 IN_N.n155 IN_N.n154 4.894
R22250 IN_N.n57 IN_N.n56 4.894
R22251 IN_N.n159 IN_N.n158 4.82
R22252 IN_N.n61 IN_N.n60 4.82
R22253 IN_N.n199 IN_N.n198 4.65
R22254 IN_N.n101 IN_N.n100 4.65
R22255 IN_N.n193 IN_N.n192 4.574
R22256 IN_N.n208 IN_N.n207 4.574
R22257 IN_N.n271 IN_N.n270 4.574
R22258 IN_N.n110 IN_N.n109 4.574
R22259 IN_N.n95 IN_N.n94 4.574
R22260 IN_N.n337 IN_N.n336 4.574
R22261 IN_N.n148 IN_N.n147 4.131
R22262 IN_N.n158 IN_N.n157 4.131
R22263 IN_N.n292 IN_N.n291 4.131
R22264 IN_N.n17 IN_N.n16 4.131
R22265 IN_N.n51 IN_N.n50 4.131
R22266 IN_N.n60 IN_N.n59 4.131
R22267 IN_N.n2 IN_N.n1 4.131
R22268 IN_N.n362 IN_N.n361 4.131
R22269 IN_N.n249 IN_N.n18 4.11
R22270 IN_N.n364 IN_N.n363 4.109
R22271 IN_N.n294 IN_N.n293 4.109
R22272 IN_N.n316 IN_N.n3 4.109
R22273 IN_N.n151 IN_N.n150 3.737
R22274 IN_N.n53 IN_N.n52 3.737
R22275 IN_N.n146 IN_N.n145 3.544
R22276 IN_N.n164 IN_N.n163 3
R22277 IN_N.n210 IN_N.n209 3
R22278 IN_N.n66 IN_N.n65 3
R22279 IN_N.n112 IN_N.n111 3
R22280 IN_N.n244 IN_N.n243 2.73
R22281 IN_N.n183 IN_N.n182 1.377
R22282 IN_N.n206 IN_N.n205 1.377
R22283 IN_N.n280 IN_N.n279 1.377
R22284 IN_N.n261 IN_N.n260 1.377
R22285 IN_N.n85 IN_N.n84 1.377
R22286 IN_N.n108 IN_N.n107 1.377
R22287 IN_N.n329 IN_N.n328 1.377
R22288 IN_N.n376 IN_N.n375 1.377
R22289 IN_N.n316 IN_N.n315 1.19
R22290 IN_N.n364 IN_N.n359 1.185
R22291 IN_N.n295 IN_N.n294 1.185
R22292 IN_N.n249 IN_N.n248 1.185
R22293 IN_N.n231 IN_N.n151 1.181
R22294 IN_N.n133 IN_N.n53 1.181
R22295 IN_N.n315 IN_N.n314 1.152
R22296 IN_N.n232 IN_N.n231 1.151
R22297 IN_N.n134 IN_N.n133 1.141
R22298 IN_N.n301 IN_N.n300 1.137
R22299 IN_N.n32 IN_N.n31 1.137
R22300 IN_N.n46 IN_N.n45 1.137
R22301 IN_N.n247 IN_N.n246 1.137
R22302 IN_N.n184 IN_N.n179 0.752
R22303 IN_N.n207 IN_N.n202 0.752
R22304 IN_N.n156 IN_N.n155 0.752
R22305 IN_N.n160 IN_N.n156 0.752
R22306 IN_N.n281 IN_N.n276 0.752
R22307 IN_N.n262 IN_N.n257 0.752
R22308 IN_N.n86 IN_N.n81 0.752
R22309 IN_N.n109 IN_N.n104 0.752
R22310 IN_N.n58 IN_N.n57 0.752
R22311 IN_N.n62 IN_N.n58 0.752
R22312 IN_N.n330 IN_N.n325 0.752
R22313 IN_N.n377 IN_N.n372 0.752
R22314 IN_N.n303 IN_N.n302 0.355
R22315 IN_N.n245 IN_N.n244 0.302
R22316 IN_N.n244 IN_N.n146 0.23
R22317 IN_N.n146 IN_N 0.072
R22318 IN_N.n289 IN_N.n288 0.054
R22319 IN_N.n273 IN_N.n272 0.054
R22320 IN_N.n318 IN_N.n317 0.054
R22321 IN_N.n334 IN_N.n333 0.054
R22322 IN_N.n251 IN_N.n250 0.051
R22323 IN_N.n366 IN_N.n365 0.051
R22324 IN_N.n172 IN_N.n171 0.047
R22325 IN_N.n74 IN_N.n73 0.047
R22326 IN_N.n188 IN_N.n187 0.045
R22327 IN_N.n90 IN_N.n89 0.045
R22328 IN_N.n317 IN_N.n316 0.039
R22329 IN_N.n294 IN_N.n289 0.039
R22330 IN_N.n267 IN_N.n266 0.039
R22331 IN_N.n340 IN_N.n339 0.039
R22332 IN_N.n250 IN_N.n249 0.038
R22333 IN_N.n365 IN_N.n364 0.038
R22334 IN_N.n347 IN_N.n346 0.038
R22335 IN_N IN_N.n195 0.037
R22336 IN_N.n272 IN_N.n271 0.037
R22337 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE IN_N.n97 0.037
R22338 IN_N.n337 IN_N.n334 0.037
R22339 IN_N.n314 IN_N.n313 0.037
R22340 IN_N.n21 IN_N.n13 0.037
R22341 IN_N.n298 IN_N.n297 0.036
R22342 IN_N.n29 IN_N.n28 0.036
R22343 IN_N.n11 IN_N.n10 0.036
R22344 IN_N.n344 IN_N.n343 0.036
R22345 IN_N.n306 IN_N.n305 0.035
R22346 IN_N.n48 IN_N.n47 0.035
R22347 IN_N.n171 IN_N.n151 0.035
R22348 IN_N.n73 IN_N.n53 0.035
R22349 IN_N.n190 IN_N.n189 0.034
R22350 IN_N.n92 IN_N.n91 0.034
R22351 IN_N.n266 IN_N 0.032
R22352 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE IN_N.n340 0.032
R22353 IN_N.n356 IN_N.n355 0.031
R22354 IN_N.n163 IN_N.n162 0.03
R22355 IN_N.n65 IN_N.n64 0.03
R22356 IN_N.n315 IN_N.n12 0.03
R22357 IN_N.n233 IN_N.n232 0.029
R22358 IN_N.n241 IN_N.n240 0.029
R22359 IN_N.n310 IN_N.n309 0.029
R22360 IN_N.n35 IN_N.n34 0.029
R22361 IN_N.n168 IN_N.n167 0.027
R22362 IN_N.n300 IN_N.n299 0.027
R22363 IN_N.n38 IN_N.n37 0.027
R22364 IN_N.n70 IN_N.n69 0.027
R22365 IN_N.n348 IN_N.n347 0.027
R22366 IN_N.n200 IN_N.n199 0.026
R22367 IN_N.n102 IN_N.n101 0.026
R22368 IN_N.n237 IN_N.n236 0.025
R22369 IN_N.n30 IN_N.n29 0.025
R22370 IN_N.n247 IN_N.n20 0.025
R22371 IN_N.n343 IN_N.n342 0.025
R22372 IN_N.n358 IN_N.n357 0.025
R22373 IN_N.n177 IN_N.n175 0.024
R22374 IN_N.n194 IN_N.n193 0.024
R22375 IN_N.n253 IN_N.n252 0.024
R22376 IN_N.n79 IN_N.n77 0.024
R22377 IN_N.n96 IN_N.n95 0.024
R22378 IN_N.n368 IN_N.n367 0.024
R22379 IN_N.n219 IN_N.n218 0.023
R22380 IN_N.n169 IN_N.n168 0.023
R22381 IN_N.n41 IN_N.n40 0.023
R22382 IN_N.n121 IN_N.n120 0.023
R22383 IN_N.n71 IN_N.n70 0.023
R22384 IN_N.n354 IN_N.n353 0.023
R22385 IN_N.n209 IN_N.n208 0.022
R22386 IN_N.n285 IN_N.n284 0.022
R22387 IN_N.n282 IN_N.n274 0.022
R22388 IN_N IN_N.n265 0.022
R22389 IN_N.n24 IN_N.n23 0.022
R22390 IN_N.n111 IN_N.n110 0.022
R22391 IN_N.n323 IN_N.n321 0.022
R22392 IN_N.n332 IN_N.n331 0.022
R22393 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE IN_N.n380 0.022
R22394 IN_N.n9 IN_N.n8 0.022
R22395 IN_N.n7 IN_N.n6 0.022
R22396 IN_N.n186 IN_N.n185 0.02
R22397 IN_N.n209 IN_N.n197 0.02
R22398 IN_N.n43 IN_N.n42 0.02
R22399 IN_N.n88 IN_N.n87 0.02
R22400 IN_N.n111 IN_N.n99 0.02
R22401 IN_N.n352 IN_N.n351 0.02
R22402 IN_N.n230 IN_N.n229 0.018
R22403 IN_N.n187 IN_N.n186 0.018
R22404 IN_N.n31 IN_N.n30 0.018
R22405 IN_N.n20 IN_N.n19 0.018
R22406 IN_N.n132 IN_N.n131 0.018
R22407 IN_N.n89 IN_N.n88 0.018
R22408 IN_N.n357 IN_N.n356 0.018
R22409 IN_N.n274 IN_N.n273 0.017
R22410 IN_N.n265 IN_N.n264 0.017
R22411 IN_N.n264 IN_N.n263 0.017
R22412 IN_N.n333 IN_N.n332 0.017
R22413 IN_N.n380 IN_N.n379 0.017
R22414 IN_N.n379 IN_N.n378 0.017
R22415 IN_N.n227 IN_N.n226 0.016
R22416 IN_N.n221 IN_N.n220 0.016
R22417 IN_N.n217 IN_N.n216 0.016
R22418 IN_N.n299 IN_N.n298 0.016
R22419 IN_N.n25 IN_N.n24 0.016
R22420 IN_N.n44 IN_N.n43 0.016
R22421 IN_N.n129 IN_N.n128 0.016
R22422 IN_N.n123 IN_N.n122 0.016
R22423 IN_N.n119 IN_N.n118 0.016
R22424 IN_N.n12 IN_N.n11 0.016
R22425 IN_N.n6 IN_N.n5 0.016
R22426 IN_N.n351 IN_N.n350 0.016
R22427 IN_N.n305 IN_N.n304 0.016
R22428 IN_N.n301 IN_N.n13 0.016
R22429 IN_N.n246 IN_N.n48 0.016
R22430 IN_N.n242 IN_N.n241 0.015
R22431 IN_N.n210 IN_N.n170 0.015
R22432 IN_N.n252 IN_N.n251 0.015
R22433 IN_N.n112 IN_N.n72 0.015
R22434 IN_N.n367 IN_N.n366 0.015
R22435 IN_N.n229 IN_N.n228 0.014
R22436 IN_N.n225 IN_N.n224 0.014
R22437 IN_N.n211 IN_N.n210 0.014
R22438 IN_N.n297 IN_N.n296 0.014
R22439 IN_N.n45 IN_N.n38 0.014
R22440 IN_N.n40 IN_N.n39 0.014
R22441 IN_N.n131 IN_N.n130 0.014
R22442 IN_N.n127 IN_N.n126 0.014
R22443 IN_N.n113 IN_N.n112 0.014
R22444 IN_N.n10 IN_N.n9 0.014
R22445 IN_N.n349 IN_N.n348 0.014
R22446 IN_N.n355 IN_N.n354 0.014
R22447 IN_N.n133 IN_N.n132 0.013
R22448 IN_N.n231 IN_N.n230 0.013
R22449 IN_N.n224 IN_N.n223 0.013
R22450 IN_N.n213 IN_N.n212 0.013
R22451 IN_N.n153 IN_N.n152 0.013
R22452 IN_N.n126 IN_N.n125 0.013
R22453 IN_N.n115 IN_N.n114 0.013
R22454 IN_N.n55 IN_N.n54 0.013
R22455 IN_N.n193 IN_N.n190 0.011
R22456 IN_N.n195 IN_N.n194 0.011
R22457 IN_N.n45 IN_N.n44 0.011
R22458 IN_N.n95 IN_N.n92 0.011
R22459 IN_N.n97 IN_N.n96 0.011
R22460 IN_N.n350 IN_N.n349 0.011
R22461 IN_N.n222 IN_N.n221 0.01
R22462 IN_N.n214 IN_N.n213 0.01
R22463 IN_N.n135 IN_N.n134 0.01
R22464 IN_N.n143 IN_N.n142 0.01
R22465 IN_N.n124 IN_N.n123 0.01
R22466 IN_N.n116 IN_N.n115 0.01
R22467 IN_N.n309 IN_N.n308 0.01
R22468 IN_N.n307 IN_N.n306 0.01
R22469 IN_N.n36 IN_N.n35 0.01
R22470 IN_N.n47 IN_N.n46 0.01
R22471 IN_N.n228 IN_N.n227 0.009
R22472 IN_N.n215 IN_N.n214 0.009
R22473 IN_N.n174 IN_N.n172 0.009
R22474 IN_N.n196 IN_N 0.009
R22475 IN_N.n288 IN_N.n287 0.009
R22476 IN_N.n31 IN_N.n25 0.009
R22477 IN_N.n130 IN_N.n129 0.009
R22478 IN_N.n117 IN_N.n116 0.009
R22479 IN_N.n76 IN_N.n74 0.009
R22480 IN_N.n98 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE 0.009
R22481 IN_N.n320 IN_N.n318 0.009
R22482 IN_N.n5 IN_N.n4 0.009
R22483 IN_N.n313 IN_N.n312 0.009
R22484 IN_N.n311 IN_N.n310 0.009
R22485 IN_N.n32 IN_N.n21 0.009
R22486 IN_N.n34 IN_N.n33 0.009
R22487 IN_N.n234 IN_N.n233 0.008
R22488 IN_N.n236 IN_N.n235 0.008
R22489 IN_N.n238 IN_N.n237 0.008
R22490 IN_N.n240 IN_N.n239 0.008
R22491 IN_N.n139 IN_N.n138 0.008
R22492 IN_N.n218 IN_N.n217 0.007
R22493 IN_N.n216 IN_N.n215 0.007
R22494 IN_N.n300 IN_N.n295 0.007
R22495 IN_N.n248 IN_N.n247 0.007
R22496 IN_N.n120 IN_N.n119 0.007
R22497 IN_N.n118 IN_N.n117 0.007
R22498 IN_N.n359 IN_N.n358 0.007
R22499 IN_N.n166 IN_N.n165 0.006
R22500 IN_N.n68 IN_N.n67 0.006
R22501 IN_N.n312 IN_N.n311 0.006
R22502 IN_N.n33 IN_N.n32 0.006
R22503 IN_N.n235 IN_N.n234 0.005
R22504 IN_N.n239 IN_N.n238 0.005
R22505 IN_N.n197 IN_N.n196 0.005
R22506 IN_N.n208 IN_N.n200 0.005
R22507 IN_N.n163 IN_N.n153 0.005
R22508 IN_N.n287 IN_N.n285 0.005
R22509 IN_N.n144 IN_N.n143 0.005
R22510 IN_N.n99 IN_N.n98 0.005
R22511 IN_N.n110 IN_N.n102 0.005
R22512 IN_N.n65 IN_N.n55 0.005
R22513 IN_N.n321 IN_N.n320 0.005
R22514 IN_N.n308 IN_N.n307 0.005
R22515 IN_N.n46 IN_N.n36 0.005
R22516 IN_N.n162 IN_N.n161 0.004
R22517 IN_N.n64 IN_N.n63 0.004
R22518 IN_N.n243 IN_N.n242 0.003
R22519 IN_N.n223 IN_N.n222 0.003
R22520 IN_N.n212 IN_N.n211 0.003
R22521 IN_N.n170 IN_N.n169 0.003
R22522 IN_N.n165 IN_N.n164 0.003
R22523 IN_N.n175 IN_N.n174 0.003
R22524 IN_N.n185 IN_N.n177 0.003
R22525 IN_N.n284 IN_N.n282 0.003
R22526 IN_N.n263 IN_N.n255 0.003
R22527 IN_N.n255 IN_N.n253 0.003
R22528 IN_N.n23 IN_N.n22 0.003
R22529 IN_N.n42 IN_N.n41 0.003
R22530 IN_N.n136 IN_N.n135 0.003
R22531 IN_N.n138 IN_N.n137 0.003
R22532 IN_N.n140 IN_N.n139 0.003
R22533 IN_N.n142 IN_N.n141 0.003
R22534 IN_N.n125 IN_N.n124 0.003
R22535 IN_N.n114 IN_N.n113 0.003
R22536 IN_N.n72 IN_N.n71 0.003
R22537 IN_N.n67 IN_N.n66 0.003
R22538 IN_N.n77 IN_N.n76 0.003
R22539 IN_N.n87 IN_N.n79 0.003
R22540 IN_N.n331 IN_N.n323 0.003
R22541 IN_N.n378 IN_N.n370 0.003
R22542 IN_N.n370 IN_N.n368 0.003
R22543 IN_N.n8 IN_N.n7 0.003
R22544 IN_N.n353 IN_N.n352 0.003
R22545 IN_N.n226 IN_N.n225 0.002
R22546 IN_N.n167 IN_N.n166 0.002
R22547 IN_N.n128 IN_N.n127 0.002
R22548 IN_N.n69 IN_N.n68 0.002
R22549 IN_N.n304 IN_N.n303 0.002
R22550 IN_N.n302 IN_N.n301 0.002
R22551 IN_N.n246 IN_N.n245 0.002
R22552 IN_N.n220 IN_N.n219 0.001
R22553 IN_N.n189 IN_N.n188 0.001
R22554 IN_N.n271 IN_N.n268 0.001
R22555 IN_N.n268 IN_N.n267 0.001
R22556 IN_N.n28 IN_N.n27 0.001
R22557 IN_N.n27 IN_N.n26 0.001
R22558 IN_N.n137 IN_N.n136 0.001
R22559 IN_N.n141 IN_N.n140 0.001
R22560 IN_N.n145 IN_N.n144 0.001
R22561 IN_N.n122 IN_N.n121 0.001
R22562 IN_N.n91 IN_N.n90 0.001
R22563 IN_N.n338 IN_N.n337 0.001
R22564 IN_N.n339 IN_N.n338 0.001
R22565 IN_N.n345 IN_N.n344 0.001
R22566 IN_N.n346 IN_N.n345 0.001
R22567 OUT_N.n33 OUT_N.n32 9.305
R22568 OUT_N.n252 OUT_N.n251 9.305
R22569 OUT_N.n96 OUT_N.n95 9.3
R22570 OUT_N.n16 OUT_N.n15 9.3
R22571 OUT_N.n94 OUT_N.n93 9.3
R22572 OUT_N.n136 OUT_N.n135 9.3
R22573 OUT_N.n127 OUT_N.n126 9.3
R22574 OUT_N.n130 OUT_N.n129 9.3
R22575 OUT_N.n132 OUT_N.n131 9.3
R22576 OUT_N.n114 OUT_N.n113 9.3
R22577 OUT_N.n110 OUT_N.n109 9.3
R22578 OUT_N.n107 OUT_N.n106 9.3
R22579 OUT_N.n103 OUT_N.n102 9.3
R22580 OUT_N.n118 OUT_N.n117 9.3
R22581 OUT_N.n121 OUT_N.n120 9.3
R22582 OUT_N.n123 OUT_N.n122 9.3
R22583 OUT_N.n26 OUT_N.n25 9.3
R22584 OUT_N.n24 OUT_N.n23 9.3
R22585 OUT_N.n38 OUT_N.n37 9.3
R22586 OUT_N.n63 OUT_N.n62 9.3
R22587 OUT_N.n61 OUT_N.n60 9.3
R22588 OUT_N.n58 OUT_N.n57 9.3
R22589 OUT_N.n41 OUT_N.n40 9.3
R22590 OUT_N.n45 OUT_N.n44 9.3
R22591 OUT_N.n49 OUT_N.n48 9.3
R22592 OUT_N.n52 OUT_N.n51 9.3
R22593 OUT_N.n54 OUT_N.n53 9.3
R22594 OUT_N.n82 OUT_N.n81 9.3
R22595 OUT_N.n67 OUT_N.n66 9.3
R22596 OUT_N.n216 OUT_N.n215 9.3
R22597 OUT_N.n210 OUT_N.n209 9.3
R22598 OUT_N.n214 OUT_N.n213 9.3
R22599 OUT_N.n220 OUT_N.n219 9.3
R22600 OUT_N.n235 OUT_N.n234 9.3
R22601 OUT_N.n178 OUT_N.n177 9.3
R22602 OUT_N.n180 OUT_N.n179 9.3
R22603 OUT_N.n206 OUT_N.n205 9.3
R22604 OUT_N.n204 OUT_N.n203 9.3
R22605 OUT_N.n200 OUT_N.n199 9.3
R22606 OUT_N.n196 OUT_N.n195 9.3
R22607 OUT_N.n191 OUT_N.n190 9.3
R22608 OUT_N.n188 OUT_N.n187 9.3
R22609 OUT_N.n183 OUT_N.n182 9.3
R22610 OUT_N.n257 OUT_N.n256 9.3
R22611 OUT_N.n265 OUT_N.n264 9.3
R22612 OUT_N.n275 OUT_N.n274 9.3
R22613 OUT_N.n285 OUT_N.n284 9.3
R22614 OUT_N.n295 OUT_N.n294 9.3
R22615 OUT_N.n269 OUT_N.n268 9.3
R22616 OUT_N.n273 OUT_N.n272 9.3
R22617 OUT_N.n279 OUT_N.n278 9.3
R22618 OUT_N.n283 OUT_N.n282 9.3
R22619 OUT_N.n289 OUT_N.n288 9.3
R22620 OUT_N.n293 OUT_N.n292 9.3
R22621 OUT_N.n168 OUT_N.n167 9.3
R22622 OUT_N.n260 OUT_N.n259 9.3
R22623 OUT_N.n104 OUT_N.n101 9
R22624 OUT_N.n112 OUT_N.n100 9
R22625 OUT_N.n43 OUT_N.n31 9
R22626 OUT_N.n50 OUT_N.n30 9
R22627 OUT_N.n119 OUT_N.n99 9
R22628 OUT_N.n17 OUT_N.n13 9
R22629 OUT_N.n86 OUT_N.n85 9
R22630 OUT_N.n6 OUT_N.n5 9
R22631 OUT_N.n138 OUT_N.n137 9
R22632 OUT_N.n59 OUT_N.n29 9
R22633 OUT_N.n128 OUT_N.n98 9
R22634 OUT_N.n83 OUT_N.n75 9
R22635 OUT_N.n35 OUT_N.n34 9
R22636 OUT_N.n68 OUT_N.n28 9
R22637 OUT_N.n185 OUT_N.n184 9
R22638 OUT_N.n194 OUT_N.n193 9
R22639 OUT_N.n202 OUT_N.n201 9
R22640 OUT_N.n170 OUT_N.n169 9
R22641 OUT_N.n271 OUT_N.n270 9
R22642 OUT_N.n281 OUT_N.n280 9
R22643 OUT_N.n291 OUT_N.n290 9
R22644 OUT_N.n231 OUT_N.n230 9
R22645 OUT_N.n237 OUT_N.n236 9
R22646 OUT_N.n212 OUT_N.n211 9
R22647 OUT_N.n222 OUT_N.n221 9
R22648 OUT_N.n299 OUT_N.n298 9
R22649 OUT_N.n263 OUT_N.n262 9
R22650 OUT_N.n254 OUT_N.n253 9
R22651 OUT_N.n9 OUT_N.n8 8.097
R22652 OUT_N.n71 OUT_N.n70 8.097
R22653 OUT_N.n239 OUT_N.n238 8.097
R22654 OUT_N.n172 OUT_N.n171 8.097
R22655 OUT_N.n3 OUT_N.n2 4.574
R22656 OUT_N.n79 OUT_N.n78 4.574
R22657 OUT_N.n227 OUT_N.n226 4.574
R22658 OUT_N.n165 OUT_N.n164 4.574
R22659 OUT_N.n2 OUT_N.n0 3.388
R22660 OUT_N.n78 OUT_N.n76 3.388
R22661 OUT_N.n226 OUT_N.n225 3.388
R22662 OUT_N.n164 OUT_N.n163 3.388
R22663 OUT_N.n9 OUT_N.t7 3.326
R22664 OUT_N.n9 OUT_N.t1 3.326
R22665 OUT_N.n71 OUT_N.t4 3.326
R22666 OUT_N.n71 OUT_N.t5 3.326
R22667 OUT_N.n239 OUT_N.t3 3.326
R22668 OUT_N.n239 OUT_N.t0 3.326
R22669 OUT_N.n172 OUT_N.t2 3.326
R22670 OUT_N.n172 OUT_N.t6 3.326
R22671 OUT_N.n90 OUT_N.n69 2.473
R22672 OUT_N.n140 OUT_N.n139 2.473
R22673 OUT_N.n248 OUT_N.n223 2.473
R22674 OUT_N.n247 OUT_N.n242 2.473
R22675 OUT_N.n303 OUT_N.n297 2.473
R22676 OUT_N.n141 OUT_N.n7 2.473
R22677 OUT_N.n248 OUT_N.n232 2.467
R22678 OUT_N.n303 OUT_N.n302 2.467
R22679 OUT_N.n90 OUT_N.n89 2.467
R22680 OUT_N.n140 OUT_N.n18 2.466
R22681 OUT_N.n90 OUT_N.n84 2.466
R22682 OUT_N.n303 OUT_N.n176 2.466
R22683 OUT_N.n155 OUT_N.n154 1.418
R22684 OUT_N.n10 OUT_N.n9 1.155
R22685 OUT_N.n72 OUT_N.n71 1.155
R22686 OUT_N.n173 OUT_N.n172 1.155
R22687 OUT_N.n240 OUT_N.n239 1.155
R22688 OUT_N.n11 OUT_N.n10 0.873
R22689 OUT_N.n73 OUT_N.n72 0.873
R22690 OUT_N.n174 OUT_N.n173 0.873
R22691 OUT_N.n241 OUT_N.n240 0.873
R22692 OUT_N.n2 OUT_N.n1 0.506
R22693 OUT_N.n78 OUT_N.n77 0.506
R22694 OUT_N.n226 OUT_N.n224 0.506
R22695 OUT_N.n164 OUT_N.n162 0.506
R22696 OUT_N.n135 OUT_N.n134 0.476
R22697 OUT_N.n66 OUT_N.n65 0.476
R22698 OUT_N.n219 OUT_N.n218 0.476
R22699 OUT_N.n288 OUT_N.n287 0.476
R22700 OUT_N.n154 OUT_N 0.466
R22701 OUT_N.n126 OUT_N.n125 0.445
R22702 OUT_N.n57 OUT_N.n56 0.445
R22703 OUT_N.n209 OUT_N.n208 0.445
R22704 OUT_N.n278 OUT_N.n277 0.445
R22705 OUT_N.n117 OUT_N.n116 0.414
R22706 OUT_N.n48 OUT_N.n47 0.414
R22707 OUT_N.n199 OUT_N.n198 0.414
R22708 OUT_N.n268 OUT_N.n267 0.414
R22709 OUT_N.n154 OUT_N.n153 0.392
R22710 OUT_N.n153 OUT_N.n145 0.231
R22711 OUT_N.n147 OUT_N.n146 0.23
R22712 OUT_N.n308 OUT_N.n161 0.23
R22713 OUT_N.n124 OUT_N.n123 0.073
R22714 OUT_N.n55 OUT_N.n54 0.073
R22715 OUT_N.n207 OUT_N.n206 0.073
R22716 OUT_N.n276 OUT_N.n275 0.073
R22717 OUT_N.n110 OUT_N.n108 0.073
R22718 OUT_N.n41 OUT_N.n39 0.073
R22719 OUT_N.n191 OUT_N.n189 0.073
R22720 OUT_N.n260 OUT_N.n258 0.073
R22721 OUT_N.n115 OUT_N.n114 0.072
R22722 OUT_N.n46 OUT_N.n45 0.072
R22723 OUT_N.n197 OUT_N.n196 0.072
R22724 OUT_N.n266 OUT_N.n265 0.072
R22725 OUT_N.n133 OUT_N.n132 0.062
R22726 OUT_N.n64 OUT_N.n63 0.062
R22727 OUT_N.n217 OUT_N.n216 0.062
R22728 OUT_N.n286 OUT_N.n285 0.062
R22729 OUT_N.n49 OUT_N.n46 0.057
R22730 OUT_N.n269 OUT_N.n266 0.057
R22731 OUT_N.n200 OUT_N.n197 0.057
R22732 OUT_N.n118 OUT_N.n115 0.057
R22733 OUT_N.n88 OUT_N.n87 0.055
R22734 OUT_N.n229 OUT_N.n228 0.055
R22735 OUT_N.n301 OUT_N.n300 0.055
R22736 OUT_N.n7 OUT_N.n4 0.055
R22737 OUT_N.n136 OUT_N.n133 0.054
R22738 OUT_N.n67 OUT_N.n64 0.054
R22739 OUT_N.n220 OUT_N.n217 0.054
R22740 OUT_N.n289 OUT_N.n286 0.054
R22741 OUT_N.n108 OUT_N.n107 0.054
R22742 OUT_N.n39 OUT_N.n38 0.054
R22743 OUT_N.n189 OUT_N.n188 0.054
R22744 OUT_N.n258 OUT_N.n257 0.054
R22745 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN OUT_N.n308 0.042
R22746 OUT_N.n12 OUT_N.n11 0.041
R22747 OUT_N.n74 OUT_N.n73 0.041
R22748 OUT_N.n242 OUT_N.n241 0.041
R22749 OUT_N.n175 OUT_N.n174 0.041
R22750 OUT_N.n242 OUT_N.n237 0.04
R22751 OUT_N.n146 OUT_N 0.04
R22752 OUT_N.n127 OUT_N.n124 0.039
R22753 OUT_N.n58 OUT_N.n55 0.039
R22754 OUT_N.n210 OUT_N.n207 0.039
R22755 OUT_N.n279 OUT_N.n276 0.039
R22756 OUT_N.n7 OUT_N.n6 0.031
R22757 OUT_N.n130 OUT_N.n128 0.031
R22758 OUT_N.n61 OUT_N.n59 0.031
R22759 OUT_N.n214 OUT_N.n212 0.031
R22760 OUT_N.n283 OUT_N.n281 0.031
R22761 OUT_N.n18 OUT_N.n17 0.029
R22762 OUT_N.n84 OUT_N.n83 0.029
R22763 OUT_N.n176 OUT_N.n170 0.029
R22764 OUT_N.n107 OUT_N.n105 0.028
R22765 OUT_N.n188 OUT_N.n186 0.028
R22766 OUT_N.n97 OUT_N.n96 0.026
R22767 OUT_N.n121 OUT_N.n119 0.026
R22768 OUT_N.n114 OUT_N.n112 0.026
R22769 OUT_N.n27 OUT_N.n26 0.026
R22770 OUT_N.n52 OUT_N.n50 0.026
R22771 OUT_N.n45 OUT_N.n43 0.026
R22772 OUT_N.n196 OUT_N.n194 0.026
R22773 OUT_N.n204 OUT_N.n202 0.026
R22774 OUT_N.n181 OUT_N.n180 0.026
R22775 OUT_N.n265 OUT_N.n263 0.026
R22776 OUT_N.n273 OUT_N.n271 0.026
R22777 OUT_N.n296 OUT_N.n295 0.026
R22778 OUT_N.n38 OUT_N.n36 0.024
R22779 OUT_N.n257 OUT_N.n255 0.024
R22780 OUT_N.n92 OUT_N.n91 0.024
R22781 OUT_N.n4 OUT_N.n3 0.023
R22782 OUT_N.n89 OUT_N.n86 0.023
R22783 OUT_N.n232 OUT_N.n231 0.023
R22784 OUT_N.n302 OUT_N.n299 0.023
R22785 OUT_N.n228 OUT_N.n227 0.023
R22786 OUT_N.n250 OUT_N.n249 0.022
R22787 OUT_N.n80 OUT_N.n79 0.021
R22788 OUT_N.n166 OUT_N.n165 0.021
R22789 OUT_N.n308 OUT_N.n307 0.02
R22790 OUT_N.n153 OUT_N.n152 0.019
R22791 OUT_N.n156 OUT_N.n155 0.019
R22792 OUT_N.n16 OUT_N.n14 0.019
R22793 OUT_N.n82 OUT_N.n80 0.019
R22794 OUT_N.n235 OUT_N.n233 0.019
R22795 OUT_N.n168 OUT_N.n166 0.019
R22796 OUT_N.n159 OUT_N.n158 0.016
R22797 OUT_N.n150 OUT_N.n149 0.016
R22798 OUT_N.n17 OUT_N.n16 0.014
R22799 OUT_N.n123 OUT_N.n121 0.014
R22800 OUT_N.n119 OUT_N.n118 0.014
R22801 OUT_N.n83 OUT_N.n82 0.014
R22802 OUT_N.n54 OUT_N.n52 0.014
R22803 OUT_N.n50 OUT_N.n49 0.014
R22804 OUT_N.n202 OUT_N.n200 0.014
R22805 OUT_N.n206 OUT_N.n204 0.014
R22806 OUT_N.n237 OUT_N.n235 0.014
R22807 OUT_N.n271 OUT_N.n269 0.014
R22808 OUT_N.n275 OUT_N.n273 0.014
R22809 OUT_N.n170 OUT_N.n168 0.014
R22810 OUT_N.n176 OUT_N.n175 0.011
R22811 OUT_N.n84 OUT_N.n74 0.011
R22812 OUT_N.n18 OUT_N.n12 0.011
R22813 OUT_N.n132 OUT_N.n130 0.009
R22814 OUT_N.n128 OUT_N.n127 0.009
R22815 OUT_N.n104 OUT_N.n103 0.009
R22816 OUT_N.n63 OUT_N.n61 0.009
R22817 OUT_N.n59 OUT_N.n58 0.009
R22818 OUT_N.n185 OUT_N.n183 0.009
R22819 OUT_N.n212 OUT_N.n210 0.009
R22820 OUT_N.n216 OUT_N.n214 0.009
R22821 OUT_N.n281 OUT_N.n279 0.009
R22822 OUT_N.n285 OUT_N.n283 0.009
R22823 OUT_N.n89 OUT_N.n88 0.009
R22824 OUT_N.n302 OUT_N.n301 0.009
R22825 OUT_N.n232 OUT_N.n229 0.009
R22826 OUT_N.n111 OUT_N.n110 0.008
R22827 OUT_N.n42 OUT_N.n41 0.008
R22828 OUT_N.n192 OUT_N.n191 0.008
R22829 OUT_N.n261 OUT_N.n260 0.008
R22830 OUT_N.n157 OUT_N.n156 0.008
R22831 OUT_N.n161 OUT_N.n160 0.008
R22832 OUT_N.n152 OUT_N.n151 0.008
R22833 OUT_N.n148 OUT_N.n147 0.008
R22834 OUT_N.n140 OUT_N.n92 0.008
R22835 OUT_N.n249 OUT_N.n248 0.008
R22836 OUT_N.n91 OUT_N.n90 0.007
R22837 OUT_N.n303 OUT_N.n250 0.007
R22838 OUT_N.n36 OUT_N.n35 0.007
R22839 OUT_N.n255 OUT_N.n254 0.007
R22840 OUT_N.n112 OUT_N.n111 0.006
R22841 OUT_N.n43 OUT_N.n42 0.006
R22842 OUT_N.n194 OUT_N.n192 0.006
R22843 OUT_N.n263 OUT_N.n261 0.006
R22844 OUT_N.n158 OUT_N.n157 0.005
R22845 OUT_N.n160 OUT_N.n159 0.005
R22846 OUT_N.n151 OUT_N.n150 0.005
R22847 OUT_N.n149 OUT_N.n148 0.005
R22848 OUT_N.n35 OUT_N.n33 0.005
R22849 OUT_N.n254 OUT_N.n252 0.005
R22850 OUT_N.n96 OUT_N.n94 0.004
R22851 OUT_N.n138 OUT_N.n136 0.004
R22852 OUT_N.n26 OUT_N.n24 0.004
R22853 OUT_N.n68 OUT_N.n67 0.004
R22854 OUT_N.n144 OUT_N.n143 0.004
R22855 OUT_N.n21 OUT_N.n20 0.004
R22856 OUT_N.n222 OUT_N.n220 0.004
R22857 OUT_N.n180 OUT_N.n178 0.004
R22858 OUT_N.n291 OUT_N.n289 0.004
R22859 OUT_N.n295 OUT_N.n293 0.004
R22860 OUT_N.n245 OUT_N.n244 0.004
R22861 OUT_N.n306 OUT_N.n305 0.004
R22862 OUT_N.n105 OUT_N.n104 0.004
R22863 OUT_N.n186 OUT_N.n185 0.004
R22864 OUT_N.n139 OUT_N.n138 0.003
R22865 OUT_N.n69 OUT_N.n68 0.003
R22866 OUT_N.n142 OUT_N.n141 0.003
R22867 OUT_N.n223 OUT_N.n222 0.003
R22868 OUT_N.n247 OUT_N.n246 0.003
R22869 OUT_N.n297 OUT_N.n291 0.003
R22870 OUT_N.n90 OUT_N.n22 0.003
R22871 OUT_N.n304 OUT_N.n303 0.003
R22872 OUT_N.n141 OUT_N.n140 0.002
R22873 OUT_N.n297 OUT_N.n296 0.002
R22874 OUT_N.n223 OUT_N.n181 0.002
R22875 OUT_N.n248 OUT_N.n247 0.002
R22876 OUT_N.n139 OUT_N.n97 0.002
R22877 OUT_N.n69 OUT_N.n27 0.002
R22878 OUT_N.n145 OUT_N.n144 0.001
R22879 OUT_N.n143 OUT_N.n142 0.001
R22880 OUT_N.n22 OUT_N.n21 0.001
R22881 OUT_N.n20 OUT_N.n19 0.001
R22882 OUT_N.n244 OUT_N.n243 0.001
R22883 OUT_N.n246 OUT_N.n245 0.001
R22884 OUT_N.n305 OUT_N.n304 0.001
R22885 OUT_N.n307 OUT_N.n306 0.001
R22886 IN_P.n61 IN_P.t3 846.712
R22887 IN_P.n30 IN_P.t6 846.712
R22888 IN_P.n7 IN_P.t0 846.712
R22889 IN_P.n45 IN_P.t4 846.712
R22890 IN_P.n323 IN_P.t5 846.712
R22891 IN_P.n353 IN_P.t1 846.712
R22892 IN_P.n338 IN_P.t2 846.712
R22893 IN_P.n2 IN_P.t7 846.712
R22894 IN_P.n46 IN_P.n45 15.887
R22895 IN_P.n9 IN_P.n7 15.887
R22896 IN_P.n90 IN_P.n89 15.887
R22897 IN_P.n187 IN_P.n186 15.887
R22898 IN_P.n3 IN_P.n2 15.887
R22899 IN_P.n339 IN_P.n338 15.887
R22900 IN_P.n100 IN_P.n99 12.054
R22901 IN_P.n197 IN_P.n196 12.054
R22902 IN_P.n63 IN_P.n62 10.328
R22903 IN_P.n32 IN_P.n31 10.328
R22904 IN_P.n122 IN_P.n121 10.328
R22905 IN_P.n145 IN_P.n144 10.328
R22906 IN_P.n219 IN_P.n218 10.328
R22907 IN_P.n242 IN_P.n241 10.328
R22908 IN_P.n325 IN_P.n324 10.328
R22909 IN_P.n355 IN_P.n354 10.328
R22910 IN_P.n55 IN_P.n54 9.3
R22911 IN_P.n24 IN_P.n5 9.3
R22912 IN_P.n66 IN_P.n65 9.3
R22913 IN_P.n65 IN_P.n64 9.3
R22914 IN_P.n35 IN_P.n34 9.3
R22915 IN_P.n34 IN_P.n33 9.3
R22916 IN_P.n147 IN_P.n146 9.3
R22917 IN_P.n114 IN_P.n113 9.3
R22918 IN_P.n125 IN_P.n124 9.3
R22919 IN_P.n124 IN_P.n123 9.3
R22920 IN_P.n211 IN_P.n210 9.3
R22921 IN_P.n244 IN_P.n243 9.3
R22922 IN_P.n222 IN_P.n221 9.3
R22923 IN_P.n221 IN_P.n220 9.3
R22924 IN_P.n347 IN_P.n346 9.3
R22925 IN_P.n358 IN_P.n357 9.3
R22926 IN_P.n357 IN_P.n356 9.3
R22927 IN_P.n328 IN_P.n327 9.3
R22928 IN_P.n327 IN_P.n326 9.3
R22929 IN_P.n318 IN_P.n317 9.3
R22930 IN_P.n117 IN_P.n116 9
R22931 IN_P.n214 IN_P.n213 9
R22932 IN_P.n350 IN_P.n349 9
R22933 IN_P.n320 IN_P.n319 9
R22934 IN_P.n27 IN_P.n26 9
R22935 IN_P.n58 IN_P.n57 9
R22936 IN_P.n72 IN_P.n71 8.764
R22937 IN_P.n132 IN_P.n131 8.764
R22938 IN_P.n229 IN_P.n228 8.764
R22939 IN_P.n332 IN_P.n331 8.764
R22940 IN_P.n48 IN_P.n47 7.008
R22941 IN_P.n341 IN_P.n340 7.008
R22942 IN_P.n62 IN_P.n61 6.885
R22943 IN_P.n31 IN_P.n30 6.885
R22944 IN_P.n121 IN_P.n120 6.885
R22945 IN_P.n144 IN_P.n143 6.885
R22946 IN_P.n218 IN_P.n217 6.885
R22947 IN_P.n241 IN_P.n240 6.885
R22948 IN_P.n324 IN_P.n323 6.885
R22949 IN_P.n354 IN_P.n353 6.885
R22950 IN_P.n46 IN_P.n43 6.276
R22951 IN_P.n9 IN_P.n8 6.276
R22952 IN_P.n90 IN_P.n87 6.276
R22953 IN_P.n187 IN_P.n184 6.276
R22954 IN_P.n3 IN_P.n0 6.276
R22955 IN_P.n339 IN_P.n336 6.276
R22956 IN_P.n60 IN_P.n59 5.647
R22957 IN_P.n29 IN_P.n28 5.647
R22958 IN_P.n119 IN_P.n118 5.647
R22959 IN_P.n142 IN_P.n141 5.647
R22960 IN_P.n216 IN_P.n215 5.647
R22961 IN_P.n239 IN_P.n238 5.647
R22962 IN_P.n322 IN_P.n321 5.647
R22963 IN_P.n352 IN_P.n351 5.647
R22964 IN_P.n101 IN_P.n100 4.934
R22965 IN_P.n198 IN_P.n197 4.934
R22966 IN_P.n95 IN_P.n94 4.894
R22967 IN_P.n192 IN_P.n191 4.894
R22968 IN_P.n99 IN_P.n98 4.82
R22969 IN_P.n196 IN_P.n195 4.82
R22970 IN_P.n139 IN_P.n138 4.65
R22971 IN_P.n236 IN_P.n235 4.65
R22972 IN_P.n148 IN_P.n147 4.574
R22973 IN_P.n133 IN_P.n132 4.574
R22974 IN_P.n245 IN_P.n244 4.574
R22975 IN_P.n230 IN_P.n229 4.574
R22976 IN_P.n333 IN_P.n332 4.574
R22977 IN_P.n73 IN_P.n72 4.574
R22978 IN_P.n45 IN_P.n44 4.131
R22979 IN_P.n7 IN_P.n6 4.131
R22980 IN_P.n89 IN_P.n88 4.131
R22981 IN_P.n98 IN_P.n97 4.131
R22982 IN_P.n186 IN_P.n185 4.131
R22983 IN_P.n195 IN_P.n194 4.131
R22984 IN_P.n2 IN_P.n1 4.131
R22985 IN_P.n338 IN_P.n337 4.131
R22986 IN_P.n316 IN_P.n3 4.129
R22987 IN_P.n21 IN_P.n9 4.11
R22988 IN_P.n91 IN_P.n90 3.739
R22989 IN_P.n188 IN_P.n187 3.737
R22990 IN_P.n104 IN_P.n103 3
R22991 IN_P.n150 IN_P.n149 3
R22992 IN_P.n201 IN_P.n200 3
R22993 IN_P.n247 IN_P.n246 3
R22994 IN_P.n281 IN_P.n280 2.606
R22995 IN_P.n75 IN_P.n74 2.473
R22996 IN_P.n39 IN_P.n38 2.473
R22997 IN_P.n282 IN_P.n183 1.905
R22998 IN_P.n283 IN_P.n282 1.705
R22999 IN_P.n64 IN_P.n63 1.377
R23000 IN_P.n33 IN_P.n32 1.377
R23001 IN_P.n123 IN_P.n122 1.377
R23002 IN_P.n146 IN_P.n145 1.377
R23003 IN_P.n220 IN_P.n219 1.377
R23004 IN_P.n243 IN_P.n242 1.377
R23005 IN_P.n326 IN_P.n325 1.377
R23006 IN_P.n356 IN_P.n355 1.377
R23007 IN_P.n316 IN_P.n315 1.37
R23008 IN_P.n21 IN_P.n20 1.185
R23009 IN_P.n171 IN_P.n91 1.182
R23010 IN_P.n268 IN_P.n188 1.181
R23011 IN_P.n296 IN_P.n295 1.152
R23012 IN_P.n172 IN_P.n171 1.151
R23013 IN_P.n269 IN_P.n268 1.141
R23014 IN_P.n301 IN_P.n300 0.859
R23015 IN_P.n65 IN_P.n60 0.752
R23016 IN_P.n34 IN_P.n29 0.752
R23017 IN_P.n124 IN_P.n119 0.752
R23018 IN_P.n147 IN_P.n142 0.752
R23019 IN_P.n96 IN_P.n95 0.752
R23020 IN_P.n100 IN_P.n96 0.752
R23021 IN_P.n221 IN_P.n216 0.752
R23022 IN_P.n244 IN_P.n239 0.752
R23023 IN_P.n193 IN_P.n192 0.752
R23024 IN_P.n197 IN_P.n193 0.752
R23025 IN_P.n327 IN_P.n322 0.752
R23026 IN_P.n357 IN_P.n352 0.752
R23027 IN_P.n284 IN_P.n283 0.369
R23028 IN_P.n86 IN_P 0.2
R23029 IN_P.n47 IN_P.n46 0.11
R23030 IN_P.n340 IN_P.n339 0.11
R23031 IN_P.n318 IN_P.n316 0.083
R23032 IN_P.n53 IN_P.n52 0.054
R23033 IN_P.n74 IN_P.n68 0.054
R23034 IN_P.n330 IN_P.n329 0.054
R23035 IN_P.n313 IN_P.n312 0.054
R23036 IN_P.n309 IN_P.n308 0.054
R23037 IN_P.n23 IN_P.n22 0.051
R23038 IN_P.n282 IN_P.n281 0.049
R23039 IN_P.n345 IN_P.n344 0.049
R23040 IN_P.n305 IN_P.n304 0.049
R23041 IN_P.n283 IN_P.n86 0.049
R23042 IN_P.n209 IN_P.n208 0.047
R23043 IN_P.n112 IN_P.n111 0.047
R23044 IN_P.n225 IN_P.n224 0.045
R23045 IN_P.n128 IN_P.n127 0.045
R23046 IN_P.n329 IN_P.n328 0.039
R23047 IN_P.n335 IN_P.n334 0.039
R23048 IN_P.n314 IN_P.n313 0.039
R23049 IN_P.n310 IN_P.n309 0.039
R23050 IN_P.n306 IN_P.n305 0.039
R23051 IN_P.n22 IN_P.n21 0.038
R23052 IN_P.n40 IN_P.n39 0.038
R23053 IN_P.n300 IN_P.n299 0.038
R23054 IN_P IN_P.n232 0.037
R23055 IN_P.n74 IN_P.n73 0.037
R23056 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE IN_P.n135 0.037
R23057 IN_P.n333 IN_P.n330 0.037
R23058 IN_P.n312 IN_P.n311 0.037
R23059 IN_P.n308 IN_P.n307 0.037
R23060 IN_P.n302 IN_P.n301 0.037
R23061 IN_P.n295 IN_P.n294 0.037
R23062 IN_P.n84 IN_P.n83 0.036
R23063 IN_P.n75 IN_P.n42 0.036
R23064 IN_P.n111 IN_P.n91 0.035
R23065 IN_P.n52 IN_P.n51 0.035
R23066 IN_P.n344 IN_P.n343 0.035
R23067 IN_P.n304 IN_P.n303 0.035
R23068 IN_P.n287 IN_P.n286 0.035
R23069 IN_P.n208 IN_P.n188 0.035
R23070 IN_P.n227 IN_P.n226 0.034
R23071 IN_P.n130 IN_P.n129 0.034
R23072 IN_P.n359 IN_P.n358 0.034
R23073 IN_P.n38 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE 0.032
R23074 IN_P IN_P.n335 0.032
R23075 IN_P.n17 IN_P.n16 0.031
R23076 IN_P.n296 IN_P.n85 0.03
R23077 IN_P.n200 IN_P.n199 0.03
R23078 IN_P.n103 IN_P.n102 0.03
R23079 IN_P.n173 IN_P.n172 0.029
R23080 IN_P.n181 IN_P.n180 0.029
R23081 IN_P.n291 IN_P.n290 0.029
R23082 IN_P.n320 IN_P.n318 0.028
R23083 IN_P.n108 IN_P.n107 0.027
R23084 IN_P.n205 IN_P.n204 0.027
R23085 IN_P.n39 IN_P.n4 0.027
R23086 IN_P.n237 IN_P.n236 0.026
R23087 IN_P.n140 IN_P.n139 0.026
R23088 IN_P.n177 IN_P.n176 0.025
R23089 IN_P.n76 IN_P.n75 0.025
R23090 IN_P.n19 IN_P.n18 0.025
R23091 IN_P.n214 IN_P.n212 0.024
R23092 IN_P.n231 IN_P.n230 0.024
R23093 IN_P.n25 IN_P.n24 0.024
R23094 IN_P.n117 IN_P.n115 0.024
R23095 IN_P.n134 IN_P.n133 0.024
R23096 IN_P.n348 IN_P.n347 0.024
R23097 IN_P.n159 IN_P.n158 0.023
R23098 IN_P.n109 IN_P.n108 0.023
R23099 IN_P.n256 IN_P.n255 0.023
R23100 IN_P.n206 IN_P.n205 0.023
R23101 IN_P.n15 IN_P.n14 0.023
R23102 IN_P.n246 IN_P.n245 0.022
R23103 IN_P.n58 IN_P.n56 0.022
R23104 IN_P.n67 IN_P.n66 0.022
R23105 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE IN_P.n37 0.022
R23106 IN_P.n149 IN_P.n148 0.022
R23107 IN_P IN_P.n359 0.022
R23108 IN_P.n82 IN_P.n81 0.022
R23109 IN_P.n80 IN_P.n79 0.022
R23110 IN_P.n223 IN_P.n222 0.02
R23111 IN_P.n246 IN_P.n234 0.02
R23112 IN_P.n126 IN_P.n125 0.02
R23113 IN_P.n149 IN_P.n137 0.02
R23114 IN_P.n13 IN_P.n12 0.02
R23115 IN_P.n224 IN_P.n223 0.018
R23116 IN_P.n127 IN_P.n126 0.018
R23117 IN_P.n170 IN_P.n169 0.018
R23118 IN_P.n267 IN_P.n266 0.018
R23119 IN_P.n77 IN_P.n76 0.018
R23120 IN_P.n18 IN_P.n17 0.018
R23121 IN_P.n68 IN_P.n67 0.017
R23122 IN_P.n37 IN_P.n36 0.017
R23123 IN_P.n36 IN_P.n35 0.017
R23124 IN_P.n167 IN_P.n166 0.016
R23125 IN_P.n161 IN_P.n160 0.016
R23126 IN_P.n157 IN_P.n156 0.016
R23127 IN_P.n264 IN_P.n263 0.016
R23128 IN_P.n258 IN_P.n257 0.016
R23129 IN_P.n254 IN_P.n253 0.016
R23130 IN_P.n85 IN_P.n84 0.016
R23131 IN_P.n79 IN_P.n78 0.016
R23132 IN_P.n12 IN_P.n11 0.016
R23133 IN_P.n286 IN_P.n285 0.016
R23134 IN_P.n24 IN_P.n23 0.015
R23135 IN_P.n150 IN_P.n110 0.015
R23136 IN_P.n182 IN_P.n181 0.015
R23137 IN_P.n247 IN_P.n207 0.015
R23138 IN_P.n347 IN_P.n345 0.015
R23139 IN_P.n169 IN_P.n168 0.014
R23140 IN_P.n165 IN_P.n164 0.014
R23141 IN_P.n151 IN_P.n150 0.014
R23142 IN_P.n266 IN_P.n265 0.014
R23143 IN_P.n262 IN_P.n261 0.014
R23144 IN_P.n248 IN_P.n247 0.014
R23145 IN_P.n83 IN_P.n82 0.014
R23146 IN_P.n10 IN_P.n4 0.014
R23147 IN_P.n16 IN_P.n15 0.014
R23148 IN_P.n171 IN_P.n170 0.014
R23149 IN_P.n268 IN_P.n267 0.013
R23150 IN_P.n190 IN_P.n189 0.013
R23151 IN_P.n93 IN_P.n92 0.013
R23152 IN_P.n164 IN_P.n163 0.013
R23153 IN_P.n153 IN_P.n152 0.013
R23154 IN_P.n261 IN_P.n260 0.013
R23155 IN_P.n250 IN_P.n249 0.013
R23156 IN_P.n230 IN_P.n227 0.011
R23157 IN_P.n232 IN_P.n231 0.011
R23158 IN_P.n133 IN_P.n130 0.011
R23159 IN_P.n135 IN_P.n134 0.011
R23160 IN_P.n11 IN_P.n10 0.011
R23161 IN_P.n162 IN_P.n161 0.01
R23162 IN_P.n154 IN_P.n153 0.01
R23163 IN_P.n270 IN_P.n269 0.01
R23164 IN_P.n278 IN_P.n277 0.01
R23165 IN_P.n259 IN_P.n258 0.01
R23166 IN_P.n251 IN_P.n250 0.01
R23167 IN_P.n290 IN_P.n289 0.01
R23168 IN_P.n288 IN_P.n287 0.01
R23169 IN_P.n342 IN_P.n341 0.01
R23170 IN_P.n49 IN_P.n48 0.01
R23171 IN_P.n211 IN_P.n209 0.009
R23172 IN_P.n233 IN_P 0.009
R23173 IN_P.n55 IN_P.n53 0.009
R23174 IN_P.n114 IN_P.n112 0.009
R23175 IN_P.n136 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE 0.009
R23176 IN_P.n168 IN_P.n167 0.009
R23177 IN_P.n155 IN_P.n154 0.009
R23178 IN_P.n265 IN_P.n264 0.009
R23179 IN_P.n252 IN_P.n251 0.009
R23180 IN_P.n78 IN_P.n77 0.009
R23181 IN_P.n294 IN_P.n293 0.009
R23182 IN_P.n292 IN_P.n291 0.009
R23183 IN_P.n174 IN_P.n173 0.008
R23184 IN_P.n176 IN_P.n175 0.008
R23185 IN_P.n178 IN_P.n177 0.008
R23186 IN_P.n180 IN_P.n179 0.008
R23187 IN_P.n274 IN_P.n273 0.008
R23188 IN_P.n158 IN_P.n157 0.007
R23189 IN_P.n156 IN_P.n155 0.007
R23190 IN_P.n255 IN_P.n254 0.007
R23191 IN_P.n253 IN_P.n252 0.007
R23192 IN_P.n343 IN_P.n342 0.007
R23193 IN_P.n303 IN_P.n302 0.007
R23194 IN_P.n20 IN_P.n19 0.007
R23195 IN_P.n106 IN_P.n105 0.006
R23196 IN_P.n203 IN_P.n202 0.006
R23197 IN_P.n293 IN_P.n292 0.006
R23198 IN_P.n297 IN_P.n296 0.006
R23199 IN_P.n234 IN_P.n233 0.005
R23200 IN_P.n245 IN_P.n237 0.005
R23201 IN_P.n200 IN_P.n190 0.005
R23202 IN_P.n56 IN_P.n55 0.005
R23203 IN_P.n137 IN_P.n136 0.005
R23204 IN_P.n148 IN_P.n140 0.005
R23205 IN_P.n103 IN_P.n93 0.005
R23206 IN_P.n175 IN_P.n174 0.005
R23207 IN_P.n179 IN_P.n178 0.005
R23208 IN_P.n279 IN_P.n278 0.005
R23209 IN_P.n289 IN_P.n288 0.005
R23210 IN_P.n199 IN_P.n198 0.004
R23211 IN_P.n102 IN_P.n101 0.004
R23212 IN_P.n212 IN_P.n211 0.003
R23213 IN_P.n222 IN_P.n214 0.003
R23214 IN_P.n50 IN_P.n49 0.003
R23215 IN_P.n51 IN_P.n50 0.003
R23216 IN_P.n66 IN_P.n58 0.003
R23217 IN_P.n35 IN_P.n27 0.003
R23218 IN_P.n27 IN_P.n25 0.003
R23219 IN_P.n115 IN_P.n114 0.003
R23220 IN_P.n125 IN_P.n117 0.003
R23221 IN_P.n163 IN_P.n162 0.003
R23222 IN_P.n152 IN_P.n151 0.003
R23223 IN_P.n110 IN_P.n109 0.003
R23224 IN_P.n105 IN_P.n104 0.003
R23225 IN_P.n183 IN_P.n182 0.003
R23226 IN_P.n271 IN_P.n270 0.003
R23227 IN_P.n273 IN_P.n272 0.003
R23228 IN_P.n275 IN_P.n274 0.003
R23229 IN_P.n277 IN_P.n276 0.003
R23230 IN_P.n260 IN_P.n259 0.003
R23231 IN_P.n249 IN_P.n248 0.003
R23232 IN_P.n207 IN_P.n206 0.003
R23233 IN_P.n202 IN_P.n201 0.003
R23234 IN_P.n328 IN_P.n320 0.003
R23235 IN_P.n334 IN_P.n333 0.003
R23236 IN_P.n358 IN_P.n350 0.003
R23237 IN_P.n350 IN_P.n348 0.003
R23238 IN_P.n315 IN_P.n314 0.003
R23239 IN_P.n311 IN_P.n310 0.003
R23240 IN_P.n307 IN_P.n306 0.003
R23241 IN_P.n299 IN_P.n298 0.003
R23242 IN_P.n298 IN_P.n297 0.003
R23243 IN_P.n81 IN_P.n80 0.003
R23244 IN_P.n14 IN_P.n13 0.003
R23245 IN_P.n166 IN_P.n165 0.002
R23246 IN_P.n107 IN_P.n106 0.002
R23247 IN_P.n263 IN_P.n262 0.002
R23248 IN_P.n204 IN_P.n203 0.002
R23249 IN_P.n285 IN_P.n284 0.002
R23250 IN_P.n226 IN_P.n225 0.001
R23251 IN_P.n73 IN_P.n70 0.001
R23252 IN_P.n70 IN_P.n69 0.001
R23253 IN_P.n129 IN_P.n128 0.001
R23254 IN_P.n160 IN_P.n159 0.001
R23255 IN_P.n272 IN_P.n271 0.001
R23256 IN_P.n276 IN_P.n275 0.001
R23257 IN_P.n280 IN_P.n279 0.001
R23258 IN_P.n257 IN_P.n256 0.001
R23259 IN_P.n42 IN_P.n41 0.001
R23260 IN_P.n41 IN_P.n40 0.001
R23261 OUT_P.n187 OUT_P.n186 9.304
R23262 OUT_P.n155 OUT_P.n154 9.304
R23263 OUT_P.n29 OUT_P.n28 9.304
R23264 OUT_P.n1 OUT_P.n0 9.304
R23265 OUT_P.n268 OUT_P.n267 9.3
R23266 OUT_P.n264 OUT_P.n263 9.3
R23267 OUT_P.n165 OUT_P.n164 9.3
R23268 OUT_P.n159 OUT_P.n158 9.3
R23269 OUT_P.n254 OUT_P.n253 9.3
R23270 OUT_P.n260 OUT_P.n259 9.3
R23271 OUT_P.n145 OUT_P.n144 9.3
R23272 OUT_P.n147 OUT_P.n146 9.3
R23273 OUT_P.n170 OUT_P.n169 9.3
R23274 OUT_P.n153 OUT_P.n152 9.3
R23275 OUT_P.n258 OUT_P.n257 9.3
R23276 OUT_P.n270 OUT_P.n269 9.3
R23277 OUT_P.n278 OUT_P.n277 9.3
R23278 OUT_P.n190 OUT_P.n189 9.3
R23279 OUT_P.n213 OUT_P.n212 9.3
R23280 OUT_P.n215 OUT_P.n214 9.3
R23281 OUT_P.n232 OUT_P.n231 9.3
R23282 OUT_P.n219 OUT_P.n218 9.3
R23283 OUT_P.n224 OUT_P.n223 9.3
R23284 OUT_P.n222 OUT_P.n221 9.3
R23285 OUT_P.n209 OUT_P.n208 9.3
R23286 OUT_P.n196 OUT_P.n195 9.3
R23287 OUT_P.n200 OUT_P.n199 9.3
R23288 OUT_P.n183 OUT_P.n182 9.3
R23289 OUT_P.n178 OUT_P.n177 9.3
R23290 OUT_P.n176 OUT_P.n175 9.3
R23291 OUT_P.n33 OUT_P.n32 9.3
R23292 OUT_P.n39 OUT_P.n38 9.3
R23293 OUT_P.n44 OUT_P.n43 9.3
R23294 OUT_P.n71 OUT_P.n70 9.3
R23295 OUT_P.n52 OUT_P.n51 9.3
R23296 OUT_P.n79 OUT_P.n78 9.3
R23297 OUT_P.n81 OUT_P.n80 9.3
R23298 OUT_P.n85 OUT_P.n84 9.3
R23299 OUT_P.n89 OUT_P.n88 9.3
R23300 OUT_P.n91 OUT_P.n90 9.3
R23301 OUT_P.n67 OUT_P.n66 9.3
R23302 OUT_P.n75 OUT_P.n74 9.3
R23303 OUT_P.n46 OUT_P.n45 9.3
R23304 OUT_P.n5 OUT_P.n4 9.3
R23305 OUT_P.n117 OUT_P.n116 9.3
R23306 OUT_P.n24 OUT_P.n23 9.3
R23307 OUT_P.n121 OUT_P.n120 9.3
R23308 OUT_P.n16 OUT_P.n15 9.3
R23309 OUT_P.n11 OUT_P.n10 9.3
R23310 OUT_P.n131 OUT_P.n130 9.3
R23311 OUT_P.n135 OUT_P.n134 9.3
R23312 OUT_P.n127 OUT_P.n126 9.3
R23313 OUT_P.n125 OUT_P.n124 9.3
R23314 OUT_P.n137 OUT_P.n136 9.3
R23315 OUT_P.n113 OUT_P.n112 9.3
R23316 OUT_P.n19 OUT_P.n18 9.3
R23317 OUT_P.n230 OUT_P.n229 9
R23318 OUT_P.n198 OUT_P.n184 9
R23319 OUT_P.n180 OUT_P.n174 9
R23320 OUT_P.n220 OUT_P.n205 9
R23321 OUT_P.n225 OUT_P.n204 9
R23322 OUT_P.n211 OUT_P.n210 9
R23323 OUT_P.n150 OUT_P.n149 9
R23324 OUT_P.n256 OUT_P.n255 9
R23325 OUT_P.n157 OUT_P.n156 9
R23326 OUT_P.n168 OUT_P.n167 9
R23327 OUT_P.n266 OUT_P.n265 9
R23328 OUT_P.n271 OUT_P.n250 9
R23329 OUT_P.n276 OUT_P.n275 9
R23330 OUT_P.n188 OUT_P.n185 9
R23331 OUT_P.n14 OUT_P.n13 9
R23332 OUT_P.n111 OUT_P.n107 9
R23333 OUT_P.n65 OUT_P.n61 9
R23334 OUT_P.n123 OUT_P.n122 9
R23335 OUT_P.n133 OUT_P.n132 9
R23336 OUT_P.n139 OUT_P.n138 9
R23337 OUT_P.n87 OUT_P.n86 9
R23338 OUT_P.n93 OUT_P.n92 9
R23339 OUT_P.n77 OUT_P.n76 9
R23340 OUT_P.n49 OUT_P.n48 9
R23341 OUT_P.n42 OUT_P.n41 9
R23342 OUT_P.n31 OUT_P.n30 9
R23343 OUT_P.n21 OUT_P.n17 9
R23344 OUT_P.n3 OUT_P.n2 9
R23345 OUT_P.n237 OUT_P.n236 4.574
R23346 OUT_P.n283 OUT_P.n282 4.574
R23347 OUT_P.n115 OUT_P.n106 4.574
R23348 OUT_P.n69 OUT_P.n60 4.574
R23349 OUT_P.n282 OUT_P.n280 3.388
R23350 OUT_P.n236 OUT_P.n234 3.388
R23351 OUT_P.n60 OUT_P.n59 3.388
R23352 OUT_P.n106 OUT_P.n105 3.388
R23353 OUT_P.n272 OUT_P.t0 3.326
R23354 OUT_P.n272 OUT_P.t2 3.326
R23355 OUT_P.n226 OUT_P.t6 3.326
R23356 OUT_P.n226 OUT_P.t5 3.326
R23357 OUT_P.n62 OUT_P.t3 3.326
R23358 OUT_P.n62 OUT_P.t4 3.326
R23359 OUT_P.n108 OUT_P.t1 3.326
R23360 OUT_P.n108 OUT_P.t7 3.326
R23361 OUT_P.n243 OUT_P.n203 2.473
R23362 OUT_P.n102 OUT_P.n27 2.473
R23363 OUT_P.n248 OUT_P.n173 2.473
R23364 OUT_P.n97 OUT_P.n55 2.473
R23365 OUT_P.n285 OUT_P.n284 2.231
R23366 OUT_P.n141 OUT_P.n140 2.231
R23367 OUT_P.n95 OUT_P.n94 2.231
R23368 OUT_P.n241 OUT_P.n238 2.231
R23369 OUT_P.n296 OUT_P.n295 1.608
R23370 OUT_P.n273 OUT_P.n272 1.155
R23371 OUT_P.n227 OUT_P.n226 1.155
R23372 OUT_P.n63 OUT_P.n62 1.155
R23373 OUT_P.n109 OUT_P.n108 1.155
R23374 OUT_P.n274 OUT_P.n273 0.921
R23375 OUT_P.n228 OUT_P.n227 0.921
R23376 OUT_P.n64 OUT_P.n63 0.921
R23377 OUT_P.n110 OUT_P.n109 0.921
R23378 OUT_P.n282 OUT_P.n281 0.506
R23379 OUT_P.n236 OUT_P.n235 0.506
R23380 OUT_P.n60 OUT_P.n58 0.506
R23381 OUT_P.n106 OUT_P.n104 0.506
R23382 OUT_P.n263 OUT_P.n262 0.476
R23383 OUT_P.n218 OUT_P.n217 0.476
R23384 OUT_P.n84 OUT_P.n83 0.476
R23385 OUT_P.n130 OUT_P.n129 0.476
R23386 OUT_P.n297 OUT_P.n296 0.453
R23387 OUT_P.n253 OUT_P.n252 0.445
R23388 OUT_P.n208 OUT_P.n207 0.445
R23389 OUT_P.n74 OUT_P.n73 0.445
R23390 OUT_P.n120 OUT_P.n119 0.445
R23391 OUT_P.n152 OUT_P.n151 0.414
R23392 OUT_P.n182 OUT_P.n181 0.414
R23393 OUT_P.n51 OUT_P.n50 0.414
R23394 OUT_P.n23 OUT_P.n22 0.414
R23395 OUT_P.n296 OUT_P 0.392
R23396 OUT_P.n164 OUT_P.n163 0.382
R23397 OUT_P.n195 OUT_P.n194 0.382
R23398 OUT_P.n38 OUT_P.n37 0.382
R23399 OUT_P.n10 OUT_P.n9 0.382
R23400 OUT_P.n295 OUT_P.n287 0.216
R23401 OUT_P.n289 OUT_P.n288 0.215
R23402 OUT_P.n304 OUT_P.n303 0.215
R23403 OUT_P.n72 OUT_P.n71 0.073
R23404 OUT_P.n118 OUT_P.n117 0.073
R23405 OUT_P.n261 OUT_P.n260 0.068
R23406 OUT_P.n216 OUT_P.n215 0.068
R23407 OUT_P.n82 OUT_P.n81 0.068
R23408 OUT_P.n128 OUT_P.n127 0.068
R23409 OUT_P.n284 OUT_P.n283 0.055
R23410 OUT_P.n140 OUT_P.n115 0.054
R23411 OUT_P.n94 OUT_P.n69 0.054
R23412 OUT_P.n238 OUT_P.n225 0.054
R23413 OUT_P.n238 OUT_P.n237 0.054
R23414 OUT_P.n94 OUT_P.n93 0.054
R23415 OUT_P.n140 OUT_P.n139 0.054
R23416 OUT_P.n284 OUT_P.n271 0.054
R23417 OUT_P.n264 OUT_P.n261 0.048
R23418 OUT_P.n219 OUT_P.n216 0.048
R23419 OUT_P.n85 OUT_P.n82 0.048
R23420 OUT_P.n131 OUT_P.n128 0.048
R23421 OUT_P.n161 OUT_P.n160 0.046
R23422 OUT_P.n192 OUT_P.n191 0.046
R23423 OUT_P.n35 OUT_P.n34 0.046
R23424 OUT_P.n7 OUT_P.n6 0.046
R23425 OUT_P.n173 OUT_P.n172 0.044
R23426 OUT_P.n203 OUT_P.n202 0.044
R23427 OUT_P.n54 OUT_P.n53 0.044
R23428 OUT_P.n26 OUT_P.n25 0.044
R23429 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN OUT_P.n304 0.043
R23430 OUT_P.n288 OUT_P 0.041
R23431 OUT_P.n254 OUT_P.n251 0.039
R23432 OUT_P.n209 OUT_P.n206 0.039
R23433 OUT_P.n75 OUT_P.n72 0.039
R23434 OUT_P.n121 OUT_P.n118 0.039
R23435 OUT_P.n165 OUT_P.n162 0.038
R23436 OUT_P.n196 OUT_P.n193 0.038
R23437 OUT_P.n39 OUT_P.n36 0.038
R23438 OUT_P.n11 OUT_P.n8 0.038
R23439 OUT_P.n172 OUT_P.n171 0.037
R23440 OUT_P.n202 OUT_P.n201 0.037
R23441 OUT_P.n55 OUT_P.n54 0.037
R23442 OUT_P.n27 OUT_P.n26 0.037
R23443 OUT_P.n230 OUT_P.n228 0.036
R23444 OUT_P.n65 OUT_P.n64 0.036
R23445 OUT_P.n111 OUT_P.n110 0.036
R23446 OUT_P.n276 OUT_P.n274 0.036
R23447 OUT_P.n162 OUT_P.n161 0.034
R23448 OUT_P.n193 OUT_P.n192 0.034
R23449 OUT_P.n36 OUT_P.n35 0.034
R23450 OUT_P.n8 OUT_P.n7 0.034
R23451 OUT_P.n173 OUT_P.n153 0.033
R23452 OUT_P.n203 OUT_P.n183 0.033
R23453 OUT_P.n53 OUT_P.n52 0.033
R23454 OUT_P.n25 OUT_P.n24 0.033
R23455 OUT_P.n268 OUT_P.n266 0.031
R23456 OUT_P.n258 OUT_P.n256 0.031
R23457 OUT_P.n159 OUT_P.n157 0.031
R23458 OUT_P.n222 OUT_P.n220 0.031
R23459 OUT_P.n213 OUT_P.n211 0.031
R23460 OUT_P.n190 OUT_P.n188 0.031
R23461 OUT_P.n33 OUT_P.n31 0.031
R23462 OUT_P.n79 OUT_P.n77 0.031
R23463 OUT_P.n89 OUT_P.n87 0.031
R23464 OUT_P.n5 OUT_P.n3 0.031
R23465 OUT_P.n125 OUT_P.n123 0.031
R23466 OUT_P.n135 OUT_P.n133 0.031
R23467 OUT_P.n170 OUT_P.n168 0.026
R23468 OUT_P.n200 OUT_P.n198 0.026
R23469 OUT_P.n44 OUT_P.n42 0.026
R23470 OUT_P.n16 OUT_P.n14 0.026
R23471 OUT_P.n100 OUT_P.n99 0.024
R23472 OUT_P.n246 OUT_P.n245 0.022
R23473 OUT_P.n283 OUT_P.n279 0.021
R23474 OUT_P.n237 OUT_P.n233 0.021
R23475 OUT_P.n69 OUT_P.n68 0.021
R23476 OUT_P.n115 OUT_P.n114 0.021
R23477 OUT_P.n148 OUT_P.n147 0.019
R23478 OUT_P.n179 OUT_P.n178 0.019
R23479 OUT_P.n47 OUT_P.n46 0.019
R23480 OUT_P.n20 OUT_P.n19 0.019
R23481 OUT_P.n304 OUT_P.n143 0.019
R23482 OUT_P.n279 OUT_P.n278 0.019
R23483 OUT_P.n271 OUT_P.n270 0.019
R23484 OUT_P.n233 OUT_P.n232 0.019
R23485 OUT_P.n225 OUT_P.n224 0.019
R23486 OUT_P.n93 OUT_P.n91 0.019
R23487 OUT_P.n68 OUT_P.n67 0.019
R23488 OUT_P.n139 OUT_P.n137 0.019
R23489 OUT_P.n114 OUT_P.n113 0.019
R23490 OUT_P.n295 OUT_P.n294 0.018
R23491 OUT_P.n298 OUT_P.n297 0.018
R23492 OUT_P.n292 OUT_P.n291 0.016
R23493 OUT_P.n301 OUT_P.n300 0.016
R23494 OUT_P.n278 OUT_P.n276 0.014
R23495 OUT_P.n147 OUT_P.n145 0.014
R23496 OUT_P.n153 OUT_P.n150 0.014
R23497 OUT_P.n232 OUT_P.n230 0.014
R23498 OUT_P.n178 OUT_P.n176 0.014
R23499 OUT_P.n183 OUT_P.n180 0.014
R23500 OUT_P.n52 OUT_P.n49 0.014
R23501 OUT_P.n67 OUT_P.n65 0.014
R23502 OUT_P.n24 OUT_P.n21 0.014
R23503 OUT_P.n113 OUT_P.n111 0.014
R23504 OUT_P.n166 OUT_P.n165 0.013
R23505 OUT_P.n197 OUT_P.n196 0.013
R23506 OUT_P.n40 OUT_P.n39 0.013
R23507 OUT_P.n12 OUT_P.n11 0.013
R23508 OUT_P.n171 OUT_P.n170 0.012
R23509 OUT_P.n201 OUT_P.n200 0.012
R23510 OUT_P.n55 OUT_P.n44 0.012
R23511 OUT_P.n27 OUT_P.n16 0.012
R23512 OUT_P.n260 OUT_P.n258 0.009
R23513 OUT_P.n256 OUT_P.n254 0.009
R23514 OUT_P.n215 OUT_P.n213 0.009
R23515 OUT_P.n211 OUT_P.n209 0.009
R23516 OUT_P.n77 OUT_P.n75 0.009
R23517 OUT_P.n81 OUT_P.n79 0.009
R23518 OUT_P.n123 OUT_P.n121 0.009
R23519 OUT_P.n127 OUT_P.n125 0.009
R23520 OUT_P.n245 OUT_P.n244 0.009
R23521 OUT_P.n101 OUT_P.n100 0.009
R23522 OUT_P.n99 OUT_P.n98 0.008
R23523 OUT_P.n294 OUT_P.n293 0.008
R23524 OUT_P.n290 OUT_P.n289 0.008
R23525 OUT_P.n299 OUT_P.n298 0.008
R23526 OUT_P.n303 OUT_P.n302 0.008
R23527 OUT_P.n247 OUT_P.n246 0.008
R23528 OUT_P.n180 OUT_P.n179 0.007
R23529 OUT_P.n150 OUT_P.n148 0.007
R23530 OUT_P.n49 OUT_P.n47 0.007
R23531 OUT_P.n21 OUT_P.n20 0.007
R23532 OUT_P.n160 OUT_P.n159 0.007
R23533 OUT_P.n191 OUT_P.n190 0.007
R23534 OUT_P.n34 OUT_P.n33 0.007
R23535 OUT_P.n6 OUT_P.n5 0.007
R23536 OUT_P.n31 OUT_P.n29 0.006
R23537 OUT_P.n3 OUT_P.n1 0.006
R23538 OUT_P.n157 OUT_P.n155 0.006
R23539 OUT_P.n188 OUT_P.n187 0.006
R23540 OUT_P.n293 OUT_P.n292 0.005
R23541 OUT_P.n291 OUT_P.n290 0.005
R23542 OUT_P.n300 OUT_P.n299 0.005
R23543 OUT_P.n302 OUT_P.n301 0.005
R23544 OUT_P.n270 OUT_P.n268 0.004
R23545 OUT_P.n266 OUT_P.n264 0.004
R23546 OUT_P.n224 OUT_P.n222 0.004
R23547 OUT_P.n220 OUT_P.n219 0.004
R23548 OUT_P.n286 OUT_P.n285 0.004
R23549 OUT_P.n241 OUT_P.n240 0.004
R23550 OUT_P.n87 OUT_P.n85 0.004
R23551 OUT_P.n91 OUT_P.n89 0.004
R23552 OUT_P.n133 OUT_P.n131 0.004
R23553 OUT_P.n137 OUT_P.n135 0.004
R23554 OUT_P.n95 OUT_P.n57 0.004
R23555 OUT_P.n142 OUT_P.n141 0.004
R23556 OUT_P.n249 OUT_P.n248 0.003
R23557 OUT_P.n97 OUT_P.n96 0.003
R23558 OUT_P.n243 OUT_P.n242 0.003
R23559 OUT_P.n103 OUT_P.n102 0.003
R23560 OUT_P.n248 OUT_P.n247 0.002
R23561 OUT_P.n98 OUT_P.n97 0.002
R23562 OUT_P.n198 OUT_P.n197 0.001
R23563 OUT_P.n168 OUT_P.n166 0.001
R23564 OUT_P.n14 OUT_P.n12 0.001
R23565 OUT_P.n42 OUT_P.n40 0.001
R23566 OUT_P.n244 OUT_P.n243 0.001
R23567 OUT_P.n102 OUT_P.n101 0.001
R23568 OUT_P.n287 OUT_P.n286 0.001
R23569 OUT_P.n285 OUT_P.n249 0.001
R23570 OUT_P.n242 OUT_P.n241 0.001
R23571 OUT_P.n240 OUT_P.n239 0.001
R23572 OUT_P.n57 OUT_P.n56 0.001
R23573 OUT_P.n96 OUT_P.n95 0.001
R23574 OUT_P.n141 OUT_P.n103 0.001
R23575 OUT_P.n143 OUT_P.n142 0.001
C26 VDD GND 11.84fF
C27 m4_2257_876# GND 0.20fF
C28 VBIAS GND 53.84fF
C29 OUT_N GND 12.90fF
C30 IN_N GND 5.57fF
C31 OUT_P GND 11.01fF
C32 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE GND 92.54fF
C33 IN_P GND 5.03fF
C34 OUT_P.n0 GND 0.01fF
C35 OUT_P.n1 GND 0.01fF
C36 OUT_P.n2 GND 0.00fF
C37 OUT_P.n3 GND 0.00fF
C38 OUT_P.n4 GND 0.01fF
C39 OUT_P.n5 GND 0.00fF
C40 OUT_P.n6 GND 0.01fF
C41 OUT_P.n7 GND 0.00fF
C42 OUT_P.n8 GND 0.01fF
C43 OUT_P.n9 GND 0.01fF
C44 OUT_P.n10 GND 0.00fF
C45 OUT_P.n11 GND 0.01fF
C46 OUT_P.n12 GND 0.00fF
C47 OUT_P.n13 GND 0.00fF
C48 OUT_P.n14 GND 0.00fF
C49 OUT_P.n15 GND 0.01fF
C50 OUT_P.n16 GND 0.00fF
C51 OUT_P.n17 GND 0.00fF
C52 OUT_P.n18 GND 0.00fF
C53 OUT_P.n19 GND 0.00fF
C54 OUT_P.n20 GND 0.00fF
C55 OUT_P.n21 GND 0.00fF
C56 OUT_P.n22 GND 0.01fF
C57 OUT_P.n23 GND 0.00fF
C58 OUT_P.n24 GND 0.01fF
C59 OUT_P.n25 GND 0.01fF
C60 OUT_P.n26 GND 0.00fF
C61 OUT_P.n27 GND 0.01fF
C62 OUT_P.n28 GND 0.01fF
C63 OUT_P.n29 GND 0.01fF
C64 OUT_P.n30 GND 0.00fF
C65 OUT_P.n31 GND 0.00fF
C66 OUT_P.n32 GND 0.01fF
C67 OUT_P.n33 GND 0.00fF
C68 OUT_P.n34 GND 0.01fF
C69 OUT_P.n35 GND 0.00fF
C70 OUT_P.n36 GND 0.01fF
C71 OUT_P.n37 GND 0.01fF
C72 OUT_P.n38 GND 0.00fF
C73 OUT_P.n39 GND 0.01fF
C74 OUT_P.n40 GND 0.00fF
C75 OUT_P.n41 GND 0.00fF
C76 OUT_P.n42 GND 0.00fF
C77 OUT_P.n43 GND 0.01fF
C78 OUT_P.n44 GND 0.00fF
C79 OUT_P.n45 GND 0.00fF
C80 OUT_P.n46 GND 0.00fF
C81 OUT_P.n47 GND 0.00fF
C82 OUT_P.n48 GND 0.00fF
C83 OUT_P.n49 GND 0.00fF
C84 OUT_P.n50 GND 0.01fF
C85 OUT_P.n51 GND 0.00fF
C86 OUT_P.n52 GND 0.01fF
C87 OUT_P.n53 GND 0.01fF
C88 OUT_P.n54 GND 0.00fF
C89 OUT_P.n55 GND 0.01fF
C90 OUT_P.n56 GND 1.07fF
C91 OUT_P.n57 GND 0.05fF
C92 OUT_P.n58 GND 0.01fF
C93 OUT_P.n59 GND 0.00fF
C94 OUT_P.n60 GND 0.00fF
C95 OUT_P.n61 GND 0.01fF
C96 OUT_P.t3 GND 0.15fF $ **FLOATING
C97 OUT_P.t4 GND 0.15fF $ **FLOATING
C98 OUT_P.n62 GND 0.43fF
C99 OUT_P.n63 GND 0.06fF
C100 OUT_P.n64 GND 0.33fF
C101 OUT_P.n65 GND 0.01fF
C102 OUT_P.n66 GND 0.00fF
C103 OUT_P.n67 GND 0.00fF
C104 OUT_P.n68 GND 0.00fF
C105 OUT_P.n69 GND 0.01fF
C106 OUT_P.n70 GND 0.01fF
C107 OUT_P.n71 GND 0.01fF
C108 OUT_P.n72 GND 0.01fF
C109 OUT_P.n73 GND 0.01fF
C110 OUT_P.n74 GND 0.00fF
C111 OUT_P.n75 GND 0.01fF
C112 OUT_P.n76 GND 0.00fF
C113 OUT_P.n77 GND 0.00fF
C114 OUT_P.n78 GND 0.00fF
C115 OUT_P.n79 GND 0.00fF
C116 OUT_P.n80 GND 0.01fF
C117 OUT_P.n81 GND 0.01fF
C118 OUT_P.n82 GND 0.01fF
C119 OUT_P.n83 GND 0.01fF
C120 OUT_P.n84 GND 0.00fF
C121 OUT_P.n85 GND 0.01fF
C122 OUT_P.n86 GND 0.00fF
C123 OUT_P.n87 GND 0.00fF
C124 OUT_P.n88 GND 0.00fF
C125 OUT_P.n89 GND 0.00fF
C126 OUT_P.n90 GND 0.00fF
C127 OUT_P.n91 GND 0.00fF
C128 OUT_P.n92 GND 0.01fF
C129 OUT_P.n93 GND 0.01fF
C130 OUT_P.n94 GND 0.01fF
C131 OUT_P.n95 GND 0.05fF
C132 OUT_P.n96 GND 0.05fF
C133 OUT_P.n98 GND 0.12fF
C134 OUT_P.n99 GND 0.23fF
C135 OUT_P.n100 GND 0.24fF
C136 OUT_P.n101 GND 0.12fF
C137 OUT_P.n103 GND 0.05fF
C138 OUT_P.n104 GND 0.01fF
C139 OUT_P.n105 GND 0.00fF
C140 OUT_P.n106 GND 0.00fF
C141 OUT_P.n107 GND 0.01fF
C142 OUT_P.t1 GND 0.15fF $ **FLOATING
C143 OUT_P.t7 GND 0.15fF $ **FLOATING
C144 OUT_P.n108 GND 0.43fF
C145 OUT_P.n109 GND 0.06fF
C146 OUT_P.n110 GND 0.33fF
C147 OUT_P.n111 GND 0.01fF
C148 OUT_P.n112 GND 0.00fF
C149 OUT_P.n113 GND 0.00fF
C150 OUT_P.n114 GND 0.00fF
C151 OUT_P.n115 GND 0.01fF
C152 OUT_P.n116 GND 0.01fF
C153 OUT_P.n117 GND 0.01fF
C154 OUT_P.n118 GND 0.01fF
C155 OUT_P.n119 GND 0.01fF
C156 OUT_P.n120 GND 0.00fF
C157 OUT_P.n121 GND 0.01fF
C158 OUT_P.n122 GND 0.00fF
C159 OUT_P.n123 GND 0.00fF
C160 OUT_P.n124 GND 0.00fF
C161 OUT_P.n125 GND 0.00fF
C162 OUT_P.n126 GND 0.01fF
C163 OUT_P.n127 GND 0.01fF
C164 OUT_P.n128 GND 0.01fF
C165 OUT_P.n129 GND 0.01fF
C166 OUT_P.n130 GND 0.00fF
C167 OUT_P.n131 GND 0.01fF
C168 OUT_P.n132 GND 0.00fF
C169 OUT_P.n133 GND 0.00fF
C170 OUT_P.n134 GND 0.00fF
C171 OUT_P.n135 GND 0.00fF
C172 OUT_P.n136 GND 0.00fF
C173 OUT_P.n137 GND 0.00fF
C174 OUT_P.n138 GND 0.01fF
C175 OUT_P.n139 GND 0.01fF
C176 OUT_P.n140 GND 0.01fF
C177 OUT_P.n141 GND 0.05fF
C178 OUT_P.n142 GND 0.05fF
C179 OUT_P.n143 GND 0.35fF
C180 OUT_P.n144 GND 0.01fF
C181 OUT_P.n145 GND 0.01fF
C182 OUT_P.n146 GND 0.00fF
C183 OUT_P.n147 GND 0.00fF
C184 OUT_P.n148 GND 0.00fF
C185 OUT_P.n149 GND 0.00fF
C186 OUT_P.n150 GND 0.00fF
C187 OUT_P.n151 GND 0.01fF
C188 OUT_P.n152 GND 0.00fF
C189 OUT_P.n153 GND 0.01fF
C190 OUT_P.n154 GND 0.01fF
C191 OUT_P.n155 GND 0.01fF
C192 OUT_P.n156 GND 0.00fF
C193 OUT_P.n157 GND 0.00fF
C194 OUT_P.n158 GND 0.01fF
C195 OUT_P.n159 GND 0.00fF
C196 OUT_P.n160 GND 0.01fF
C197 OUT_P.n161 GND 0.00fF
C198 OUT_P.n162 GND 0.01fF
C199 OUT_P.n163 GND 0.01fF
C200 OUT_P.n164 GND 0.00fF
C201 OUT_P.n165 GND 0.01fF
C202 OUT_P.n166 GND 0.00fF
C203 OUT_P.n167 GND 0.00fF
C204 OUT_P.n168 GND 0.00fF
C205 OUT_P.n169 GND 0.01fF
C206 OUT_P.n170 GND 0.00fF
C207 OUT_P.n171 GND 0.01fF
C208 OUT_P.n172 GND 0.00fF
C209 OUT_P.n173 GND 0.01fF
C210 OUT_P.n174 GND 0.00fF
C211 OUT_P.n175 GND 0.01fF
C212 OUT_P.n176 GND 0.01fF
C213 OUT_P.n177 GND 0.00fF
C214 OUT_P.n178 GND 0.00fF
C215 OUT_P.n179 GND 0.00fF
C216 OUT_P.n180 GND 0.00fF
C217 OUT_P.n181 GND 0.01fF
C218 OUT_P.n182 GND 0.00fF
C219 OUT_P.n183 GND 0.01fF
C220 OUT_P.n184 GND 0.00fF
C221 OUT_P.n185 GND 0.00fF
C222 OUT_P.n186 GND 0.01fF
C223 OUT_P.n187 GND 0.01fF
C224 OUT_P.n188 GND 0.00fF
C225 OUT_P.n189 GND 0.01fF
C226 OUT_P.n190 GND 0.00fF
C227 OUT_P.n191 GND 0.01fF
C228 OUT_P.n192 GND 0.00fF
C229 OUT_P.n193 GND 0.01fF
C230 OUT_P.n194 GND 0.01fF
C231 OUT_P.n195 GND 0.00fF
C232 OUT_P.n196 GND 0.01fF
C233 OUT_P.n197 GND 0.00fF
C234 OUT_P.n198 GND 0.00fF
C235 OUT_P.n199 GND 0.01fF
C236 OUT_P.n200 GND 0.00fF
C237 OUT_P.n201 GND 0.01fF
C238 OUT_P.n202 GND 0.00fF
C239 OUT_P.n203 GND 0.01fF
C240 OUT_P.n204 GND 0.01fF
C241 OUT_P.n205 GND 0.00fF
C242 OUT_P.n206 GND 0.01fF
C243 OUT_P.n207 GND 0.01fF
C244 OUT_P.n208 GND 0.00fF
C245 OUT_P.n209 GND 0.01fF
C246 OUT_P.n210 GND 0.00fF
C247 OUT_P.n211 GND 0.00fF
C248 OUT_P.n212 GND 0.00fF
C249 OUT_P.n213 GND 0.00fF
C250 OUT_P.n214 GND 0.01fF
C251 OUT_P.n215 GND 0.01fF
C252 OUT_P.n216 GND 0.01fF
C253 OUT_P.n217 GND 0.01fF
C254 OUT_P.n218 GND 0.00fF
C255 OUT_P.n219 GND 0.01fF
C256 OUT_P.n220 GND 0.00fF
C257 OUT_P.n221 GND 0.00fF
C258 OUT_P.n222 GND 0.00fF
C259 OUT_P.n223 GND 0.00fF
C260 OUT_P.n224 GND 0.00fF
C261 OUT_P.n225 GND 0.01fF
C262 OUT_P.t6 GND 0.15fF $ **FLOATING
C263 OUT_P.t5 GND 0.15fF $ **FLOATING
C264 OUT_P.n226 GND 0.43fF
C265 OUT_P.n227 GND 0.06fF
C266 OUT_P.n228 GND 0.33fF
C267 OUT_P.n229 GND 0.01fF
C268 OUT_P.n230 GND 0.01fF
C269 OUT_P.n231 GND 0.00fF
C270 OUT_P.n232 GND 0.00fF
C271 OUT_P.n233 GND 0.00fF
C272 OUT_P.n234 GND 0.00fF
C273 OUT_P.n235 GND 0.01fF
C274 OUT_P.n236 GND 0.00fF
C275 OUT_P.n237 GND 0.01fF
C276 OUT_P.n238 GND 0.01fF
C277 OUT_P.n239 GND 0.34fF
C278 OUT_P.n240 GND 0.05fF
C279 OUT_P.n241 GND 0.05fF
C280 OUT_P.n242 GND 0.05fF
C281 OUT_P.n244 GND 0.12fF
C282 OUT_P.n245 GND 0.22fF
C283 OUT_P.n246 GND 0.25fF
C284 OUT_P.n247 GND 0.11fF
C285 OUT_P.n249 GND 0.05fF
C286 OUT_P.n250 GND 0.01fF
C287 OUT_P.n251 GND 0.01fF
C288 OUT_P.n252 GND 0.01fF
C289 OUT_P.n253 GND 0.00fF
C290 OUT_P.n254 GND 0.01fF
C291 OUT_P.n255 GND 0.00fF
C292 OUT_P.n256 GND 0.00fF
C293 OUT_P.n257 GND 0.00fF
C294 OUT_P.n258 GND 0.00fF
C295 OUT_P.n259 GND 0.01fF
C296 OUT_P.n260 GND 0.01fF
C297 OUT_P.n261 GND 0.01fF
C298 OUT_P.n262 GND 0.01fF
C299 OUT_P.n263 GND 0.00fF
C300 OUT_P.n264 GND 0.01fF
C301 OUT_P.n265 GND 0.00fF
C302 OUT_P.n266 GND 0.00fF
C303 OUT_P.n267 GND 0.00fF
C304 OUT_P.n268 GND 0.00fF
C305 OUT_P.n269 GND 0.00fF
C306 OUT_P.n270 GND 0.00fF
C307 OUT_P.n271 GND 0.01fF
C308 OUT_P.t0 GND 0.15fF $ **FLOATING
C309 OUT_P.t2 GND 0.15fF $ **FLOATING
C310 OUT_P.n272 GND 0.43fF
C311 OUT_P.n273 GND 0.06fF
C312 OUT_P.n274 GND 0.33fF
C313 OUT_P.n275 GND 0.01fF
C314 OUT_P.n276 GND 0.01fF
C315 OUT_P.n277 GND 0.00fF
C316 OUT_P.n278 GND 0.00fF
C317 OUT_P.n279 GND 0.00fF
C318 OUT_P.n280 GND 0.00fF
C319 OUT_P.n281 GND 0.01fF
C320 OUT_P.n282 GND 0.00fF
C321 OUT_P.n283 GND 0.01fF
C322 OUT_P.n284 GND 0.01fF
C323 OUT_P.n285 GND 0.05fF
C324 OUT_P.n286 GND 0.05fF
C325 OUT_P.n287 GND 1.07fF
C326 OUT_P.n288 GND 0.43fF
C327 OUT_P.n289 GND 1.84fF
C328 OUT_P.n290 GND 0.06fF
C329 OUT_P.n291 GND 0.11fF
C330 OUT_P.n292 GND 0.11fF
C331 OUT_P.n293 GND 0.06fF
C332 OUT_P.n294 GND 0.18fF
C333 OUT_P.n295 GND 4.48fF
C334 OUT_P.n296 GND 7.96fF
C335 OUT_P.n297 GND 2.08fF
C336 OUT_P.n298 GND 0.18fF
C337 OUT_P.n299 GND 0.06fF
C338 OUT_P.n300 GND 0.11fF
C339 OUT_P.n301 GND 0.11fF
C340 OUT_P.n302 GND 0.06fF
C341 OUT_P.n303 GND 0.50fF
C342 OUT_P.n304 GND 0.35fF
C343 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN GND 0.47fF
C344 IN_P.n0 GND 0.02fF
C345 IN_P.t7 GND 0.28fF $ **FLOATING
C346 IN_P.n1 GND 0.04fF
C347 IN_P.n2 GND 0.17fF
C348 IN_P.n3 GND 0.04fF
C349 IN_P.n4 GND 0.01fF
C350 IN_P.n5 GND 0.02fF
C351 IN_P.t0 GND 0.28fF $ **FLOATING
C352 IN_P.n6 GND 0.04fF
C353 IN_P.n7 GND 0.17fF
C354 IN_P.n8 GND 0.02fF
C355 IN_P.n9 GND 0.04fF
C356 IN_P.n10 GND 0.01fF
C357 IN_P.n11 GND 0.01fF
C358 IN_P.n12 GND 0.01fF
C359 IN_P.n13 GND 0.01fF
C360 IN_P.n14 GND 0.01fF
C361 IN_P.n15 GND 0.01fF
C362 IN_P.n16 GND 0.02fF
C363 IN_P.n17 GND 0.02fF
C364 IN_P.n18 GND 0.01fF
C365 IN_P.n19 GND 0.01fF
C366 IN_P.n20 GND 0.04fF
C367 IN_P.n21 GND 0.06fF
C368 IN_P.n22 GND 0.03fF
C369 IN_P.n23 GND 0.02fF
C370 IN_P.n24 GND 0.01fF
C371 IN_P.n25 GND 0.01fF
C372 IN_P.n26 GND 0.01fF
C373 IN_P.n27 GND 0.00fF
C374 IN_P.n28 GND 0.02fF
C375 IN_P.n29 GND 0.01fF
C376 IN_P.t6 GND 0.28fF $ **FLOATING
C377 IN_P.n30 GND 0.17fF
C378 IN_P.n31 GND 0.02fF
C379 IN_P.n32 GND 0.01fF
C380 IN_P.n33 GND 0.03fF
C381 IN_P.n34 GND 0.00fF
C382 IN_P.n35 GND 0.01fF
C383 IN_P.n36 GND 0.01fF
C384 IN_P.n37 GND 0.01fF
C385 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE GND 0.03fF
C386 IN_P.n38 GND 0.02fF
C387 IN_P.n39 GND 0.02fF
C388 IN_P.n40 GND 0.01fF
C389 IN_P.n41 GND 0.00fF
C390 IN_P.n42 GND 0.01fF
C391 IN_P.n43 GND 0.02fF
C392 IN_P.n44 GND 0.04fF
C393 IN_P.t4 GND 0.28fF $ **FLOATING
C394 IN_P.n45 GND 0.17fF
C395 IN_P.n46 GND 0.02fF
C396 IN_P.n47 GND 0.02fF
C397 IN_P.n48 GND 0.03fF
C398 IN_P.n49 GND 0.01fF
C399 IN_P.n50 GND 0.00fF
C400 IN_P.n51 GND 0.01fF
C401 IN_P.n52 GND 0.03fF
C402 IN_P.n53 GND 0.02fF
C403 IN_P.n54 GND 0.02fF
C404 IN_P.n55 GND 0.00fF
C405 IN_P.n56 GND 0.01fF
C406 IN_P.n57 GND 0.01fF
C407 IN_P.n58 GND 0.01fF
C408 IN_P.n59 GND 0.02fF
C409 IN_P.n60 GND 0.01fF
C410 IN_P.t3 GND 0.28fF $ **FLOATING
C411 IN_P.n61 GND 0.17fF
C412 IN_P.n62 GND 0.02fF
C413 IN_P.n63 GND 0.01fF
C414 IN_P.n64 GND 0.03fF
C415 IN_P.n65 GND 0.00fF
C416 IN_P.n66 GND 0.01fF
C417 IN_P.n67 GND 0.01fF
C418 IN_P.n68 GND 0.02fF
C419 IN_P.n69 GND 0.01fF
C420 IN_P.n70 GND 0.00fF
C421 IN_P.n71 GND 0.05fF
C422 IN_P.n72 GND 0.03fF
C423 IN_P.n73 GND 0.01fF
C424 IN_P.n74 GND 0.03fF
C425 IN_P.n75 GND 0.02fF
C426 IN_P.n76 GND 0.01fF
C427 IN_P.n77 GND 0.01fF
C428 IN_P.n78 GND 0.01fF
C429 IN_P.n79 GND 0.01fF
C430 IN_P.n80 GND 0.01fF
C431 IN_P.n81 GND 0.01fF
C432 IN_P.n82 GND 0.01fF
C433 IN_P.n83 GND 0.02fF
C434 IN_P.n84 GND 0.02fF
C435 IN_P.n85 GND 0.02fF
C436 IN_P.n86 GND 0.23fF
C437 IN_P.n87 GND 0.02fF
C438 IN_P.n88 GND 0.04fF
C439 IN_P.n89 GND 0.17fF
C440 IN_P.n90 GND 0.03fF
C441 IN_P.n91 GND 0.06fF
C442 IN_P.n92 GND 0.02fF
C443 IN_P.n93 GND 0.01fF
C444 IN_P.n94 GND 0.01fF
C445 IN_P.n95 GND 0.00fF
C446 IN_P.n96 GND 0.00fF
C447 IN_P.n97 GND 0.04fF
C448 IN_P.n98 GND 0.15fF
C449 IN_P.n99 GND 0.04fF
C450 IN_P.n100 GND 0.02fF
C451 IN_P.n101 GND 0.05fF
C452 IN_P.n102 GND 0.01fF
C453 IN_P.n103 GND 0.01fF
C454 IN_P.n104 GND 0.09fF
C455 IN_P.n105 GND 0.01fF
C456 IN_P.n106 GND 0.01fF
C457 IN_P.n107 GND 0.02fF
C458 IN_P.n108 GND 0.03fF
C459 IN_P.n109 GND 0.02fF
C460 IN_P.n110 GND 0.01fF
C461 IN_P.n111 GND 0.03fF
C462 IN_P.n112 GND 0.02fF
C463 IN_P.n113 GND 0.02fF
C464 IN_P.n114 GND 0.00fF
C465 IN_P.n115 GND 0.01fF
C466 IN_P.n116 GND 0.01fF
C467 IN_P.n117 GND 0.01fF
C468 IN_P.n118 GND 0.02fF
C469 IN_P.n119 GND 0.01fF
C470 IN_P.n120 GND 0.17fF
C471 IN_P.n121 GND 0.02fF
C472 IN_P.n122 GND 0.01fF
C473 IN_P.n123 GND 0.03fF
C474 IN_P.n124 GND 0.00fF
C475 IN_P.n125 GND 0.01fF
C476 IN_P.n126 GND 0.01fF
C477 IN_P.n127 GND 0.02fF
C478 IN_P.n128 GND 0.01fF
C479 IN_P.n129 GND 0.01fF
C480 IN_P.n130 GND 0.01fF
C481 IN_P.n131 GND 0.05fF
C482 IN_P.n132 GND 0.03fF
C483 IN_P.n133 GND 0.01fF
C484 IN_P.n134 GND 0.01fF
C485 IN_P.n135 GND 0.02fF
C486 IN_P.n136 GND 0.00fF
C487 IN_P.n137 GND 0.01fF
C488 IN_P.n138 GND 0.02fF
C489 IN_P.n139 GND 0.02fF
C490 IN_P.n140 GND 0.01fF
C491 IN_P.n141 GND 0.02fF
C492 IN_P.n142 GND 0.01fF
C493 IN_P.n143 GND 0.17fF
C494 IN_P.n144 GND 0.02fF
C495 IN_P.n145 GND 0.01fF
C496 IN_P.n146 GND 0.03fF
C497 IN_P.n147 GND 0.01fF
C498 IN_P.n148 GND 0.01fF
C499 IN_P.n149 GND 0.01fF
C500 IN_P.n150 GND 0.02fF
C501 IN_P.n151 GND 0.01fF
C502 IN_P.n152 GND 0.01fF
C503 IN_P.n153 GND 0.02fF
C504 IN_P.n154 GND 0.01fF
C505 IN_P.n155 GND 0.01fF
C506 IN_P.n156 GND 0.02fF
C507 IN_P.n157 GND 0.02fF
C508 IN_P.n158 GND 0.02fF
C509 IN_P.n159 GND 0.02fF
C510 IN_P.n160 GND 0.01fF
C511 IN_P.n161 GND 0.02fF
C512 IN_P.n162 GND 0.01fF
C513 IN_P.n163 GND 0.01fF
C514 IN_P.n164 GND 0.02fF
C515 IN_P.n165 GND 0.01fF
C516 IN_P.n166 GND 0.01fF
C517 IN_P.n167 GND 0.02fF
C518 IN_P.n168 GND 0.02fF
C519 IN_P.n169 GND 0.02fF
C520 IN_P.n170 GND 0.02fF
C521 IN_P.n171 GND 0.09fF
C522 IN_P.n172 GND 0.11fF
C523 IN_P.n173 GND 0.04fF
C524 IN_P.n174 GND 0.01fF
C525 IN_P.n175 GND 0.01fF
C526 IN_P.n176 GND 0.03fF
C527 IN_P.n177 GND 0.03fF
C528 IN_P.n178 GND 0.01fF
C529 IN_P.n179 GND 0.01fF
C530 IN_P.n180 GND 0.04fF
C531 IN_P.n181 GND 0.04fF
C532 IN_P.n182 GND 0.02fF
C533 IN_P.n183 GND 0.98fF
C534 IN_P.n184 GND 0.02fF
C535 IN_P.n185 GND 0.04fF
C536 IN_P.n186 GND 0.17fF
C537 IN_P.n187 GND 0.03fF
C538 IN_P.n188 GND 0.06fF
C539 IN_P.n189 GND 0.02fF
C540 IN_P.n190 GND 0.01fF
C541 IN_P.n191 GND 0.01fF
C542 IN_P.n192 GND 0.00fF
C543 IN_P.n193 GND 0.00fF
C544 IN_P.n194 GND 0.04fF
C545 IN_P.n195 GND 0.15fF
C546 IN_P.n196 GND 0.04fF
C547 IN_P.n197 GND 0.02fF
C548 IN_P.n198 GND 0.05fF
C549 IN_P.n199 GND 0.01fF
C550 IN_P.n200 GND 0.01fF
C551 IN_P.n201 GND 0.09fF
C552 IN_P.n202 GND 0.01fF
C553 IN_P.n203 GND 0.01fF
C554 IN_P.n204 GND 0.02fF
C555 IN_P.n205 GND 0.03fF
C556 IN_P.n206 GND 0.02fF
C557 IN_P.n207 GND 0.01fF
C558 IN_P.n208 GND 0.03fF
C559 IN_P.n209 GND 0.02fF
C560 IN_P.n210 GND 0.02fF
C561 IN_P.n211 GND 0.00fF
C562 IN_P.n212 GND 0.01fF
C563 IN_P.n213 GND 0.01fF
C564 IN_P.n214 GND 0.01fF
C565 IN_P.n215 GND 0.02fF
C566 IN_P.n216 GND 0.01fF
C567 IN_P.n217 GND 0.17fF
C568 IN_P.n218 GND 0.02fF
C569 IN_P.n219 GND 0.01fF
C570 IN_P.n220 GND 0.03fF
C571 IN_P.n221 GND 0.00fF
C572 IN_P.n222 GND 0.01fF
C573 IN_P.n223 GND 0.01fF
C574 IN_P.n224 GND 0.02fF
C575 IN_P.n225 GND 0.01fF
C576 IN_P.n226 GND 0.01fF
C577 IN_P.n227 GND 0.01fF
C578 IN_P.n228 GND 0.05fF
C579 IN_P.n229 GND 0.03fF
C580 IN_P.n230 GND 0.01fF
C581 IN_P.n231 GND 0.01fF
C582 IN_P.n232 GND 0.02fF
C583 IN_P.n233 GND 0.00fF
C584 IN_P.n234 GND 0.01fF
C585 IN_P.n235 GND 0.02fF
C586 IN_P.n236 GND 0.02fF
C587 IN_P.n237 GND 0.01fF
C588 IN_P.n238 GND 0.02fF
C589 IN_P.n239 GND 0.01fF
C590 IN_P.n240 GND 0.17fF
C591 IN_P.n241 GND 0.02fF
C592 IN_P.n242 GND 0.01fF
C593 IN_P.n243 GND 0.03fF
C594 IN_P.n244 GND 0.01fF
C595 IN_P.n245 GND 0.01fF
C596 IN_P.n246 GND 0.01fF
C597 IN_P.n247 GND 0.02fF
C598 IN_P.n248 GND 0.01fF
C599 IN_P.n249 GND 0.01fF
C600 IN_P.n250 GND 0.02fF
C601 IN_P.n251 GND 0.01fF
C602 IN_P.n252 GND 0.01fF
C603 IN_P.n253 GND 0.02fF
C604 IN_P.n254 GND 0.02fF
C605 IN_P.n255 GND 0.02fF
C606 IN_P.n256 GND 0.02fF
C607 IN_P.n257 GND 0.01fF
C608 IN_P.n258 GND 0.02fF
C609 IN_P.n259 GND 0.01fF
C610 IN_P.n260 GND 0.01fF
C611 IN_P.n261 GND 0.02fF
C612 IN_P.n262 GND 0.01fF
C613 IN_P.n263 GND 0.01fF
C614 IN_P.n264 GND 0.02fF
C615 IN_P.n265 GND 0.02fF
C616 IN_P.n266 GND 0.02fF
C617 IN_P.n267 GND 0.02fF
C618 IN_P.n268 GND 0.09fF
C619 IN_P.n269 GND 0.33fF
C620 IN_P.n270 GND 0.10fF
C621 IN_P.n271 GND 0.04fF
C622 IN_P.n272 GND 0.04fF
C623 IN_P.n273 GND 0.09fF
C624 IN_P.n274 GND 0.09fF
C625 IN_P.n275 GND 0.04fF
C626 IN_P.n276 GND 0.04fF
C627 IN_P.n277 GND 0.10fF
C628 IN_P.n278 GND 0.12fF
C629 IN_P.n279 GND 0.05fF
C630 IN_P.n280 GND 1.93fF
C631 IN_P.n281 GND 1.92fF
C632 IN_P.n282 GND 1.41fF
C633 IN_P.n283 GND 0.37fF
C634 IN_P.n284 GND 0.31fF
C635 IN_P.n285 GND 0.02fF
C636 IN_P.n286 GND 0.05fF
C637 IN_P.n287 GND 0.04fF
C638 IN_P.n288 GND 0.01fF
C639 IN_P.n289 GND 0.01fF
C640 IN_P.n290 GND 0.03fF
C641 IN_P.n291 GND 0.03fF
C642 IN_P.n292 GND 0.01fF
C643 IN_P.n293 GND 0.01fF
C644 IN_P.n294 GND 0.04fF
C645 IN_P.n295 GND 0.01fF
C646 IN_P.n296 GND 0.01fF
C647 IN_P.n297 GND 0.00fF
C648 IN_P.n298 GND 0.00fF
C649 IN_P.n299 GND 0.01fF
C650 IN_P.n300 GND 0.32fF
C651 IN_P.n301 GND 0.32fF
C652 IN_P.n302 GND 0.01fF
C653 IN_P.n303 GND 0.01fF
C654 IN_P.n304 GND 0.03fF
C655 IN_P.n305 GND 0.03fF
C656 IN_P.n306 GND 0.01fF
C657 IN_P.n307 GND 0.01fF
C658 IN_P.n308 GND 0.03fF
C659 IN_P.n309 GND 0.03fF
C660 IN_P.n310 GND 0.01fF
C661 IN_P.n311 GND 0.01fF
C662 IN_P.n312 GND 0.03fF
C663 IN_P.n313 GND 0.03fF
C664 IN_P.n314 GND 0.01fF
C665 IN_P.n315 GND 0.11fF
C666 IN_P.n316 GND 0.08fF
C667 IN_P.n317 GND 0.02fF
C668 IN_P.n318 GND 0.04fF
C669 IN_P.n319 GND 0.01fF
C670 IN_P.n320 GND 0.01fF
C671 IN_P.n321 GND 0.02fF
C672 IN_P.n322 GND 0.01fF
C673 IN_P.t5 GND 0.28fF $ **FLOATING
C674 IN_P.n323 GND 0.17fF
C675 IN_P.n324 GND 0.02fF
C676 IN_P.n325 GND 0.01fF
C677 IN_P.n326 GND 0.03fF
C678 IN_P.n327 GND 0.00fF
C679 IN_P.n328 GND 0.01fF
C680 IN_P.n329 GND 0.03fF
C681 IN_P.n330 GND 0.03fF
C682 IN_P.n331 GND 0.05fF
C683 IN_P.n332 GND 0.03fF
C684 IN_P.n333 GND 0.01fF
C685 IN_P.n334 GND 0.01fF
C686 IN_P.n335 GND 0.02fF
C687 IN_P.n336 GND 0.02fF
C688 IN_P.t2 GND 0.28fF $ **FLOATING
C689 IN_P.n337 GND 0.04fF
C690 IN_P.n338 GND 0.17fF
C691 IN_P.n339 GND 0.02fF
C692 IN_P.n340 GND 0.02fF
C693 IN_P.n341 GND 0.03fF
C694 IN_P.n342 GND 0.01fF
C695 IN_P.n343 GND 0.01fF
C696 IN_P.n344 GND 0.03fF
C697 IN_P.n345 GND 0.02fF
C698 IN_P.n346 GND 0.02fF
C699 IN_P.n347 GND 0.01fF
C700 IN_P.n348 GND 0.01fF
C701 IN_P.n349 GND 0.01fF
C702 IN_P.n350 GND 0.00fF
C703 IN_P.n351 GND 0.02fF
C704 IN_P.n352 GND 0.01fF
C705 IN_P.t1 GND 0.28fF $ **FLOATING
C706 IN_P.n353 GND 0.17fF
C707 IN_P.n354 GND 0.02fF
C708 IN_P.n355 GND 0.01fF
C709 IN_P.n356 GND 0.03fF
C710 IN_P.n357 GND 0.00fF
C711 IN_P.n358 GND 0.01fF
C712 IN_P.n359 GND 0.02fF
C713 OUT_N.n0 GND 0.00fF
C714 OUT_N.n1 GND 0.01fF
C715 OUT_N.n2 GND 0.00fF
C716 OUT_N.n3 GND 0.01fF
C717 OUT_N.n4 GND 0.01fF
C718 OUT_N.n5 GND 0.01fF
C719 OUT_N.n6 GND 0.01fF
C720 OUT_N.n7 GND 0.01fF
C721 OUT_N.t7 GND 0.16fF $ **FLOATING
C722 OUT_N.n8 GND 0.01fF
C723 OUT_N.t1 GND 0.16fF $ **FLOATING
C724 OUT_N.n9 GND 0.46fF
C725 OUT_N.n10 GND 0.04fF
C726 OUT_N.n11 GND 0.37fF
C727 OUT_N.n12 GND 0.01fF
C728 OUT_N.n13 GND 0.01fF
C729 OUT_N.n14 GND 0.00fF
C730 OUT_N.n15 GND 0.00fF
C731 OUT_N.n16 GND 0.00fF
C732 OUT_N.n17 GND 0.01fF
C733 OUT_N.n19 GND 0.38fF
C734 OUT_N.n20 GND 0.06fF
C735 OUT_N.n21 GND 0.06fF
C736 OUT_N.n22 GND 0.06fF
C737 OUT_N.n23 GND 0.00fF
C738 OUT_N.n24 GND 0.00fF
C739 OUT_N.n25 GND 0.00fF
C740 OUT_N.n26 GND 0.00fF
C741 OUT_N.n27 GND 0.00fF
C742 OUT_N.n28 GND 0.00fF
C743 OUT_N.n29 GND 0.00fF
C744 OUT_N.n30 GND 0.00fF
C745 OUT_N.n31 GND 0.00fF
C746 OUT_N.n32 GND 0.01fF
C747 OUT_N.n33 GND 0.02fF
C748 OUT_N.n34 GND 0.00fF
C749 OUT_N.n35 GND 0.00fF
C750 OUT_N.n36 GND 0.00fF
C751 OUT_N.n37 GND 0.01fF
C752 OUT_N.n38 GND 0.01fF
C753 OUT_N.n39 GND 0.01fF
C754 OUT_N.n40 GND 0.00fF
C755 OUT_N.n41 GND 0.01fF
C756 OUT_N.n42 GND 0.00fF
C757 OUT_N.n43 GND 0.00fF
C758 OUT_N.n44 GND 0.01fF
C759 OUT_N.n45 GND 0.01fF
C760 OUT_N.n46 GND 0.01fF
C761 OUT_N.n47 GND 0.01fF
C762 OUT_N.n48 GND 0.00fF
C763 OUT_N.n49 GND 0.01fF
C764 OUT_N.n50 GND 0.00fF
C765 OUT_N.n51 GND 0.00fF
C766 OUT_N.n52 GND 0.00fF
C767 OUT_N.n53 GND 0.01fF
C768 OUT_N.n54 GND 0.01fF
C769 OUT_N.n55 GND 0.01fF
C770 OUT_N.n56 GND 0.01fF
C771 OUT_N.n57 GND 0.00fF
C772 OUT_N.n58 GND 0.01fF
C773 OUT_N.n59 GND 0.00fF
C774 OUT_N.n60 GND 0.00fF
C775 OUT_N.n61 GND 0.00fF
C776 OUT_N.n62 GND 0.01fF
C777 OUT_N.n63 GND 0.01fF
C778 OUT_N.n64 GND 0.01fF
C779 OUT_N.n65 GND 0.01fF
C780 OUT_N.n66 GND 0.00fF
C781 OUT_N.n67 GND 0.01fF
C782 OUT_N.n68 GND 0.00fF
C783 OUT_N.t4 GND 0.16fF $ **FLOATING
C784 OUT_N.n70 GND 0.01fF
C785 OUT_N.t5 GND 0.16fF $ **FLOATING
C786 OUT_N.n71 GND 0.46fF
C787 OUT_N.n72 GND 0.04fF
C788 OUT_N.n73 GND 0.37fF
C789 OUT_N.n74 GND 0.01fF
C790 OUT_N.n75 GND 0.01fF
C791 OUT_N.n76 GND 0.00fF
C792 OUT_N.n77 GND 0.01fF
C793 OUT_N.n78 GND 0.00fF
C794 OUT_N.n79 GND 0.01fF
C795 OUT_N.n80 GND 0.00fF
C796 OUT_N.n81 GND 0.00fF
C797 OUT_N.n82 GND 0.00fF
C798 OUT_N.n83 GND 0.01fF
C799 OUT_N.n85 GND 0.01fF
C800 OUT_N.n86 GND 0.01fF
C801 OUT_N.n87 GND 0.01fF
C802 OUT_N.n88 GND 0.01fF
C803 OUT_N.n90 GND 0.12fF
C804 OUT_N.n91 GND 0.27fF
C805 OUT_N.n92 GND 0.25fF
C806 OUT_N.n93 GND 0.00fF
C807 OUT_N.n94 GND 0.00fF
C808 OUT_N.n95 GND 0.00fF
C809 OUT_N.n96 GND 0.00fF
C810 OUT_N.n97 GND 0.00fF
C811 OUT_N.n98 GND 0.00fF
C812 OUT_N.n99 GND 0.00fF
C813 OUT_N.n100 GND 0.00fF
C814 OUT_N.n101 GND 0.00fF
C815 OUT_N.n102 GND 0.01fF
C816 OUT_N.n103 GND 0.02fF
C817 OUT_N.n104 GND 0.00fF
C818 OUT_N.n105 GND 0.00fF
C819 OUT_N.n106 GND 0.01fF
C820 OUT_N.n107 GND 0.01fF
C821 OUT_N.n108 GND 0.01fF
C822 OUT_N.n109 GND 0.00fF
C823 OUT_N.n110 GND 0.01fF
C824 OUT_N.n111 GND 0.00fF
C825 OUT_N.n112 GND 0.00fF
C826 OUT_N.n113 GND 0.01fF
C827 OUT_N.n114 GND 0.01fF
C828 OUT_N.n115 GND 0.01fF
C829 OUT_N.n116 GND 0.01fF
C830 OUT_N.n117 GND 0.00fF
C831 OUT_N.n118 GND 0.01fF
C832 OUT_N.n119 GND 0.00fF
C833 OUT_N.n120 GND 0.00fF
C834 OUT_N.n121 GND 0.00fF
C835 OUT_N.n122 GND 0.01fF
C836 OUT_N.n123 GND 0.01fF
C837 OUT_N.n124 GND 0.01fF
C838 OUT_N.n125 GND 0.01fF
C839 OUT_N.n126 GND 0.00fF
C840 OUT_N.n127 GND 0.01fF
C841 OUT_N.n128 GND 0.00fF
C842 OUT_N.n129 GND 0.00fF
C843 OUT_N.n130 GND 0.00fF
C844 OUT_N.n131 GND 0.01fF
C845 OUT_N.n132 GND 0.01fF
C846 OUT_N.n133 GND 0.01fF
C847 OUT_N.n134 GND 0.01fF
C848 OUT_N.n135 GND 0.00fF
C849 OUT_N.n136 GND 0.01fF
C850 OUT_N.n137 GND 0.00fF
C851 OUT_N.n138 GND 0.00fF
C852 OUT_N.n140 GND 0.12fF
C853 OUT_N.n142 GND 0.06fF
C854 OUT_N.n143 GND 0.06fF
C855 OUT_N.n144 GND 0.06fF
C856 OUT_N.n145 GND 1.17fF
C857 OUT_N.n146 GND 0.39fF
C858 OUT_N.n147 GND 0.54fF
C859 OUT_N.n148 GND 0.07fF
C860 OUT_N.n149 GND 0.12fF
C861 OUT_N.n150 GND 0.12fF
C862 OUT_N.n151 GND 0.07fF
C863 OUT_N.n152 GND 0.20fF
C864 OUT_N.n153 GND 1.96fF
C865 OUT_N.n154 GND 7.87fF
C866 OUT_N.n155 GND 3.91fF
C867 OUT_N.n156 GND 0.20fF
C868 OUT_N.n157 GND 0.07fF
C869 OUT_N.n158 GND 0.12fF
C870 OUT_N.n159 GND 0.12fF
C871 OUT_N.n160 GND 0.07fF
C872 OUT_N.n161 GND 2.00fF
C873 OUT_N.n162 GND 0.01fF
C874 OUT_N.n163 GND 0.00fF
C875 OUT_N.n164 GND 0.00fF
C876 OUT_N.n165 GND 0.01fF
C877 OUT_N.n166 GND 0.00fF
C878 OUT_N.n167 GND 0.00fF
C879 OUT_N.n168 GND 0.00fF
C880 OUT_N.n169 GND 0.01fF
C881 OUT_N.n170 GND 0.01fF
C882 OUT_N.t2 GND 0.16fF $ **FLOATING
C883 OUT_N.n171 GND 0.01fF
C884 OUT_N.t6 GND 0.16fF $ **FLOATING
C885 OUT_N.n172 GND 0.46fF
C886 OUT_N.n173 GND 0.04fF
C887 OUT_N.n174 GND 0.37fF
C888 OUT_N.n175 GND 0.01fF
C889 OUT_N.n177 GND 0.00fF
C890 OUT_N.n178 GND 0.00fF
C891 OUT_N.n179 GND 0.00fF
C892 OUT_N.n180 GND 0.00fF
C893 OUT_N.n181 GND 0.00fF
C894 OUT_N.n182 GND 0.01fF
C895 OUT_N.n183 GND 0.02fF
C896 OUT_N.n184 GND 0.00fF
C897 OUT_N.n185 GND 0.00fF
C898 OUT_N.n186 GND 0.00fF
C899 OUT_N.n187 GND 0.01fF
C900 OUT_N.n188 GND 0.01fF
C901 OUT_N.n189 GND 0.01fF
C902 OUT_N.n190 GND 0.00fF
C903 OUT_N.n191 GND 0.01fF
C904 OUT_N.n192 GND 0.00fF
C905 OUT_N.n193 GND 0.00fF
C906 OUT_N.n194 GND 0.00fF
C907 OUT_N.n195 GND 0.01fF
C908 OUT_N.n196 GND 0.01fF
C909 OUT_N.n197 GND 0.01fF
C910 OUT_N.n198 GND 0.01fF
C911 OUT_N.n199 GND 0.00fF
C912 OUT_N.n200 GND 0.01fF
C913 OUT_N.n201 GND 0.00fF
C914 OUT_N.n202 GND 0.00fF
C915 OUT_N.n203 GND 0.00fF
C916 OUT_N.n204 GND 0.00fF
C917 OUT_N.n205 GND 0.01fF
C918 OUT_N.n206 GND 0.01fF
C919 OUT_N.n207 GND 0.01fF
C920 OUT_N.n208 GND 0.01fF
C921 OUT_N.n209 GND 0.00fF
C922 OUT_N.n210 GND 0.01fF
C923 OUT_N.n211 GND 0.00fF
C924 OUT_N.n212 GND 0.00fF
C925 OUT_N.n213 GND 0.00fF
C926 OUT_N.n214 GND 0.00fF
C927 OUT_N.n215 GND 0.01fF
C928 OUT_N.n216 GND 0.01fF
C929 OUT_N.n217 GND 0.01fF
C930 OUT_N.n218 GND 0.01fF
C931 OUT_N.n219 GND 0.00fF
C932 OUT_N.n220 GND 0.01fF
C933 OUT_N.n221 GND 0.00fF
C934 OUT_N.n222 GND 0.00fF
C935 OUT_N.n224 GND 0.01fF
C936 OUT_N.n225 GND 0.00fF
C937 OUT_N.n226 GND 0.00fF
C938 OUT_N.n227 GND 0.01fF
C939 OUT_N.n228 GND 0.01fF
C940 OUT_N.n229 GND 0.01fF
C941 OUT_N.n230 GND 0.01fF
C942 OUT_N.n231 GND 0.01fF
C943 OUT_N.n233 GND 0.00fF
C944 OUT_N.n234 GND 0.00fF
C945 OUT_N.n235 GND 0.00fF
C946 OUT_N.n236 GND 0.01fF
C947 OUT_N.n237 GND 0.01fF
C948 OUT_N.t3 GND 0.16fF $ **FLOATING
C949 OUT_N.n238 GND 0.01fF
C950 OUT_N.t0 GND 0.16fF $ **FLOATING
C951 OUT_N.n239 GND 0.46fF
C952 OUT_N.n240 GND 0.04fF
C953 OUT_N.n241 GND 0.37fF
C954 OUT_N.n242 GND 0.01fF
C955 OUT_N.n243 GND 1.17fF
C956 OUT_N.n244 GND 0.06fF
C957 OUT_N.n245 GND 0.06fF
C958 OUT_N.n246 GND 0.06fF
C959 OUT_N.n248 GND 0.12fF
C960 OUT_N.n249 GND 0.26fF
C961 OUT_N.n250 GND 0.26fF
C962 OUT_N.n251 GND 0.01fF
C963 OUT_N.n252 GND 0.02fF
C964 OUT_N.n253 GND 0.00fF
C965 OUT_N.n254 GND 0.00fF
C966 OUT_N.n255 GND 0.00fF
C967 OUT_N.n256 GND 0.01fF
C968 OUT_N.n257 GND 0.01fF
C969 OUT_N.n258 GND 0.01fF
C970 OUT_N.n259 GND 0.00fF
C971 OUT_N.n260 GND 0.01fF
C972 OUT_N.n261 GND 0.00fF
C973 OUT_N.n262 GND 0.00fF
C974 OUT_N.n263 GND 0.00fF
C975 OUT_N.n264 GND 0.01fF
C976 OUT_N.n265 GND 0.01fF
C977 OUT_N.n266 GND 0.01fF
C978 OUT_N.n267 GND 0.01fF
C979 OUT_N.n268 GND 0.00fF
C980 OUT_N.n269 GND 0.01fF
C981 OUT_N.n270 GND 0.00fF
C982 OUT_N.n271 GND 0.00fF
C983 OUT_N.n272 GND 0.00fF
C984 OUT_N.n273 GND 0.00fF
C985 OUT_N.n274 GND 0.01fF
C986 OUT_N.n275 GND 0.01fF
C987 OUT_N.n276 GND 0.01fF
C988 OUT_N.n277 GND 0.01fF
C989 OUT_N.n278 GND 0.00fF
C990 OUT_N.n279 GND 0.01fF
C991 OUT_N.n280 GND 0.00fF
C992 OUT_N.n281 GND 0.00fF
C993 OUT_N.n282 GND 0.00fF
C994 OUT_N.n283 GND 0.00fF
C995 OUT_N.n284 GND 0.01fF
C996 OUT_N.n285 GND 0.01fF
C997 OUT_N.n286 GND 0.01fF
C998 OUT_N.n287 GND 0.01fF
C999 OUT_N.n288 GND 0.00fF
C1000 OUT_N.n289 GND 0.01fF
C1001 OUT_N.n290 GND 0.00fF
C1002 OUT_N.n291 GND 0.00fF
C1003 OUT_N.n292 GND 0.00fF
C1004 OUT_N.n293 GND 0.00fF
C1005 OUT_N.n294 GND 0.00fF
C1006 OUT_N.n295 GND 0.00fF
C1007 OUT_N.n296 GND 0.00fF
C1008 OUT_N.n298 GND 0.01fF
C1009 OUT_N.n299 GND 0.01fF
C1010 OUT_N.n300 GND 0.01fF
C1011 OUT_N.n301 GND 0.01fF
C1012 OUT_N.n303 GND 0.12fF
C1013 OUT_N.n304 GND 0.06fF
C1014 OUT_N.n305 GND 0.06fF
C1015 OUT_N.n306 GND 0.06fF
C1016 OUT_N.n307 GND 0.39fF
C1017 OUT_N.n308 GND 0.46fF
C1018 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN GND 0.55fF
C1019 IN_N.n0 GND 0.02fF
C1020 IN_N.t4 GND 0.27fF $ **FLOATING
C1021 IN_N.n1 GND 0.04fF
C1022 IN_N.n2 GND 0.17fF
C1023 IN_N.n3 GND 0.03fF
C1024 IN_N.n4 GND 0.01fF
C1025 IN_N.n5 GND 0.01fF
C1026 IN_N.n6 GND 0.01fF
C1027 IN_N.n7 GND 0.01fF
C1028 IN_N.n8 GND 0.01fF
C1029 IN_N.n9 GND 0.01fF
C1030 IN_N.n10 GND 0.02fF
C1031 IN_N.n11 GND 0.02fF
C1032 IN_N.n12 GND 0.02fF
C1033 IN_N.n13 GND 0.05fF
C1034 IN_N.n14 GND 0.02fF
C1035 IN_N.n15 GND 0.02fF
C1036 IN_N.t2 GND 0.27fF $ **FLOATING
C1037 IN_N.n16 GND 0.04fF
C1038 IN_N.n17 GND 0.17fF
C1039 IN_N.n18 GND 0.03fF
C1040 IN_N.n19 GND 0.02fF
C1041 IN_N.n20 GND 0.01fF
C1042 IN_N.n21 GND 0.04fF
C1043 IN_N.n22 GND 0.01fF
C1044 IN_N.n23 GND 0.01fF
C1045 IN_N.n24 GND 0.01fF
C1046 IN_N.n25 GND 0.01fF
C1047 IN_N.n26 GND 0.01fF
C1048 IN_N.n27 GND 0.00fF
C1049 IN_N.n28 GND 0.01fF
C1050 IN_N.n29 GND 0.02fF
C1051 IN_N.n30 GND 0.01fF
C1052 IN_N.n31 GND 0.01fF
C1053 IN_N.n32 GND 0.01fF
C1054 IN_N.n33 GND 0.01fF
C1055 IN_N.n34 GND 0.03fF
C1056 IN_N.n35 GND 0.03fF
C1057 IN_N.n36 GND 0.01fF
C1058 IN_N.n37 GND 0.02fF
C1059 IN_N.n38 GND 0.01fF
C1060 IN_N.n39 GND 0.01fF
C1061 IN_N.n40 GND 0.01fF
C1062 IN_N.n41 GND 0.01fF
C1063 IN_N.n42 GND 0.01fF
C1064 IN_N.n43 GND 0.01fF
C1065 IN_N.n44 GND 0.01fF
C1066 IN_N.n45 GND 0.01fF
C1067 IN_N.n46 GND 0.01fF
C1068 IN_N.n47 GND 0.04fF
C1069 IN_N.n48 GND 0.04fF
C1070 IN_N.n49 GND 0.02fF
C1071 IN_N.n50 GND 0.04fF
C1072 IN_N.n51 GND 0.17fF
C1073 IN_N.n52 GND 0.03fF
C1074 IN_N.n53 GND 0.06fF
C1075 IN_N.n54 GND 0.02fF
C1076 IN_N.n55 GND 0.01fF
C1077 IN_N.n56 GND 0.01fF
C1078 IN_N.n57 GND 0.00fF
C1079 IN_N.n58 GND 0.00fF
C1080 IN_N.n59 GND 0.04fF
C1081 IN_N.n60 GND 0.15fF
C1082 IN_N.n61 GND 0.04fF
C1083 IN_N.n62 GND 0.02fF
C1084 IN_N.n63 GND 0.04fF
C1085 IN_N.n64 GND 0.01fF
C1086 IN_N.n65 GND 0.01fF
C1087 IN_N.n66 GND 0.09fF
C1088 IN_N.n67 GND 0.01fF
C1089 IN_N.n68 GND 0.01fF
C1090 IN_N.n69 GND 0.02fF
C1091 IN_N.n70 GND 0.03fF
C1092 IN_N.n71 GND 0.02fF
C1093 IN_N.n72 GND 0.01fF
C1094 IN_N.n73 GND 0.03fF
C1095 IN_N.n74 GND 0.02fF
C1096 IN_N.n75 GND 0.02fF
C1097 IN_N.n76 GND 0.00fF
C1098 IN_N.n77 GND 0.01fF
C1099 IN_N.n78 GND 0.01fF
C1100 IN_N.n79 GND 0.01fF
C1101 IN_N.n80 GND 0.02fF
C1102 IN_N.n81 GND 0.01fF
C1103 IN_N.n82 GND 0.17fF
C1104 IN_N.n83 GND 0.02fF
C1105 IN_N.n84 GND 0.01fF
C1106 IN_N.n85 GND 0.03fF
C1107 IN_N.n86 GND 0.00fF
C1108 IN_N.n87 GND 0.01fF
C1109 IN_N.n88 GND 0.01fF
C1110 IN_N.n89 GND 0.02fF
C1111 IN_N.n90 GND 0.01fF
C1112 IN_N.n91 GND 0.01fF
C1113 IN_N.n92 GND 0.01fF
C1114 IN_N.n93 GND 0.05fF
C1115 IN_N.n94 GND 0.03fF
C1116 IN_N.n95 GND 0.01fF
C1117 IN_N.n96 GND 0.01fF
C1118 IN_N.n97 GND 0.01fF
C1119 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE GND 0.03fF
C1120 IN_N.n98 GND 0.00fF
C1121 IN_N.n99 GND 0.01fF
C1122 IN_N.n100 GND 0.02fF
C1123 IN_N.n101 GND 0.02fF
C1124 IN_N.n102 GND 0.01fF
C1125 IN_N.n103 GND 0.02fF
C1126 IN_N.n104 GND 0.01fF
C1127 IN_N.n105 GND 0.17fF
C1128 IN_N.n106 GND 0.02fF
C1129 IN_N.n107 GND 0.01fF
C1130 IN_N.n108 GND 0.03fF
C1131 IN_N.n109 GND 0.01fF
C1132 IN_N.n110 GND 0.01fF
C1133 IN_N.n111 GND 0.01fF
C1134 IN_N.n112 GND 0.02fF
C1135 IN_N.n113 GND 0.01fF
C1136 IN_N.n114 GND 0.01fF
C1137 IN_N.n115 GND 0.01fF
C1138 IN_N.n116 GND 0.01fF
C1139 IN_N.n117 GND 0.01fF
C1140 IN_N.n118 GND 0.02fF
C1141 IN_N.n119 GND 0.02fF
C1142 IN_N.n120 GND 0.02fF
C1143 IN_N.n121 GND 0.02fF
C1144 IN_N.n122 GND 0.01fF
C1145 IN_N.n123 GND 0.02fF
C1146 IN_N.n124 GND 0.01fF
C1147 IN_N.n125 GND 0.01fF
C1148 IN_N.n126 GND 0.02fF
C1149 IN_N.n127 GND 0.01fF
C1150 IN_N.n128 GND 0.01fF
C1151 IN_N.n129 GND 0.02fF
C1152 IN_N.n130 GND 0.01fF
C1153 IN_N.n131 GND 0.02fF
C1154 IN_N.n132 GND 0.02fF
C1155 IN_N.n133 GND 0.09fF
C1156 IN_N.n134 GND 0.32fF
C1157 IN_N.n135 GND 0.10fF
C1158 IN_N.n136 GND 0.04fF
C1159 IN_N.n137 GND 0.04fF
C1160 IN_N.n138 GND 0.09fF
C1161 IN_N.n139 GND 0.09fF
C1162 IN_N.n140 GND 0.04fF
C1163 IN_N.n141 GND 0.04fF
C1164 IN_N.n142 GND 0.10fF
C1165 IN_N.n143 GND 0.12fF
C1166 IN_N.n144 GND 0.05fF
C1167 IN_N.n145 GND 2.48fF
C1168 IN_N.n146 GND 1.82fF
C1169 IN_N.n147 GND 0.04fF
C1170 IN_N.n148 GND 0.17fF
C1171 IN_N.n149 GND 0.02fF
C1172 IN_N.n150 GND 0.03fF
C1173 IN_N.n151 GND 0.06fF
C1174 IN_N.n152 GND 0.02fF
C1175 IN_N.n153 GND 0.01fF
C1176 IN_N.n154 GND 0.01fF
C1177 IN_N.n155 GND 0.00fF
C1178 IN_N.n156 GND 0.00fF
C1179 IN_N.n157 GND 0.04fF
C1180 IN_N.n158 GND 0.15fF
C1181 IN_N.n159 GND 0.04fF
C1182 IN_N.n160 GND 0.02fF
C1183 IN_N.n161 GND 0.04fF
C1184 IN_N.n162 GND 0.01fF
C1185 IN_N.n163 GND 0.01fF
C1186 IN_N.n164 GND 0.09fF
C1187 IN_N.n165 GND 0.01fF
C1188 IN_N.n166 GND 0.01fF
C1189 IN_N.n167 GND 0.02fF
C1190 IN_N.n168 GND 0.03fF
C1191 IN_N.n169 GND 0.02fF
C1192 IN_N.n170 GND 0.01fF
C1193 IN_N.n171 GND 0.03fF
C1194 IN_N.n172 GND 0.02fF
C1195 IN_N.n173 GND 0.02fF
C1196 IN_N.n174 GND 0.00fF
C1197 IN_N.n175 GND 0.01fF
C1198 IN_N.n176 GND 0.01fF
C1199 IN_N.n177 GND 0.01fF
C1200 IN_N.n178 GND 0.02fF
C1201 IN_N.n179 GND 0.01fF
C1202 IN_N.n180 GND 0.17fF
C1203 IN_N.n181 GND 0.02fF
C1204 IN_N.n182 GND 0.01fF
C1205 IN_N.n183 GND 0.03fF
C1206 IN_N.n184 GND 0.00fF
C1207 IN_N.n185 GND 0.01fF
C1208 IN_N.n186 GND 0.01fF
C1209 IN_N.n187 GND 0.02fF
C1210 IN_N.n188 GND 0.01fF
C1211 IN_N.n189 GND 0.01fF
C1212 IN_N.n190 GND 0.01fF
C1213 IN_N.n191 GND 0.05fF
C1214 IN_N.n192 GND 0.03fF
C1215 IN_N.n193 GND 0.01fF
C1216 IN_N.n194 GND 0.01fF
C1217 IN_N.n195 GND 0.01fF
C1218 IN_N.n196 GND 0.00fF
C1219 IN_N.n197 GND 0.01fF
C1220 IN_N.n198 GND 0.02fF
C1221 IN_N.n199 GND 0.02fF
C1222 IN_N.n200 GND 0.01fF
C1223 IN_N.n201 GND 0.02fF
C1224 IN_N.n202 GND 0.01fF
C1225 IN_N.n203 GND 0.17fF
C1226 IN_N.n204 GND 0.02fF
C1227 IN_N.n205 GND 0.01fF
C1228 IN_N.n206 GND 0.03fF
C1229 IN_N.n207 GND 0.01fF
C1230 IN_N.n208 GND 0.01fF
C1231 IN_N.n209 GND 0.01fF
C1232 IN_N.n210 GND 0.02fF
C1233 IN_N.n211 GND 0.01fF
C1234 IN_N.n212 GND 0.01fF
C1235 IN_N.n213 GND 0.01fF
C1236 IN_N.n214 GND 0.01fF
C1237 IN_N.n215 GND 0.01fF
C1238 IN_N.n216 GND 0.02fF
C1239 IN_N.n217 GND 0.02fF
C1240 IN_N.n218 GND 0.02fF
C1241 IN_N.n219 GND 0.02fF
C1242 IN_N.n220 GND 0.01fF
C1243 IN_N.n221 GND 0.02fF
C1244 IN_N.n222 GND 0.01fF
C1245 IN_N.n223 GND 0.01fF
C1246 IN_N.n224 GND 0.02fF
C1247 IN_N.n225 GND 0.01fF
C1248 IN_N.n226 GND 0.01fF
C1249 IN_N.n227 GND 0.02fF
C1250 IN_N.n228 GND 0.01fF
C1251 IN_N.n229 GND 0.02fF
C1252 IN_N.n230 GND 0.02fF
C1253 IN_N.n231 GND 0.09fF
C1254 IN_N.n232 GND 0.11fF
C1255 IN_N.n233 GND 0.03fF
C1256 IN_N.n234 GND 0.01fF
C1257 IN_N.n235 GND 0.01fF
C1258 IN_N.n236 GND 0.03fF
C1259 IN_N.n237 GND 0.03fF
C1260 IN_N.n238 GND 0.01fF
C1261 IN_N.n239 GND 0.01fF
C1262 IN_N.n240 GND 0.03fF
C1263 IN_N.n241 GND 0.04fF
C1264 IN_N.n242 GND 0.02fF
C1265 IN_N.n243 GND 1.39fF
C1266 IN_N.n244 GND 1.47fF
C1267 IN_N.n245 GND 0.25fF
C1268 IN_N.n246 GND 0.02fF
C1269 IN_N.n247 GND 0.01fF
C1270 IN_N.n248 GND 0.04fF
C1271 IN_N.n249 GND 0.05fF
C1272 IN_N.n250 GND 0.03fF
C1273 IN_N.n251 GND 0.02fF
C1274 IN_N.n252 GND 0.01fF
C1275 IN_N.n253 GND 0.01fF
C1276 IN_N.n254 GND 0.01fF
C1277 IN_N.n255 GND 0.00fF
C1278 IN_N.n256 GND 0.02fF
C1279 IN_N.n257 GND 0.01fF
C1280 IN_N.t3 GND 0.27fF $ **FLOATING
C1281 IN_N.n258 GND 0.17fF
C1282 IN_N.n259 GND 0.02fF
C1283 IN_N.n260 GND 0.01fF
C1284 IN_N.n261 GND 0.03fF
C1285 IN_N.n262 GND 0.00fF
C1286 IN_N.n263 GND 0.01fF
C1287 IN_N.n264 GND 0.01fF
C1288 IN_N.n265 GND 0.01fF
C1289 IN_N.n266 GND 0.02fF
C1290 IN_N.n267 GND 0.01fF
C1291 IN_N.n268 GND 0.00fF
C1292 IN_N.n269 GND 0.05fF
C1293 IN_N.n270 GND 0.03fF
C1294 IN_N.n271 GND 0.01fF
C1295 IN_N.n272 GND 0.03fF
C1296 IN_N.n273 GND 0.02fF
C1297 IN_N.n274 GND 0.01fF
C1298 IN_N.n275 GND 0.02fF
C1299 IN_N.n276 GND 0.01fF
C1300 IN_N.t6 GND 0.27fF $ **FLOATING
C1301 IN_N.n277 GND 0.17fF
C1302 IN_N.n278 GND 0.02fF
C1303 IN_N.n279 GND 0.01fF
C1304 IN_N.n280 GND 0.03fF
C1305 IN_N.n281 GND 0.00fF
C1306 IN_N.n282 GND 0.01fF
C1307 IN_N.n283 GND 0.01fF
C1308 IN_N.n284 GND 0.01fF
C1309 IN_N.n285 GND 0.01fF
C1310 IN_N.n286 GND 0.02fF
C1311 IN_N.n287 GND 0.00fF
C1312 IN_N.n288 GND 0.02fF
C1313 IN_N.n289 GND 0.03fF
C1314 IN_N.n290 GND 0.02fF
C1315 IN_N.t0 GND 0.27fF $ **FLOATING
C1316 IN_N.n291 GND 0.04fF
C1317 IN_N.n292 GND 0.17fF
C1318 IN_N.n293 GND 0.03fF
C1319 IN_N.n294 GND 0.05fF
C1320 IN_N.n295 GND 0.04fF
C1321 IN_N.n296 GND 0.01fF
C1322 IN_N.n297 GND 0.02fF
C1323 IN_N.n298 GND 0.02fF
C1324 IN_N.n299 GND 0.01fF
C1325 IN_N.n300 GND 0.01fF
C1326 IN_N.n301 GND 0.02fF
C1327 IN_N.n302 GND 1.24fF
C1328 IN_N.n303 GND 0.98fF
C1329 IN_N.n304 GND 0.02fF
C1330 IN_N.n305 GND 0.04fF
C1331 IN_N.n306 GND 0.04fF
C1332 IN_N.n307 GND 0.01fF
C1333 IN_N.n308 GND 0.01fF
C1334 IN_N.n309 GND 0.03fF
C1335 IN_N.n310 GND 0.03fF
C1336 IN_N.n311 GND 0.01fF
C1337 IN_N.n312 GND 0.01fF
C1338 IN_N.n313 GND 0.04fF
C1339 IN_N.n315 GND 0.04fF
C1340 IN_N.n316 GND 0.05fF
C1341 IN_N.n317 GND 0.03fF
C1342 IN_N.n318 GND 0.02fF
C1343 IN_N.n319 GND 0.02fF
C1344 IN_N.n320 GND 0.00fF
C1345 IN_N.n321 GND 0.01fF
C1346 IN_N.n322 GND 0.01fF
C1347 IN_N.n323 GND 0.01fF
C1348 IN_N.n324 GND 0.02fF
C1349 IN_N.n325 GND 0.01fF
C1350 IN_N.t7 GND 0.27fF $ **FLOATING
C1351 IN_N.n326 GND 0.17fF
C1352 IN_N.n327 GND 0.02fF
C1353 IN_N.n328 GND 0.01fF
C1354 IN_N.n329 GND 0.03fF
C1355 IN_N.n330 GND 0.00fF
C1356 IN_N.n331 GND 0.01fF
C1357 IN_N.n332 GND 0.01fF
C1358 IN_N.n333 GND 0.02fF
C1359 IN_N.n334 GND 0.03fF
C1360 IN_N.n335 GND 0.05fF
C1361 IN_N.n336 GND 0.03fF
C1362 IN_N.n337 GND 0.01fF
C1363 IN_N.n338 GND 0.00fF
C1364 IN_N.n339 GND 0.01fF
C1365 IN_N.n340 GND 0.02fF
C1366 IN_N.n341 GND 0.02fF
C1367 IN_N.n342 GND 0.01fF
C1368 IN_N.n343 GND 0.02fF
C1369 IN_N.n344 GND 0.01fF
C1370 IN_N.n345 GND 0.00fF
C1371 IN_N.n346 GND 0.01fF
C1372 IN_N.n347 GND 0.02fF
C1373 IN_N.n348 GND 0.01fF
C1374 IN_N.n349 GND 0.01fF
C1375 IN_N.n350 GND 0.01fF
C1376 IN_N.n351 GND 0.01fF
C1377 IN_N.n352 GND 0.01fF
C1378 IN_N.n353 GND 0.01fF
C1379 IN_N.n354 GND 0.01fF
C1380 IN_N.n355 GND 0.01fF
C1381 IN_N.n356 GND 0.02fF
C1382 IN_N.n357 GND 0.01fF
C1383 IN_N.n358 GND 0.01fF
C1384 IN_N.n359 GND 0.04fF
C1385 IN_N.n360 GND 0.02fF
C1386 IN_N.t1 GND 0.27fF $ **FLOATING
C1387 IN_N.n361 GND 0.04fF
C1388 IN_N.n362 GND 0.17fF
C1389 IN_N.n363 GND 0.03fF
C1390 IN_N.n364 GND 0.05fF
C1391 IN_N.n365 GND 0.03fF
C1392 IN_N.n366 GND 0.02fF
C1393 IN_N.n367 GND 0.01fF
C1394 IN_N.n368 GND 0.01fF
C1395 IN_N.n369 GND 0.01fF
C1396 IN_N.n370 GND 0.00fF
C1397 IN_N.n371 GND 0.02fF
C1398 IN_N.n372 GND 0.01fF
C1399 IN_N.t5 GND 0.27fF $ **FLOATING
C1400 IN_N.n373 GND 0.17fF
C1401 IN_N.n374 GND 0.02fF
C1402 IN_N.n375 GND 0.01fF
C1403 IN_N.n376 GND 0.03fF
C1404 IN_N.n377 GND 0.00fF
C1405 IN_N.n378 GND 0.01fF
C1406 IN_N.n379 GND 0.01fF
C1407 IN_N.n380 GND 0.01fF
C1408 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n0 GND 0.37fF
C1409 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1 GND 7.36fF
C1410 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n2 GND 0.24fF
C1411 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n3 GND 0.24fF
C1412 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n4 GND 0.55fF
C1413 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n5 GND 0.55fF
C1414 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n6 GND 0.55fF
C1415 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n7 GND 0.55fF
C1416 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n8 GND 0.55fF
C1417 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n9 GND 0.55fF
C1418 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n10 GND 0.55fF
C1419 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n11 GND 0.00fF
C1420 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n12 GND 0.04fF
C1421 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n13 GND 0.01fF
C1422 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n14 GND 0.00fF
C1423 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n15 GND 0.00fF
C1424 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n16 GND 0.04fF
C1425 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n17 GND 0.01fF
C1426 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n18 GND 0.00fF
C1427 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n19 GND 0.00fF
C1428 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n20 GND 0.04fF
C1429 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n21 GND 0.01fF
C1430 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n22 GND 0.00fF
C1431 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n23 GND 0.00fF
C1432 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n24 GND 0.04fF
C1433 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n25 GND 0.01fF
C1434 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n26 GND 0.00fF
C1435 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n27 GND 0.00fF
C1436 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n28 GND 0.04fF
C1437 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n29 GND 0.01fF
C1438 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n30 GND 0.00fF
C1439 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n31 GND 0.00fF
C1440 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n32 GND 0.04fF
C1441 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n33 GND 0.01fF
C1442 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n34 GND 0.00fF
C1443 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n35 GND 0.00fF
C1444 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n36 GND 0.04fF
C1445 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n37 GND 0.01fF
C1446 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n38 GND 0.00fF
C1447 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n39 GND 0.01fF
C1448 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n40 GND 0.00fF
C1449 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n41 GND 0.01fF
C1450 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n42 GND 0.00fF
C1451 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n43 GND 0.01fF
C1452 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n44 GND 0.01fF
C1453 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n45 GND 0.01fF
C1454 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n46 GND 0.01fF
C1455 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n47 GND 0.01fF
C1456 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n48 GND 0.01fF
C1457 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n49 GND 0.01fF
C1458 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n50 GND 0.01fF
C1459 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n51 GND 0.01fF
C1460 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n52 GND 0.01fF
C1461 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n53 GND 0.01fF
C1462 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n54 GND 0.01fF
C1463 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n55 GND 0.01fF
C1464 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n56 GND 0.01fF
C1465 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n57 GND 0.01fF
C1466 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n58 GND 0.01fF
C1467 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n59 GND 0.01fF
C1468 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n60 GND 0.01fF
C1469 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n61 GND 0.01fF
C1470 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n62 GND 0.01fF
C1471 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n63 GND 0.01fF
C1472 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n64 GND 0.01fF
C1473 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n65 GND 0.01fF
C1474 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n66 GND 0.01fF
C1475 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n67 GND 0.01fF
C1476 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n68 GND 0.01fF
C1477 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n69 GND 0.01fF
C1478 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n70 GND 0.01fF
C1479 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n71 GND 0.01fF
C1480 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n72 GND 0.01fF
C1481 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n73 GND 0.01fF
C1482 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n74 GND 0.01fF
C1483 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n75 GND 0.01fF
C1484 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n76 GND 0.01fF
C1485 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n77 GND 0.01fF
C1486 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n78 GND 0.01fF
C1487 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n79 GND 0.01fF
C1488 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n80 GND 0.01fF
C1489 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n81 GND 0.01fF
C1490 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n82 GND 0.01fF
C1491 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n83 GND 0.01fF
C1492 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n84 GND 0.01fF
C1493 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n85 GND 0.01fF
C1494 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n86 GND 0.01fF
C1495 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n87 GND 0.01fF
C1496 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n88 GND 0.01fF
C1497 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n89 GND 0.01fF
C1498 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n90 GND 0.01fF
C1499 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n91 GND 0.01fF
C1500 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n92 GND 0.01fF
C1501 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n93 GND 0.01fF
C1502 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n94 GND 0.01fF
C1503 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n95 GND 0.01fF
C1504 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n96 GND 0.01fF
C1505 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n97 GND 0.01fF
C1506 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n98 GND 0.01fF
C1507 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n99 GND 0.01fF
C1508 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n100 GND 0.01fF
C1509 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n101 GND 0.01fF
C1510 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n102 GND 0.01fF
C1511 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n103 GND 0.01fF
C1512 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n104 GND 0.01fF
C1513 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n105 GND 0.01fF
C1514 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n106 GND 0.00fF
C1515 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n107 GND 0.00fF
C1516 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n108 GND 0.00fF
C1517 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n109 GND 0.01fF
C1518 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n110 GND 0.00fF
C1519 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n111 GND 0.01fF
C1520 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n112 GND 0.00fF
C1521 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n113 GND 0.01fF
C1522 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n114 GND 0.00fF
C1523 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n115 GND 0.01fF
C1524 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n116 GND 0.00fF
C1525 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n117 GND 0.01fF
C1526 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n118 GND 0.00fF
C1527 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n119 GND 0.00fF
C1528 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n120 GND 0.00fF
C1529 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n121 GND 0.00fF
C1530 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n122 GND 0.00fF
C1531 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n123 GND 0.00fF
C1532 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n124 GND 0.00fF
C1533 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n125 GND 0.61fF
C1534 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n126 GND 0.72fF
C1535 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n127 GND 2.09fF
C1536 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n128 GND 0.72fF
C1537 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n129 GND 0.61fF
C1538 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n130 GND 2.09fF
C1539 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n131 GND 1.00fF
C1540 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n132 GND 3.75fF
C1541 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n133 GND 1.00fF
C1542 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n134 GND 4.36fF
C1543 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n135 GND 1.00fF
C1544 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n136 GND 4.36fF
C1545 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n137 GND 1.00fF
C1546 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n138 GND 0.87fF
C1547 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n139 GND 2.44fF
C1548 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n140 GND 1.00fF
C1549 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n141 GND 4.36fF
C1550 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n142 GND 1.00fF
C1551 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n143 GND 4.36fF
C1552 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n144 GND 1.00fF
C1553 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n145 GND 0.87fF
C1554 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n146 GND 2.44fF
C1555 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n147 GND 0.01fF
C1556 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n148 GND 0.00fF
C1557 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n149 GND 0.00fF
C1558 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n150 GND 0.01fF
C1559 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n151 GND 0.01fF
C1560 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n152 GND 0.00fF
C1561 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n153 GND 0.00fF
C1562 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n154 GND 0.00fF
C1563 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n155 GND 0.00fF
C1564 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n156 GND 0.00fF
C1565 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n157 GND 0.00fF
C1566 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n158 GND 0.01fF
C1567 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n159 GND 0.01fF
C1568 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n160 GND 0.01fF
C1569 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n161 GND 0.01fF
C1570 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n162 GND 0.01fF
C1571 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n163 GND 0.00fF
C1572 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n164 GND 0.00fF
C1573 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n165 GND 0.00fF
C1574 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n166 GND 0.00fF
C1575 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n167 GND 0.00fF
C1576 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n168 GND 0.01fF
C1577 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n169 GND 0.01fF
C1578 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n170 GND 0.01fF
C1579 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n171 GND 0.01fF
C1580 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n172 GND 0.01fF
C1581 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n173 GND 0.00fF
C1582 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n174 GND 0.00fF
C1583 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n175 GND 0.00fF
C1584 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n176 GND 0.00fF
C1585 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n177 GND 0.01fF
C1586 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t10 GND 0.13fF $
+ **FLOATING
C1587 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t6 GND 0.13fF $
+ **FLOATING
C1588 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n178 GND 0.37fF
C1589 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n179 GND 0.04fF
C1590 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n180 GND 0.29fF
C1591 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n181 GND 0.01fF
C1592 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n182 GND 0.01fF
C1593 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n183 GND 0.00fF
C1594 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n184 GND 0.00fF
C1595 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n185 GND 0.00fF
C1596 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n186 GND 0.00fF
C1597 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n187 GND 0.00fF
C1598 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n188 GND 0.00fF
C1599 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n189 GND 0.01fF
C1600 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n190 GND 0.00fF
C1601 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n191 GND 0.00fF
C1602 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n192 GND 0.00fF
C1603 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n193 GND 0.01fF
C1604 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n194 GND 0.01fF
C1605 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n195 GND 0.01fF
C1606 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n196 GND 0.01fF
C1607 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n197 GND 0.01fF
C1608 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n198 GND 0.00fF
C1609 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n199 GND 0.01fF
C1610 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n200 GND 0.00fF
C1611 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n201 GND 0.01fF
C1612 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n202 GND 0.00fF
C1613 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n203 GND 0.01fF
C1614 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n204 GND 0.00fF
C1615 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n205 GND 0.97fF
C1616 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n206 GND 0.00fF
C1617 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n207 GND 0.00fF
C1618 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n208 GND 0.00fF
C1619 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n209 GND 0.00fF
C1620 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n210 GND 0.00fF
C1621 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n211 GND 0.00fF
C1622 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n212 GND 0.00fF
C1623 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n213 GND 0.00fF
C1624 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n214 GND 0.00fF
C1625 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n215 GND 0.42fF
C1626 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n216 GND 0.42fF
C1627 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n217 GND 0.42fF
C1628 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n218 GND 0.42fF
C1629 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n219 GND 0.42fF
C1630 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n220 GND 0.42fF
C1631 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n221 GND 0.42fF
C1632 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n222 GND 1.22fF
C1633 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n223 GND 0.01fF
C1634 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n224 GND 0.00fF
C1635 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n225 GND 0.00fF
C1636 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n226 GND 0.00fF
C1637 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n227 GND 0.01fF
C1638 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n228 GND 0.01fF
C1639 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n229 GND 0.01fF
C1640 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n230 GND 0.01fF
C1641 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n231 GND 0.01fF
C1642 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n232 GND 0.00fF
C1643 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n233 GND 0.01fF
C1644 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n234 GND 0.00fF
C1645 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n235 GND 0.01fF
C1646 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n236 GND 0.00fF
C1647 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n237 GND 0.01fF
C1648 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n238 GND 0.00fF
C1649 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n239 GND 0.01fF
C1650 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n240 GND 0.01fF
C1651 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n241 GND 0.00fF
C1652 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n242 GND 0.00fF
C1653 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n243 GND 0.00fF
C1654 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n244 GND 0.00fF
C1655 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n245 GND 0.00fF
C1656 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n246 GND 0.00fF
C1657 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n247 GND 0.01fF
C1658 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n248 GND 0.01fF
C1659 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n249 GND 0.01fF
C1660 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n250 GND 0.01fF
C1661 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n251 GND 0.01fF
C1662 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n252 GND 0.00fF
C1663 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n253 GND 0.00fF
C1664 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n254 GND 0.00fF
C1665 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n255 GND 0.00fF
C1666 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n256 GND 0.00fF
C1667 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n257 GND 0.00fF
C1668 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n258 GND 0.01fF
C1669 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n259 GND 0.01fF
C1670 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n260 GND 0.01fF
C1671 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n261 GND 0.01fF
C1672 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n262 GND 0.01fF
C1673 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n263 GND 0.00fF
C1674 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n264 GND 0.00fF
C1675 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n265 GND 0.00fF
C1676 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n266 GND 0.00fF
C1677 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n267 GND 0.01fF
C1678 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t2 GND 0.13fF $
+ **FLOATING
C1679 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n268 GND 0.49fF
C1680 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n269 GND 0.05fF
C1681 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n270 GND 0.28fF
C1682 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n271 GND 0.01fF
C1683 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n272 GND 0.01fF
C1684 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n273 GND 0.00fF
C1685 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n274 GND 0.00fF
C1686 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n275 GND 0.00fF
C1687 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n276 GND 0.00fF
C1688 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n277 GND 0.00fF
C1689 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n278 GND 0.00fF
C1690 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n279 GND 0.01fF
C1691 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n280 GND 0.14fF
C1692 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n281 GND 0.01fF
C1693 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n282 GND 0.00fF
C1694 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n283 GND 0.01fF
C1695 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n284 GND 0.00fF
C1696 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n285 GND 0.00fF
C1697 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n286 GND 0.01fF
C1698 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n287 GND 0.01fF
C1699 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n288 GND 0.01fF
C1700 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n289 GND 0.01fF
C1701 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n290 GND 0.01fF
C1702 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n291 GND 0.00fF
C1703 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n292 GND 0.00fF
C1704 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n293 GND 0.00fF
C1705 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n294 GND 0.00fF
C1706 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n295 GND 0.01fF
C1707 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n296 GND 0.01fF
C1708 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n297 GND 0.01fF
C1709 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n298 GND 0.00fF
C1710 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n299 GND 0.01fF
C1711 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n300 GND 0.00fF
C1712 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n301 GND 0.00fF
C1713 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n302 GND 0.00fF
C1714 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n303 GND 0.00fF
C1715 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n304 GND 0.01fF
C1716 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n305 GND 0.00fF
C1717 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n306 GND 0.01fF
C1718 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n307 GND 0.01fF
C1719 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n308 GND 0.00fF
C1720 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n309 GND 0.01fF
C1721 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n310 GND 0.00fF
C1722 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n311 GND 0.01fF
C1723 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n312 GND 0.00fF
C1724 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n313 GND 0.00fF
C1725 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n314 GND 0.00fF
C1726 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n315 GND 0.00fF
C1727 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n316 GND 0.01fF
C1728 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n317 GND 0.00fF
C1729 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n318 GND 0.01fF
C1730 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n319 GND 0.01fF
C1731 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n320 GND 0.01fF
C1732 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n321 GND 0.00fF
C1733 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n322 GND 0.00fF
C1734 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n323 GND 0.01fF
C1735 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n324 GND 0.01fF
C1736 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n325 GND 0.00fF
C1737 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n326 GND 0.00fF
C1738 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n327 GND 0.00fF
C1739 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n328 GND 0.00fF
C1740 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n329 GND 0.00fF
C1741 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n330 GND 0.01fF
C1742 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t38 GND 0.13fF $
+ **FLOATING
C1743 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t23 GND 0.13fF $
+ **FLOATING
C1744 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n331 GND 0.37fF
C1745 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n332 GND 0.05fF
C1746 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n333 GND 0.28fF
C1747 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n334 GND 0.01fF
C1748 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n335 GND 0.00fF
C1749 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n336 GND 0.00fF
C1750 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n337 GND 0.00fF
C1751 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n338 GND 0.01fF
C1752 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n339 GND 0.01fF
C1753 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n340 GND 0.01fF
C1754 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n341 GND 0.01fF
C1755 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n342 GND 0.00fF
C1756 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n343 GND 0.00fF
C1757 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n344 GND 0.00fF
C1758 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n345 GND 0.00fF
C1759 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n346 GND 0.01fF
C1760 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n347 GND 0.01fF
C1761 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n348 GND 0.01fF
C1762 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n349 GND 0.01fF
C1763 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n350 GND 0.01fF
C1764 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n351 GND 0.00fF
C1765 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n352 GND 0.00fF
C1766 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n353 GND 0.00fF
C1767 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n354 GND 0.00fF
C1768 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n355 GND 0.01fF
C1769 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n356 GND 0.01fF
C1770 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n357 GND 0.01fF
C1771 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n358 GND 0.01fF
C1772 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n359 GND 0.01fF
C1773 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n360 GND 0.00fF
C1774 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n361 GND 0.00fF
C1775 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n362 GND 0.01fF
C1776 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n363 GND 0.00fF
C1777 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n364 GND 0.01fF
C1778 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n365 GND 0.00fF
C1779 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n366 GND 0.01fF
C1780 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n367 GND 0.17fF
C1781 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n368 GND 1.44fF
C1782 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n369 GND 0.53fF
C1783 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN GND 0.45fF
C1784 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n370 GND 0.00fF
C1785 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n371 GND 0.00fF
C1786 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n372 GND 0.00fF
C1787 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n373 GND 0.01fF
C1788 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t27 GND 0.13fF $
+ **FLOATING
C1789 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t44 GND 0.13fF $
+ **FLOATING
C1790 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n374 GND 0.37fF
C1791 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n375 GND 0.05fF
C1792 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n376 GND 0.28fF
C1793 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n377 GND 0.01fF
C1794 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n378 GND 0.00fF
C1795 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n379 GND 0.00fF
C1796 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n380 GND 0.00fF
C1797 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n381 GND 0.01fF
C1798 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n382 GND 0.01fF
C1799 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n383 GND 0.00fF
C1800 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n384 GND 0.00fF
C1801 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n385 GND 0.00fF
C1802 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n386 GND 0.01fF
C1803 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n387 GND 0.01fF
C1804 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n388 GND 0.01fF
C1805 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n389 GND 0.01fF
C1806 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n390 GND 0.01fF
C1807 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n391 GND 0.00fF
C1808 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n392 GND 0.00fF
C1809 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n393 GND 0.00fF
C1810 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n394 GND 0.00fF
C1811 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n395 GND 0.01fF
C1812 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n396 GND 0.01fF
C1813 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n397 GND 0.01fF
C1814 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n398 GND 0.00fF
C1815 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n399 GND 0.01fF
C1816 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n400 GND 0.01fF
C1817 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n401 GND 0.00fF
C1818 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n402 GND 0.00fF
C1819 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n403 GND 0.00fF
C1820 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n404 GND 0.00fF
C1821 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n405 GND 0.04fF
C1822 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n406 GND 0.01fF
C1823 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n407 GND 0.01fF
C1824 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n408 GND 0.01fF
C1825 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n409 GND 0.00fF
C1826 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n410 GND 0.00fF
C1827 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n411 GND 0.00fF
C1828 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n412 GND 0.00fF
C1829 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n413 GND 0.01fF
C1830 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n414 GND 0.01fF
C1831 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n415 GND 0.01fF
C1832 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n416 GND 0.00fF
C1833 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n417 GND 0.01fF
C1834 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n418 GND 0.00fF
C1835 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n419 GND 0.00fF
C1836 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n420 GND 0.01fF
C1837 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n421 GND 0.01fF
C1838 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n422 GND 0.01fF
C1839 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n423 GND 0.01fF
C1840 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n424 GND 0.00fF
C1841 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n425 GND 0.00fF
C1842 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n426 GND 0.00fF
C1843 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n427 GND 0.01fF
C1844 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t45 GND 0.13fF $
+ **FLOATING
C1845 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t20 GND 0.13fF $
+ **FLOATING
C1846 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n428 GND 0.37fF
C1847 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n429 GND 0.05fF
C1848 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n430 GND 0.28fF
C1849 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n431 GND 0.01fF
C1850 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n432 GND 0.00fF
C1851 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n433 GND 0.00fF
C1852 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n434 GND 0.00fF
C1853 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n435 GND 0.01fF
C1854 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n436 GND 0.01fF
C1855 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n437 GND 0.00fF
C1856 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n438 GND 0.00fF
C1857 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n439 GND 0.00fF
C1858 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n440 GND 0.00fF
C1859 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n441 GND 0.01fF
C1860 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n442 GND 0.01fF
C1861 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n443 GND 0.01fF
C1862 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n444 GND 0.01fF
C1863 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n445 GND 0.01fF
C1864 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n446 GND 0.00fF
C1865 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n447 GND 0.00fF
C1866 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n448 GND 0.00fF
C1867 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n449 GND 0.00fF
C1868 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n450 GND 0.01fF
C1869 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n451 GND 0.01fF
C1870 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n452 GND 0.01fF
C1871 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n453 GND 0.00fF
C1872 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n454 GND 0.00fF
C1873 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n455 GND 0.01fF
C1874 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n456 GND 0.01fF
C1875 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n457 GND 0.01fF
C1876 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n458 GND 0.01fF
C1877 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n459 GND 0.00fF
C1878 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n460 GND 0.00fF
C1879 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n461 GND 0.01fF
C1880 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n462 GND 0.00fF
C1881 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n463 GND 0.01fF
C1882 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n464 GND 0.00fF
C1883 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n465 GND 0.01fF
C1884 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n466 GND 0.01fF
C1885 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n467 GND 0.00fF
C1886 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n468 GND 0.01fF
C1887 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n469 GND 0.00fF
C1888 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n470 GND 0.00fF
C1889 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n471 GND 0.00fF
C1890 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n472 GND 0.00fF
C1891 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n473 GND 0.53fF
C1892 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/DRAIN GND 0.45fF
C1893 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n474 GND 0.00fF
C1894 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n475 GND 0.00fF
C1895 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n476 GND 0.00fF
C1896 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n477 GND 0.01fF
C1897 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t36 GND 0.13fF $
+ **FLOATING
C1898 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t37 GND 0.13fF $
+ **FLOATING
C1899 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n478 GND 0.37fF
C1900 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n479 GND 0.05fF
C1901 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n480 GND 0.28fF
C1902 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n481 GND 0.01fF
C1903 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n482 GND 0.00fF
C1904 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n483 GND 0.00fF
C1905 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n484 GND 0.00fF
C1906 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n485 GND 0.01fF
C1907 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n486 GND 0.01fF
C1908 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n487 GND 0.00fF
C1909 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n488 GND 0.00fF
C1910 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n489 GND 0.00fF
C1911 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n490 GND 0.01fF
C1912 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n491 GND 0.01fF
C1913 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n492 GND 0.01fF
C1914 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n493 GND 0.01fF
C1915 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n494 GND 0.01fF
C1916 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n495 GND 0.00fF
C1917 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n496 GND 0.00fF
C1918 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n497 GND 0.00fF
C1919 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n498 GND 0.00fF
C1920 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n499 GND 0.01fF
C1921 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n500 GND 0.01fF
C1922 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n501 GND 0.01fF
C1923 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n502 GND 0.00fF
C1924 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n503 GND 0.01fF
C1925 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n504 GND 0.01fF
C1926 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n505 GND 0.00fF
C1927 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n506 GND 0.00fF
C1928 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n507 GND 0.00fF
C1929 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n508 GND 0.00fF
C1930 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n509 GND 0.04fF
C1931 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n510 GND 0.01fF
C1932 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n511 GND 0.01fF
C1933 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n512 GND 0.01fF
C1934 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n513 GND 0.00fF
C1935 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n514 GND 0.00fF
C1936 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n515 GND 0.00fF
C1937 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n516 GND 0.00fF
C1938 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n517 GND 0.01fF
C1939 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n518 GND 0.01fF
C1940 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n519 GND 0.01fF
C1941 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n520 GND 0.00fF
C1942 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n521 GND 0.01fF
C1943 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n522 GND 0.00fF
C1944 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n523 GND 0.00fF
C1945 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n524 GND 0.01fF
C1946 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n525 GND 0.01fF
C1947 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n526 GND 0.01fF
C1948 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n527 GND 0.01fF
C1949 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n528 GND 0.00fF
C1950 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n529 GND 0.00fF
C1951 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n530 GND 0.00fF
C1952 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n531 GND 0.01fF
C1953 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t40 GND 0.13fF $
+ **FLOATING
C1954 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t25 GND 0.13fF $
+ **FLOATING
C1955 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n532 GND 0.37fF
C1956 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n533 GND 0.05fF
C1957 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n534 GND 0.28fF
C1958 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n535 GND 0.01fF
C1959 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n536 GND 0.00fF
C1960 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n537 GND 0.00fF
C1961 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n538 GND 0.00fF
C1962 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n539 GND 0.01fF
C1963 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n540 GND 0.01fF
C1964 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n541 GND 0.00fF
C1965 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n542 GND 0.00fF
C1966 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n543 GND 0.00fF
C1967 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n544 GND 0.00fF
C1968 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n545 GND 0.01fF
C1969 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n546 GND 0.01fF
C1970 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n547 GND 0.01fF
C1971 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n548 GND 0.01fF
C1972 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n549 GND 0.01fF
C1973 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n550 GND 0.00fF
C1974 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n551 GND 0.00fF
C1975 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n552 GND 0.00fF
C1976 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n553 GND 0.00fF
C1977 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n554 GND 0.01fF
C1978 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n555 GND 0.01fF
C1979 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n556 GND 0.01fF
C1980 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n557 GND 0.00fF
C1981 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n558 GND 0.00fF
C1982 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n559 GND 0.01fF
C1983 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n560 GND 0.01fF
C1984 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n561 GND 0.01fF
C1985 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n562 GND 0.01fF
C1986 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n563 GND 0.00fF
C1987 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n564 GND 0.00fF
C1988 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n565 GND 0.01fF
C1989 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n566 GND 0.00fF
C1990 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n567 GND 0.01fF
C1991 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n568 GND 0.00fF
C1992 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n569 GND 0.01fF
C1993 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n570 GND 0.01fF
C1994 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n571 GND 0.00fF
C1995 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n572 GND 0.01fF
C1996 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n573 GND 0.00fF
C1997 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n574 GND 0.00fF
C1998 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n575 GND 0.00fF
C1999 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n576 GND 0.00fF
C2000 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n577 GND 0.53fF
C2001 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN GND 0.45fF
C2002 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n578 GND 0.00fF
C2003 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n579 GND 0.00fF
C2004 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n580 GND 0.00fF
C2005 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n581 GND 0.01fF
C2006 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t34 GND 0.13fF $
+ **FLOATING
C2007 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t35 GND 0.13fF $
+ **FLOATING
C2008 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n582 GND 0.37fF
C2009 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n583 GND 0.05fF
C2010 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n584 GND 0.28fF
C2011 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n585 GND 0.01fF
C2012 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n586 GND 0.00fF
C2013 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n587 GND 0.00fF
C2014 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n588 GND 0.00fF
C2015 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n589 GND 0.01fF
C2016 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n590 GND 0.01fF
C2017 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n591 GND 0.00fF
C2018 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n592 GND 0.00fF
C2019 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n593 GND 0.00fF
C2020 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n594 GND 0.01fF
C2021 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n595 GND 0.01fF
C2022 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n596 GND 0.01fF
C2023 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n597 GND 0.01fF
C2024 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n598 GND 0.01fF
C2025 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n599 GND 0.00fF
C2026 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n600 GND 0.00fF
C2027 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n601 GND 0.00fF
C2028 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n602 GND 0.00fF
C2029 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n603 GND 0.01fF
C2030 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n604 GND 0.01fF
C2031 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n605 GND 0.01fF
C2032 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n606 GND 0.00fF
C2033 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n607 GND 0.01fF
C2034 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n608 GND 0.01fF
C2035 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n609 GND 0.00fF
C2036 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n610 GND 0.00fF
C2037 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n611 GND 0.00fF
C2038 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n612 GND 0.00fF
C2039 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n613 GND 0.04fF
C2040 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n614 GND 0.01fF
C2041 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n615 GND 0.01fF
C2042 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n616 GND 0.01fF
C2043 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n617 GND 0.00fF
C2044 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n618 GND 0.00fF
C2045 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n619 GND 0.00fF
C2046 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n620 GND 0.00fF
C2047 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n621 GND 0.01fF
C2048 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n622 GND 0.01fF
C2049 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n623 GND 0.01fF
C2050 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n624 GND 0.00fF
C2051 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n625 GND 0.01fF
C2052 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n626 GND 0.00fF
C2053 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n627 GND 0.00fF
C2054 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n628 GND 0.01fF
C2055 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n629 GND 0.01fF
C2056 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n630 GND 0.01fF
C2057 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n631 GND 0.01fF
C2058 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n632 GND 0.00fF
C2059 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n633 GND 0.00fF
C2060 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n634 GND 0.00fF
C2061 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n635 GND 0.01fF
C2062 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t47 GND 0.13fF $
+ **FLOATING
C2063 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t22 GND 0.13fF $
+ **FLOATING
C2064 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n636 GND 0.37fF
C2065 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n637 GND 0.05fF
C2066 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n638 GND 0.28fF
C2067 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n639 GND 0.01fF
C2068 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n640 GND 0.00fF
C2069 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n641 GND 0.00fF
C2070 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n642 GND 0.00fF
C2071 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n643 GND 0.01fF
C2072 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n644 GND 0.01fF
C2073 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n645 GND 0.00fF
C2074 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n646 GND 0.00fF
C2075 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n647 GND 0.00fF
C2076 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n648 GND 0.00fF
C2077 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n649 GND 0.01fF
C2078 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n650 GND 0.01fF
C2079 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n651 GND 0.01fF
C2080 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n652 GND 0.01fF
C2081 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n653 GND 0.01fF
C2082 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n654 GND 0.00fF
C2083 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n655 GND 0.00fF
C2084 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n656 GND 0.00fF
C2085 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n657 GND 0.00fF
C2086 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n658 GND 0.01fF
C2087 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n659 GND 0.01fF
C2088 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n660 GND 0.01fF
C2089 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n661 GND 0.00fF
C2090 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n662 GND 0.00fF
C2091 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n663 GND 0.01fF
C2092 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n664 GND 0.01fF
C2093 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n665 GND 0.01fF
C2094 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n666 GND 0.01fF
C2095 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n667 GND 0.00fF
C2096 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n668 GND 0.00fF
C2097 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n669 GND 0.01fF
C2098 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n670 GND 0.00fF
C2099 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n671 GND 0.01fF
C2100 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n672 GND 0.00fF
C2101 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n673 GND 0.01fF
C2102 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n674 GND 0.01fF
C2103 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n675 GND 0.00fF
C2104 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n676 GND 0.01fF
C2105 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n677 GND 0.00fF
C2106 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n678 GND 0.00fF
C2107 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n679 GND 0.00fF
C2108 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n680 GND 0.00fF
C2109 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n681 GND 4.87fF
C2110 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n682 GND 2.90fF
C2111 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n683 GND 0.35fF
C2112 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE GND 0.27fF
C2113 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n684 GND 0.00fF
C2114 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n685 GND 0.00fF
C2115 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n686 GND 0.01fF
C2116 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n687 GND 0.00fF
C2117 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n688 GND 0.00fF
C2118 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n689 GND 0.01fF
C2119 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n690 GND 0.01fF
C2120 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n691 GND 0.01fF
C2121 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n692 GND 0.01fF
C2122 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n693 GND 0.00fF
C2123 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n694 GND 0.01fF
C2124 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n695 GND 0.00fF
C2125 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n696 GND 0.01fF
C2126 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n697 GND 0.00fF
C2127 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n698 GND 0.01fF
C2128 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n699 GND 0.00fF
C2129 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n700 GND 0.01fF
C2130 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n701 GND 0.01fF
C2131 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n702 GND 0.00fF
C2132 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n703 GND 0.00fF
C2133 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n704 GND 0.00fF
C2134 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n705 GND 0.00fF
C2135 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n706 GND 0.00fF
C2136 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n707 GND 0.00fF
C2137 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n708 GND 0.00fF
C2138 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n709 GND 0.01fF
C2139 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n710 GND 0.01fF
C2140 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n711 GND 0.01fF
C2141 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n712 GND 0.01fF
C2142 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n713 GND 0.01fF
C2143 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n714 GND 0.00fF
C2144 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n715 GND 0.00fF
C2145 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n716 GND 0.00fF
C2146 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n717 GND 0.00fF
C2147 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n718 GND 0.00fF
C2148 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n719 GND 0.00fF
C2149 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n720 GND 0.01fF
C2150 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n721 GND 0.01fF
C2151 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n722 GND 0.01fF
C2152 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n723 GND 0.01fF
C2153 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n724 GND 0.01fF
C2154 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n725 GND 0.00fF
C2155 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n726 GND 0.00fF
C2156 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n727 GND 0.00fF
C2157 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n728 GND 0.01fF
C2158 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n729 GND 0.01fF
C2159 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t5 GND 0.13fF $
+ **FLOATING
C2160 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n730 GND 0.49fF
C2161 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n731 GND 0.05fF
C2162 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n732 GND 0.28fF
C2163 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n733 GND 0.01fF
C2164 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n734 GND 0.01fF
C2165 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n735 GND 0.00fF
C2166 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n736 GND 0.00fF
C2167 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n737 GND 0.00fF
C2168 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n738 GND 0.00fF
C2169 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n739 GND 0.00fF
C2170 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n740 GND 0.00fF
C2171 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n741 GND 0.01fF
C2172 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n742 GND 0.01fF
C2173 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n743 GND 0.35fF
C2174 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n744 GND 1.56fF
C2175 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n745 GND 0.35fF
C2176 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n746 GND 0.35fF
C2177 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n747 GND 0.44fF
C2178 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n748 GND 0.00fF
C2179 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n749 GND 0.00fF
C2180 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n750 GND 0.00fF
C2181 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n751 GND 0.01fF
C2182 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n752 GND 0.01fF
C2183 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n753 GND 0.01fF
C2184 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n754 GND 0.01fF
C2185 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n755 GND 0.01fF
C2186 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n756 GND 0.00fF
C2187 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n757 GND 0.01fF
C2188 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n758 GND 0.00fF
C2189 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n759 GND 0.00fF
C2190 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n760 GND 0.01fF
C2191 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n761 GND 0.00fF
C2192 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n762 GND 0.01fF
C2193 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n763 GND 0.00fF
C2194 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n764 GND 0.01fF
C2195 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n765 GND 0.01fF
C2196 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n766 GND 0.00fF
C2197 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n767 GND 0.00fF
C2198 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n768 GND 0.00fF
C2199 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n769 GND 0.00fF
C2200 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n770 GND 0.00fF
C2201 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n771 GND 0.00fF
C2202 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n772 GND 0.00fF
C2203 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n773 GND 0.01fF
C2204 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n774 GND 0.01fF
C2205 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n775 GND 0.01fF
C2206 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n776 GND 0.01fF
C2207 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n777 GND 0.01fF
C2208 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n778 GND 0.00fF
C2209 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n779 GND 0.00fF
C2210 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n780 GND 0.00fF
C2211 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n781 GND 0.00fF
C2212 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n782 GND 0.00fF
C2213 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n783 GND 0.01fF
C2214 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n784 GND 0.01fF
C2215 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n785 GND 0.01fF
C2216 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n786 GND 0.01fF
C2217 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n787 GND 0.01fF
C2218 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n788 GND 0.00fF
C2219 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n789 GND 0.00fF
C2220 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n790 GND 0.00fF
C2221 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n791 GND 0.01fF
C2222 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n792 GND 0.01fF
C2223 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t11 GND 0.13fF $
+ **FLOATING
C2224 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n793 GND 0.49fF
C2225 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n794 GND 0.05fF
C2226 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n795 GND 0.28fF
C2227 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n796 GND 0.01fF
C2228 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n797 GND 0.01fF
C2229 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n798 GND 0.00fF
C2230 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n799 GND 0.00fF
C2231 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n800 GND 0.00fF
C2232 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n801 GND 0.00fF
C2233 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n802 GND 0.00fF
C2234 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n803 GND 0.00fF
C2235 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n804 GND 0.01fF
C2236 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n805 GND 0.01fF
C2237 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n806 GND 0.35fF
C2238 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE GND 0.27fF
C2239 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t13 GND 0.13fF $
+ **FLOATING
C2240 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n807 GND 0.49fF
C2241 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n808 GND 0.05fF
C2242 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n809 GND 0.28fF
C2243 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n810 GND 0.01fF
C2244 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n811 GND 0.01fF
C2245 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n812 GND 0.00fF
C2246 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n813 GND 0.00fF
C2247 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n814 GND 0.00fF
C2248 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n815 GND 0.00fF
C2249 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n816 GND 0.00fF
C2250 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n817 GND 0.00fF
C2251 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n818 GND 0.01fF
C2252 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n819 GND 0.01fF
C2253 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n820 GND 0.00fF
C2254 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n821 GND 0.01fF
C2255 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n822 GND 0.01fF
C2256 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n823 GND 0.00fF
C2257 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n824 GND 0.00fF
C2258 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n825 GND 0.00fF
C2259 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n826 GND 0.00fF
C2260 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n827 GND 0.00fF
C2261 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n828 GND 0.00fF
C2262 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n829 GND 0.01fF
C2263 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n830 GND 0.01fF
C2264 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n831 GND 0.01fF
C2265 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n832 GND 0.01fF
C2266 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n833 GND 0.01fF
C2267 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n834 GND 0.00fF
C2268 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n835 GND 0.00fF
C2269 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n836 GND 0.00fF
C2270 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n837 GND 0.01fF
C2271 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n838 GND 0.13fF
C2272 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n839 GND 0.35fF
C2273 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n840 GND 1.53fF
C2274 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n841 GND 0.35fF
C2275 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n842 GND 0.01fF
C2276 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n843 GND 0.45fF
C2277 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n844 GND 0.01fF
C2278 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n845 GND 0.01fF
C2279 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n846 GND 0.01fF
C2280 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n847 GND 0.00fF
C2281 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n848 GND 0.00fF
C2282 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n849 GND 0.00fF
C2283 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n850 GND 0.00fF
C2284 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n851 GND 0.00fF
C2285 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n852 GND 0.01fF
C2286 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n853 GND 0.00fF
C2287 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n854 GND 0.00fF
C2288 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n855 GND 0.01fF
C2289 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n856 GND 0.00fF
C2290 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n857 GND 0.00fF
C2291 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n858 GND 0.00fF
C2292 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n859 GND 0.01fF
C2293 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n860 GND 0.01fF
C2294 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n861 GND 0.01fF
C2295 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n862 GND 0.01fF
C2296 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n863 GND 0.01fF
C2297 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n864 GND 0.00fF
C2298 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n865 GND 0.01fF
C2299 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n866 GND 0.00fF
C2300 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n867 GND 0.01fF
C2301 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n868 GND 0.00fF
C2302 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n869 GND 0.00fF
C2303 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n870 GND 0.00fF
C2304 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n871 GND 0.01fF
C2305 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n872 GND 0.01fF
C2306 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n873 GND 0.01fF
C2307 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n874 GND 0.01fF
C2308 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n875 GND 0.01fF
C2309 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n876 GND 0.00fF
C2310 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n877 GND 0.01fF
C2311 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n878 GND 0.00fF
C2312 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n879 GND 0.01fF
C2313 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n880 GND 0.00fF
C2314 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n881 GND 0.01fF
C2315 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n882 GND 0.00fF
C2316 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n883 GND 0.26fF
C2317 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n884 GND 0.33fF
C2318 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n885 GND 0.00fF
C2319 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n886 GND 0.00fF
C2320 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n887 GND 0.01fF
C2321 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n888 GND 0.01fF
C2322 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n889 GND 0.00fF
C2323 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n890 GND 0.00fF
C2324 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n891 GND 0.00fF
C2325 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n892 GND 0.00fF
C2326 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n893 GND 0.00fF
C2327 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n894 GND 0.00fF
C2328 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n895 GND 0.01fF
C2329 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n896 GND 0.01fF
C2330 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n897 GND 0.01fF
C2331 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n898 GND 0.01fF
C2332 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n899 GND 0.01fF
C2333 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n900 GND 0.00fF
C2334 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n901 GND 0.00fF
C2335 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n902 GND 0.00fF
C2336 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n903 GND 0.00fF
C2337 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n904 GND 0.00fF
C2338 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n905 GND 0.00fF
C2339 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n906 GND 0.01fF
C2340 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n907 GND 0.01fF
C2341 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n908 GND 0.01fF
C2342 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n909 GND 0.01fF
C2343 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n910 GND 0.01fF
C2344 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n911 GND 0.00fF
C2345 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n912 GND 0.00fF
C2346 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n913 GND 0.00fF
C2347 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n914 GND 0.01fF
C2348 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n915 GND 0.01fF
C2349 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t8 GND 0.13fF $
+ **FLOATING
C2350 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t1 GND 0.13fF $
+ **FLOATING
C2351 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n916 GND 0.37fF
C2352 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n917 GND 0.05fF
C2353 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n918 GND 0.28fF
C2354 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n919 GND 0.01fF
C2355 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n920 GND 0.01fF
C2356 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n921 GND 0.00fF
C2357 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n922 GND 0.00fF
C2358 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n923 GND 0.00fF
C2359 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n924 GND 0.00fF
C2360 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n925 GND 0.00fF
C2361 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n926 GND 0.00fF
C2362 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n927 GND 0.01fF
C2363 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n928 GND 0.00fF
C2364 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n929 GND 0.35fF
C2365 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n930 GND 0.40fF
C2366 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n931 GND 1.88fF
C2367 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n932 GND 0.35fF
C2368 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n933 GND 0.08fF
C2369 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n934 GND 0.33fF
C2370 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n935 GND 0.01fF
C2371 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n936 GND 0.00fF
C2372 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n937 GND 0.00fF
C2373 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n938 GND 0.01fF
C2374 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n939 GND 0.01fF
C2375 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n940 GND 0.01fF
C2376 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n941 GND 0.01fF
C2377 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n942 GND 0.00fF
C2378 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n943 GND 0.01fF
C2379 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n944 GND 0.00fF
C2380 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n945 GND 0.00fF
C2381 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n946 GND 0.01fF
C2382 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n947 GND 0.00fF
C2383 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n948 GND 0.01fF
C2384 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n949 GND 0.00fF
C2385 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n950 GND 0.01fF
C2386 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n951 GND 0.01fF
C2387 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n952 GND 0.00fF
C2388 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n953 GND 0.00fF
C2389 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n954 GND 0.00fF
C2390 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n955 GND 0.00fF
C2391 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n956 GND 0.00fF
C2392 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n957 GND 0.00fF
C2393 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n958 GND 0.00fF
C2394 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n959 GND 0.01fF
C2395 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n960 GND 0.01fF
C2396 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n961 GND 0.01fF
C2397 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n962 GND 0.01fF
C2398 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n963 GND 0.01fF
C2399 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n964 GND 0.00fF
C2400 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n965 GND 0.00fF
C2401 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n966 GND 0.00fF
C2402 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n967 GND 0.00fF
C2403 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n968 GND 0.00fF
C2404 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n969 GND 0.00fF
C2405 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n970 GND 0.01fF
C2406 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n971 GND 0.01fF
C2407 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n972 GND 0.01fF
C2408 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n973 GND 0.01fF
C2409 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n974 GND 0.01fF
C2410 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n975 GND 0.00fF
C2411 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n976 GND 0.00fF
C2412 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n977 GND 0.00fF
C2413 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n978 GND 0.00fF
C2414 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n979 GND 0.00fF
C2415 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n980 GND 0.00fF
C2416 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n981 GND 0.00fF
C2417 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n982 GND 0.01fF
C2418 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t7 GND 0.13fF $
+ **FLOATING
C2419 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n983 GND 0.49fF
C2420 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n984 GND 0.05fF
C2421 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n985 GND 0.28fF
C2422 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n986 GND 0.01fF
C2423 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n987 GND 0.00fF
C2424 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n988 GND 0.00fF
C2425 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n989 GND 0.00fF
C2426 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n990 GND 0.01fF
C2427 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n991 GND 0.01fF
C2428 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n992 GND 0.01fF
C2429 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n993 GND 0.01fF
C2430 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n994 GND 0.26fF
C2431 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n995 GND 0.33fF
C2432 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n996 GND 0.01fF
C2433 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n997 GND 0.00fF
C2434 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n998 GND 0.00fF
C2435 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n999 GND 0.01fF
C2436 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1000 GND 0.01fF
C2437 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1001 GND 0.01fF
C2438 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1002 GND 0.01fF
C2439 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1003 GND 0.00fF
C2440 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1004 GND 0.01fF
C2441 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1005 GND 0.00fF
C2442 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1006 GND 0.00fF
C2443 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1007 GND 0.01fF
C2444 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1008 GND 0.00fF
C2445 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1009 GND 0.01fF
C2446 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1010 GND 0.00fF
C2447 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1011 GND 0.00fF
C2448 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1012 GND 0.00fF
C2449 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1013 GND 0.00fF
C2450 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1014 GND 0.01fF
C2451 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t9 GND 0.13fF $
+ **FLOATING
C2452 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t3 GND 0.13fF $
+ **FLOATING
C2453 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1015 GND 0.37fF
C2454 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1016 GND 0.05fF
C2455 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1017 GND 0.28fF
C2456 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1018 GND 0.01fF
C2457 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1019 GND 0.00fF
C2458 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1020 GND 0.00fF
C2459 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1021 GND 0.00fF
C2460 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1022 GND 0.01fF
C2461 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1023 GND 0.01fF
C2462 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1024 GND 0.01fF
C2463 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1025 GND 0.00fF
C2464 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1026 GND 0.00fF
C2465 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1027 GND 0.00fF
C2466 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1028 GND 0.00fF
C2467 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1029 GND 0.00fF
C2468 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1030 GND 0.00fF
C2469 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1031 GND 0.00fF
C2470 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1032 GND 0.01fF
C2471 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1033 GND 0.01fF
C2472 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1034 GND 0.01fF
C2473 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1035 GND 0.01fF
C2474 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1036 GND 0.01fF
C2475 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1037 GND 0.00fF
C2476 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1038 GND 0.00fF
C2477 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1039 GND 0.00fF
C2478 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1040 GND 0.00fF
C2479 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1041 GND 0.00fF
C2480 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1042 GND 0.00fF
C2481 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1043 GND 0.01fF
C2482 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1044 GND 0.01fF
C2483 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1045 GND 0.01fF
C2484 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1046 GND 0.01fF
C2485 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1047 GND 0.01fF
C2486 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1048 GND 0.00fF
C2487 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1049 GND 0.00fF
C2488 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1050 GND 0.00fF
C2489 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1051 GND 0.00fF
C2490 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1052 GND 0.01fF
C2491 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1053 GND 0.01fF
C2492 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1054 GND 0.00fF
C2493 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1055 GND 0.35fF
C2494 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1056 GND 0.40fF
C2495 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1057 GND 4.39fF
C2496 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1058 GND 3.07fF
C2497 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1059 GND 0.01fF
C2498 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t4 GND 0.13fF $
+ **FLOATING
C2499 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1060 GND 0.49fF
C2500 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1061 GND 0.05fF
C2501 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1062 GND 0.28fF
C2502 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1063 GND 0.01fF
C2503 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1064 GND 0.00fF
C2504 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1065 GND 0.00fF
C2505 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1066 GND 0.00fF
C2506 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1067 GND 0.00fF
C2507 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1068 GND 0.00fF
C2508 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1069 GND 0.00fF
C2509 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1070 GND 0.01fF
C2510 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1071 GND 0.01fF
C2511 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1072 GND 0.00fF
C2512 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1073 GND 0.00fF
C2513 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1074 GND 0.01fF
C2514 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1075 GND 0.01fF
C2515 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1076 GND 0.01fF
C2516 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1077 GND 0.01fF
C2517 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1078 GND 0.00fF
C2518 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1079 GND 0.01fF
C2519 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1080 GND 0.00fF
C2520 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1081 GND 0.00fF
C2521 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1082 GND 0.01fF
C2522 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1083 GND 0.00fF
C2523 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1084 GND 0.01fF
C2524 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1085 GND 0.00fF
C2525 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1086 GND 0.01fF
C2526 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1087 GND 0.01fF
C2527 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1088 GND 0.00fF
C2528 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1089 GND 0.00fF
C2529 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1090 GND 0.00fF
C2530 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1091 GND 0.00fF
C2531 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1092 GND 0.00fF
C2532 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1093 GND 0.00fF
C2533 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1094 GND 0.00fF
C2534 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1095 GND 0.01fF
C2535 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1096 GND 0.01fF
C2536 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1097 GND 0.01fF
C2537 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1098 GND 0.01fF
C2538 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1099 GND 0.01fF
C2539 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1100 GND 0.00fF
C2540 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1101 GND 0.00fF
C2541 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1102 GND 0.00fF
C2542 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1103 GND 0.00fF
C2543 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1104 GND 0.00fF
C2544 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1105 GND 0.00fF
C2545 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1106 GND 0.01fF
C2546 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1107 GND 0.01fF
C2547 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1108 GND 0.01fF
C2548 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1109 GND 0.01fF
C2549 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1110 GND 0.01fF
C2550 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1111 GND 0.00fF
C2551 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1112 GND 0.00fF
C2552 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1113 GND 0.00fF
C2553 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1114 GND 0.00fF
C2554 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1115 GND 0.01fF
C2555 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1116 GND 0.01fF
C2556 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1117 GND 0.01fF
C2557 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1118 GND 0.35fF
C2558 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE GND 0.27fF
C2559 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1119 GND 1.88fF
C2560 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1120 GND 0.35fF
C2561 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1121 GND 0.08fF
C2562 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1122 GND 0.33fF
C2563 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1123 GND 0.01fF
C2564 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1124 GND 0.00fF
C2565 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1125 GND 0.00fF
C2566 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1126 GND 0.01fF
C2567 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1127 GND 0.01fF
C2568 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1128 GND 0.01fF
C2569 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1129 GND 0.01fF
C2570 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1130 GND 0.00fF
C2571 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1131 GND 0.01fF
C2572 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1132 GND 0.00fF
C2573 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1133 GND 0.00fF
C2574 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1134 GND 0.01fF
C2575 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1135 GND 0.00fF
C2576 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1136 GND 0.01fF
C2577 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1137 GND 0.00fF
C2578 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1138 GND 0.01fF
C2579 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1139 GND 0.01fF
C2580 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1140 GND 0.00fF
C2581 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1141 GND 0.00fF
C2582 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1142 GND 0.00fF
C2583 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1143 GND 0.00fF
C2584 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1144 GND 0.00fF
C2585 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1145 GND 0.00fF
C2586 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1146 GND 0.00fF
C2587 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1147 GND 0.01fF
C2588 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1148 GND 0.01fF
C2589 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1149 GND 0.01fF
C2590 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1150 GND 0.01fF
C2591 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1151 GND 0.01fF
C2592 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1152 GND 0.00fF
C2593 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1153 GND 0.00fF
C2594 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1154 GND 0.00fF
C2595 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1155 GND 0.00fF
C2596 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1156 GND 0.00fF
C2597 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1157 GND 0.00fF
C2598 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1158 GND 0.01fF
C2599 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1159 GND 0.01fF
C2600 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1160 GND 0.01fF
C2601 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1161 GND 0.01fF
C2602 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1162 GND 0.01fF
C2603 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1163 GND 0.00fF
C2604 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1164 GND 0.00fF
C2605 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1165 GND 0.00fF
C2606 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1166 GND 0.00fF
C2607 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1167 GND 0.00fF
C2608 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1168 GND 0.00fF
C2609 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1169 GND 0.00fF
C2610 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1170 GND 0.01fF
C2611 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t0 GND 0.13fF $
+ **FLOATING
C2612 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1171 GND 0.49fF
C2613 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1172 GND 0.05fF
C2614 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1173 GND 0.28fF
C2615 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1174 GND 0.01fF
C2616 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1175 GND 0.00fF
C2617 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1176 GND 0.00fF
C2618 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1177 GND 0.00fF
C2619 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1178 GND 0.01fF
C2620 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1179 GND 0.01fF
C2621 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1180 GND 0.01fF
C2622 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1181 GND 0.01fF
C2623 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1182 GND 0.26fF
C2624 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1183 GND 0.33fF
C2625 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1184 GND 0.01fF
C2626 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1185 GND 0.00fF
C2627 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1186 GND 0.00fF
C2628 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1187 GND 0.01fF
C2629 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1188 GND 0.01fF
C2630 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1189 GND 0.01fF
C2631 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1190 GND 0.01fF
C2632 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1191 GND 0.00fF
C2633 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1192 GND 0.01fF
C2634 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1193 GND 0.00fF
C2635 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1194 GND 0.00fF
C2636 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1195 GND 0.01fF
C2637 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1196 GND 0.00fF
C2638 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1197 GND 0.01fF
C2639 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1198 GND 0.00fF
C2640 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1199 GND 0.00fF
C2641 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1200 GND 0.00fF
C2642 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1201 GND 0.00fF
C2643 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1202 GND 0.01fF
C2644 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t14 GND 0.13fF $
+ **FLOATING
C2645 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t12 GND 0.13fF $
+ **FLOATING
C2646 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1203 GND 0.37fF
C2647 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1204 GND 0.05fF
C2648 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1205 GND 0.28fF
C2649 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1206 GND 0.01fF
C2650 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1207 GND 0.00fF
C2651 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1208 GND 0.00fF
C2652 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1209 GND 0.00fF
C2653 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1210 GND 0.01fF
C2654 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1211 GND 0.01fF
C2655 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1212 GND 0.01fF
C2656 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1213 GND 0.00fF
C2657 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1214 GND 0.00fF
C2658 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1215 GND 0.00fF
C2659 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1216 GND 0.00fF
C2660 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1217 GND 0.00fF
C2661 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1218 GND 0.00fF
C2662 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1219 GND 0.00fF
C2663 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1220 GND 0.01fF
C2664 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1221 GND 0.01fF
C2665 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1222 GND 0.01fF
C2666 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1223 GND 0.01fF
C2667 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1224 GND 0.01fF
C2668 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1225 GND 0.00fF
C2669 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1226 GND 0.00fF
C2670 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1227 GND 0.00fF
C2671 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1228 GND 0.00fF
C2672 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1229 GND 0.00fF
C2673 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1230 GND 0.00fF
C2674 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1231 GND 0.01fF
C2675 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1232 GND 0.01fF
C2676 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1233 GND 0.01fF
C2677 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1234 GND 0.01fF
C2678 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1235 GND 0.01fF
C2679 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1236 GND 0.00fF
C2680 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1237 GND 0.00fF
C2681 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1238 GND 0.00fF
C2682 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1239 GND 0.00fF
C2683 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1240 GND 0.01fF
C2684 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1241 GND 0.01fF
C2685 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1242 GND 0.00fF
C2686 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1243 GND 0.35fF
C2687 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1244 GND 0.40fF
C2688 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1245 GND 0.01fF
C2689 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t15 GND 0.13fF $
+ **FLOATING
C2690 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1246 GND 0.49fF
C2691 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1247 GND 0.05fF
C2692 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1248 GND 0.28fF
C2693 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1249 GND 0.01fF
C2694 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1250 GND 0.00fF
C2695 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1251 GND 0.00fF
C2696 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1252 GND 0.00fF
C2697 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1253 GND 0.00fF
C2698 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1254 GND 0.00fF
C2699 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1255 GND 0.00fF
C2700 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1256 GND 0.01fF
C2701 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1257 GND 0.01fF
C2702 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1258 GND 0.00fF
C2703 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1259 GND 0.00fF
C2704 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1260 GND 0.01fF
C2705 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1261 GND 0.01fF
C2706 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1262 GND 0.01fF
C2707 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1263 GND 0.01fF
C2708 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1264 GND 0.00fF
C2709 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1265 GND 0.01fF
C2710 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1266 GND 0.00fF
C2711 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1267 GND 0.00fF
C2712 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1268 GND 0.01fF
C2713 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1269 GND 0.00fF
C2714 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1270 GND 0.01fF
C2715 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1271 GND 0.00fF
C2716 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1272 GND 0.01fF
C2717 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1273 GND 0.01fF
C2718 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1274 GND 0.00fF
C2719 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1275 GND 0.00fF
C2720 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1276 GND 0.00fF
C2721 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1277 GND 0.00fF
C2722 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1278 GND 0.00fF
C2723 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1279 GND 0.00fF
C2724 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1280 GND 0.00fF
C2725 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1281 GND 0.01fF
C2726 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1282 GND 0.01fF
C2727 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1283 GND 0.01fF
C2728 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1284 GND 0.01fF
C2729 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1285 GND 0.01fF
C2730 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1286 GND 0.00fF
C2731 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1287 GND 0.00fF
C2732 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1288 GND 0.00fF
C2733 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1289 GND 0.00fF
C2734 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1290 GND 0.00fF
C2735 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1291 GND 0.00fF
C2736 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1292 GND 0.01fF
C2737 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1293 GND 0.01fF
C2738 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1294 GND 0.01fF
C2739 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1295 GND 0.01fF
C2740 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1296 GND 0.01fF
C2741 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1297 GND 0.00fF
C2742 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1298 GND 0.00fF
C2743 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1299 GND 0.00fF
C2744 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1300 GND 0.00fF
C2745 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1301 GND 0.01fF
C2746 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1302 GND 0.01fF
C2747 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1303 GND 0.01fF
C2748 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1304 GND 0.35fF
C2749 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1305 GND 8.40fF
C2750 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1306 GND 0.53fF
C2751 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN GND 0.45fF
C2752 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1307 GND 0.00fF
C2753 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1308 GND 0.00fF
C2754 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1309 GND 0.00fF
C2755 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1310 GND 0.01fF
C2756 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t19 GND 0.13fF $
+ **FLOATING
C2757 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t43 GND 0.13fF $
+ **FLOATING
C2758 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1311 GND 0.37fF
C2759 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1312 GND 0.05fF
C2760 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1313 GND 0.28fF
C2761 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1314 GND 0.01fF
C2762 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1315 GND 0.00fF
C2763 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1316 GND 0.00fF
C2764 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1317 GND 0.00fF
C2765 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1318 GND 0.01fF
C2766 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1319 GND 0.01fF
C2767 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1320 GND 0.00fF
C2768 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1321 GND 0.00fF
C2769 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1322 GND 0.00fF
C2770 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1323 GND 0.01fF
C2771 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1324 GND 0.01fF
C2772 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1325 GND 0.01fF
C2773 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1326 GND 0.01fF
C2774 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1327 GND 0.01fF
C2775 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1328 GND 0.00fF
C2776 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1329 GND 0.00fF
C2777 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1330 GND 0.00fF
C2778 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1331 GND 0.00fF
C2779 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1332 GND 0.01fF
C2780 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1333 GND 0.01fF
C2781 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1334 GND 0.01fF
C2782 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1335 GND 0.00fF
C2783 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1336 GND 0.01fF
C2784 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1337 GND 0.01fF
C2785 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1338 GND 0.00fF
C2786 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1339 GND 0.00fF
C2787 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1340 GND 0.00fF
C2788 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1341 GND 0.00fF
C2789 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1342 GND 0.04fF
C2790 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1343 GND 0.01fF
C2791 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1344 GND 0.01fF
C2792 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1345 GND 0.01fF
C2793 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1346 GND 0.00fF
C2794 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1347 GND 0.00fF
C2795 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1348 GND 0.00fF
C2796 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1349 GND 0.00fF
C2797 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1350 GND 0.01fF
C2798 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1351 GND 0.01fF
C2799 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1352 GND 0.01fF
C2800 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1353 GND 0.00fF
C2801 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1354 GND 0.01fF
C2802 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1355 GND 0.00fF
C2803 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1356 GND 0.00fF
C2804 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1357 GND 0.01fF
C2805 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1358 GND 0.01fF
C2806 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1359 GND 0.01fF
C2807 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1360 GND 0.01fF
C2808 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1361 GND 0.00fF
C2809 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1362 GND 0.00fF
C2810 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1363 GND 0.00fF
C2811 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1364 GND 0.01fF
C2812 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t31 GND 0.13fF $
+ **FLOATING
C2813 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t18 GND 0.13fF $
+ **FLOATING
C2814 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1365 GND 0.37fF
C2815 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1366 GND 0.05fF
C2816 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1367 GND 0.28fF
C2817 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1368 GND 0.01fF
C2818 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1369 GND 0.00fF
C2819 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1370 GND 0.00fF
C2820 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1371 GND 0.00fF
C2821 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1372 GND 0.01fF
C2822 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1373 GND 0.01fF
C2823 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1374 GND 0.00fF
C2824 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1375 GND 0.00fF
C2825 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1376 GND 0.00fF
C2826 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1377 GND 0.00fF
C2827 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1378 GND 0.01fF
C2828 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1379 GND 0.01fF
C2829 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1380 GND 0.01fF
C2830 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1381 GND 0.01fF
C2831 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1382 GND 0.01fF
C2832 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1383 GND 0.00fF
C2833 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1384 GND 0.00fF
C2834 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1385 GND 0.00fF
C2835 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1386 GND 0.00fF
C2836 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1387 GND 0.01fF
C2837 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1388 GND 0.01fF
C2838 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1389 GND 0.01fF
C2839 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1390 GND 0.00fF
C2840 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1391 GND 0.00fF
C2841 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1392 GND 0.01fF
C2842 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1393 GND 0.01fF
C2843 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1394 GND 0.01fF
C2844 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1395 GND 0.01fF
C2845 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1396 GND 0.00fF
C2846 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1397 GND 0.00fF
C2847 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1398 GND 0.01fF
C2848 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1399 GND 0.00fF
C2849 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1400 GND 0.01fF
C2850 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1401 GND 0.00fF
C2851 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1402 GND 0.01fF
C2852 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1403 GND 0.01fF
C2853 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1404 GND 0.00fF
C2854 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1405 GND 0.01fF
C2855 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1406 GND 0.00fF
C2856 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1407 GND 0.00fF
C2857 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1408 GND 0.00fF
C2858 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1409 GND 0.00fF
C2859 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1410 GND 0.53fF
C2860 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN GND 0.45fF
C2861 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1411 GND 0.00fF
C2862 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1412 GND 0.00fF
C2863 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1413 GND 0.00fF
C2864 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1414 GND 0.01fF
C2865 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t26 GND 0.13fF $
+ **FLOATING
C2866 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t39 GND 0.13fF $
+ **FLOATING
C2867 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1415 GND 0.37fF
C2868 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1416 GND 0.05fF
C2869 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1417 GND 0.28fF
C2870 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1418 GND 0.01fF
C2871 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1419 GND 0.00fF
C2872 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1420 GND 0.00fF
C2873 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1421 GND 0.00fF
C2874 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1422 GND 0.01fF
C2875 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1423 GND 0.01fF
C2876 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1424 GND 0.00fF
C2877 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1425 GND 0.00fF
C2878 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1426 GND 0.00fF
C2879 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1427 GND 0.01fF
C2880 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1428 GND 0.01fF
C2881 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1429 GND 0.01fF
C2882 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1430 GND 0.01fF
C2883 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1431 GND 0.01fF
C2884 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1432 GND 0.00fF
C2885 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1433 GND 0.00fF
C2886 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1434 GND 0.00fF
C2887 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1435 GND 0.00fF
C2888 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1436 GND 0.01fF
C2889 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1437 GND 0.01fF
C2890 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1438 GND 0.01fF
C2891 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1439 GND 0.00fF
C2892 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1440 GND 0.01fF
C2893 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1441 GND 0.01fF
C2894 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1442 GND 0.00fF
C2895 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1443 GND 0.00fF
C2896 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1444 GND 0.00fF
C2897 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1445 GND 0.00fF
C2898 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1446 GND 0.04fF
C2899 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1447 GND 0.01fF
C2900 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1448 GND 0.01fF
C2901 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1449 GND 0.01fF
C2902 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1450 GND 0.00fF
C2903 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1451 GND 0.00fF
C2904 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1452 GND 0.00fF
C2905 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1453 GND 0.00fF
C2906 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1454 GND 0.01fF
C2907 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1455 GND 0.01fF
C2908 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1456 GND 0.01fF
C2909 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1457 GND 0.00fF
C2910 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1458 GND 0.01fF
C2911 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1459 GND 0.00fF
C2912 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1460 GND 0.00fF
C2913 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1461 GND 0.01fF
C2914 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1462 GND 0.01fF
C2915 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1463 GND 0.01fF
C2916 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1464 GND 0.01fF
C2917 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1465 GND 0.00fF
C2918 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1466 GND 0.00fF
C2919 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1467 GND 0.00fF
C2920 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1468 GND 0.01fF
C2921 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t41 GND 0.13fF $
+ **FLOATING
C2922 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t16 GND 0.13fF $
+ **FLOATING
C2923 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1469 GND 0.37fF
C2924 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1470 GND 0.05fF
C2925 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1471 GND 0.28fF
C2926 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1472 GND 0.01fF
C2927 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1473 GND 0.00fF
C2928 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1474 GND 0.00fF
C2929 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1475 GND 0.00fF
C2930 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1476 GND 0.01fF
C2931 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1477 GND 0.01fF
C2932 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1478 GND 0.00fF
C2933 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1479 GND 0.00fF
C2934 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1480 GND 0.00fF
C2935 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1481 GND 0.00fF
C2936 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1482 GND 0.01fF
C2937 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1483 GND 0.01fF
C2938 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1484 GND 0.01fF
C2939 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1485 GND 0.01fF
C2940 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1486 GND 0.01fF
C2941 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1487 GND 0.00fF
C2942 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1488 GND 0.00fF
C2943 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1489 GND 0.00fF
C2944 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1490 GND 0.00fF
C2945 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1491 GND 0.01fF
C2946 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1492 GND 0.01fF
C2947 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1493 GND 0.01fF
C2948 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1494 GND 0.00fF
C2949 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1495 GND 0.00fF
C2950 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1496 GND 0.01fF
C2951 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1497 GND 0.01fF
C2952 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1498 GND 0.01fF
C2953 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1499 GND 0.01fF
C2954 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1500 GND 0.00fF
C2955 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1501 GND 0.00fF
C2956 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1502 GND 0.01fF
C2957 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1503 GND 0.00fF
C2958 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1504 GND 0.01fF
C2959 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1505 GND 0.00fF
C2960 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1506 GND 0.01fF
C2961 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1507 GND 0.01fF
C2962 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1508 GND 0.00fF
C2963 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1509 GND 0.01fF
C2964 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1510 GND 0.00fF
C2965 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1511 GND 0.00fF
C2966 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1512 GND 0.00fF
C2967 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1513 GND 0.00fF
C2968 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1514 GND 0.53fF
C2969 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN GND 0.45fF
C2970 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1515 GND 0.00fF
C2971 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1516 GND 0.00fF
C2972 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1517 GND 0.00fF
C2973 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1518 GND 0.01fF
C2974 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t28 GND 0.13fF $
+ **FLOATING
C2975 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t32 GND 0.13fF $
+ **FLOATING
C2976 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1519 GND 0.37fF
C2977 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1520 GND 0.05fF
C2978 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1521 GND 0.28fF
C2979 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1522 GND 0.01fF
C2980 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1523 GND 0.00fF
C2981 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1524 GND 0.00fF
C2982 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1525 GND 0.00fF
C2983 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1526 GND 0.01fF
C2984 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1527 GND 0.01fF
C2985 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1528 GND 0.00fF
C2986 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1529 GND 0.00fF
C2987 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1530 GND 0.00fF
C2988 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1531 GND 0.01fF
C2989 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1532 GND 0.01fF
C2990 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1533 GND 0.01fF
C2991 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1534 GND 0.01fF
C2992 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1535 GND 0.01fF
C2993 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1536 GND 0.00fF
C2994 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1537 GND 0.00fF
C2995 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1538 GND 0.00fF
C2996 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1539 GND 0.00fF
C2997 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1540 GND 0.01fF
C2998 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1541 GND 0.01fF
C2999 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1542 GND 0.01fF
C3000 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1543 GND 0.00fF
C3001 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1544 GND 0.01fF
C3002 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1545 GND 0.01fF
C3003 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1546 GND 0.00fF
C3004 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1547 GND 0.00fF
C3005 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1548 GND 0.00fF
C3006 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1549 GND 0.00fF
C3007 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1550 GND 0.04fF
C3008 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1551 GND 0.01fF
C3009 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1552 GND 0.01fF
C3010 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1553 GND 0.01fF
C3011 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1554 GND 0.00fF
C3012 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1555 GND 0.00fF
C3013 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1556 GND 0.00fF
C3014 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1557 GND 0.00fF
C3015 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1558 GND 0.01fF
C3016 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1559 GND 0.01fF
C3017 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1560 GND 0.01fF
C3018 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1561 GND 0.00fF
C3019 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1562 GND 0.01fF
C3020 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1563 GND 0.00fF
C3021 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1564 GND 0.00fF
C3022 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1565 GND 0.01fF
C3023 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1566 GND 0.01fF
C3024 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1567 GND 0.01fF
C3025 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1568 GND 0.01fF
C3026 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1569 GND 0.00fF
C3027 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1570 GND 0.00fF
C3028 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1571 GND 0.00fF
C3029 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1572 GND 0.01fF
C3030 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t33 GND 0.13fF $
+ **FLOATING
C3031 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t21 GND 0.13fF $
+ **FLOATING
C3032 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1573 GND 0.37fF
C3033 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1574 GND 0.05fF
C3034 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1575 GND 0.28fF
C3035 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1576 GND 0.01fF
C3036 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1577 GND 0.00fF
C3037 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1578 GND 0.00fF
C3038 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1579 GND 0.00fF
C3039 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1580 GND 0.01fF
C3040 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1581 GND 0.01fF
C3041 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1582 GND 0.00fF
C3042 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1583 GND 0.00fF
C3043 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1584 GND 0.00fF
C3044 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1585 GND 0.00fF
C3045 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1586 GND 0.01fF
C3046 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1587 GND 0.01fF
C3047 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1588 GND 0.01fF
C3048 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1589 GND 0.01fF
C3049 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1590 GND 0.01fF
C3050 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1591 GND 0.00fF
C3051 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1592 GND 0.00fF
C3052 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1593 GND 0.00fF
C3053 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1594 GND 0.00fF
C3054 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1595 GND 0.01fF
C3055 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1596 GND 0.01fF
C3056 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1597 GND 0.01fF
C3057 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1598 GND 0.00fF
C3058 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1599 GND 0.00fF
C3059 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1600 GND 0.01fF
C3060 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1601 GND 0.01fF
C3061 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1602 GND 0.01fF
C3062 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1603 GND 0.01fF
C3063 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1604 GND 0.00fF
C3064 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1605 GND 0.00fF
C3065 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1606 GND 0.01fF
C3066 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1607 GND 0.00fF
C3067 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1608 GND 0.01fF
C3068 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1609 GND 0.00fF
C3069 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1610 GND 0.01fF
C3070 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1611 GND 0.01fF
C3071 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1612 GND 0.00fF
C3072 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1613 GND 0.01fF
C3073 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1614 GND 0.00fF
C3074 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1615 GND 0.00fF
C3075 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1616 GND 0.00fF
C3076 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1617 GND 0.00fF
C3077 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1618 GND 0.53fF
C3078 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN GND 0.45fF
C3079 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1619 GND 0.00fF
C3080 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1620 GND 0.00fF
C3081 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1621 GND 0.00fF
C3082 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1622 GND 0.01fF
C3083 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t29 GND 0.13fF $
+ **FLOATING
C3084 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t30 GND 0.13fF $
+ **FLOATING
C3085 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1623 GND 0.37fF
C3086 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1624 GND 0.05fF
C3087 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1625 GND 0.28fF
C3088 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1626 GND 0.01fF
C3089 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1627 GND 0.00fF
C3090 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1628 GND 0.00fF
C3091 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1629 GND 0.00fF
C3092 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1630 GND 0.01fF
C3093 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1631 GND 0.01fF
C3094 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1632 GND 0.00fF
C3095 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1633 GND 0.00fF
C3096 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1634 GND 0.00fF
C3097 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1635 GND 0.01fF
C3098 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1636 GND 0.01fF
C3099 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1637 GND 0.01fF
C3100 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1638 GND 0.01fF
C3101 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1639 GND 0.01fF
C3102 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1640 GND 0.00fF
C3103 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1641 GND 0.00fF
C3104 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1642 GND 0.00fF
C3105 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1643 GND 0.00fF
C3106 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1644 GND 0.01fF
C3107 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1645 GND 0.01fF
C3108 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1646 GND 0.01fF
C3109 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1647 GND 0.00fF
C3110 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1648 GND 0.01fF
C3111 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1649 GND 0.01fF
C3112 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1650 GND 0.00fF
C3113 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1651 GND 0.00fF
C3114 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1652 GND 0.00fF
C3115 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1653 GND 0.00fF
C3116 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1654 GND 0.04fF
C3117 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1655 GND 0.01fF
C3118 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1656 GND 0.01fF
C3119 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1657 GND 0.01fF
C3120 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1658 GND 0.00fF
C3121 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1659 GND 0.00fF
C3122 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1660 GND 0.00fF
C3123 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1661 GND 0.00fF
C3124 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1662 GND 0.01fF
C3125 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1663 GND 0.01fF
C3126 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1664 GND 0.01fF
C3127 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1665 GND 0.00fF
C3128 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1666 GND 0.01fF
C3129 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1667 GND 0.00fF
C3130 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1668 GND 0.00fF
C3131 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1669 GND 0.01fF
C3132 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1670 GND 0.01fF
C3133 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1671 GND 0.01fF
C3134 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1672 GND 0.01fF
C3135 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1673 GND 0.00fF
C3136 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1674 GND 0.00fF
C3137 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1675 GND 0.00fF
C3138 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1676 GND 0.01fF
C3139 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t42 GND 0.13fF $
+ **FLOATING
C3140 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t17 GND 0.13fF $
+ **FLOATING
C3141 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1677 GND 0.37fF
C3142 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1678 GND 0.05fF
C3143 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1679 GND 0.28fF
C3144 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1680 GND 0.01fF
C3145 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1681 GND 0.00fF
C3146 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1682 GND 0.00fF
C3147 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1683 GND 0.00fF
C3148 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1684 GND 0.01fF
C3149 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1685 GND 0.01fF
C3150 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1686 GND 0.00fF
C3151 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1687 GND 0.00fF
C3152 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1688 GND 0.00fF
C3153 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1689 GND 0.00fF
C3154 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1690 GND 0.01fF
C3155 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1691 GND 0.01fF
C3156 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1692 GND 0.01fF
C3157 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1693 GND 0.01fF
C3158 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1694 GND 0.01fF
C3159 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1695 GND 0.00fF
C3160 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1696 GND 0.00fF
C3161 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1697 GND 0.00fF
C3162 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1698 GND 0.00fF
C3163 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1699 GND 0.01fF
C3164 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1700 GND 0.01fF
C3165 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1701 GND 0.01fF
C3166 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1702 GND 0.00fF
C3167 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1703 GND 0.00fF
C3168 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1704 GND 0.01fF
C3169 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1705 GND 0.01fF
C3170 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1706 GND 0.01fF
C3171 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1707 GND 0.01fF
C3172 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1708 GND 0.00fF
C3173 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1709 GND 0.00fF
C3174 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1710 GND 0.01fF
C3175 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1711 GND 0.00fF
C3176 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1712 GND 0.01fF
C3177 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1713 GND 0.00fF
C3178 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1714 GND 0.01fF
C3179 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1715 GND 0.01fF
C3180 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1716 GND 0.00fF
C3181 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1717 GND 0.01fF
C3182 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1718 GND 0.00fF
C3183 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1719 GND 0.00fF
C3184 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1720 GND 0.00fF
C3185 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1721 GND 0.00fF
C3186 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1722 GND 11.36fF
C3187 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1723 GND 0.29fF
C3188 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t24 GND 0.13fF $
+ **FLOATING
C3189 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.t46 GND 0.13fF $
+ **FLOATING
C3190 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1724 GND 0.37fF
C3191 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1725 GND 0.05fF
C3192 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1726 GND 0.28fF
C3193 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1727 GND 0.01fF
C3194 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1728 GND 0.01fF
C3195 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1729 GND 0.00fF
C3196 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1730 GND 0.00fF
C3197 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1731 GND 0.00fF
C3198 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1732 GND 0.00fF
C3199 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1733 GND 0.00fF
C3200 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1734 GND 0.00fF
C3201 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1735 GND 0.01fF
C3202 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1736 GND 0.01fF
C3203 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1737 GND 0.01fF
C3204 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1738 GND 0.00fF
C3205 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1739 GND 0.00fF
C3206 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1740 GND 0.00fF
C3207 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1741 GND 0.00fF
C3208 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1742 GND 0.01fF
C3209 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1743 GND 0.01fF
C3210 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1744 GND 0.01fF
C3211 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1745 GND 0.01fF
C3212 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1746 GND 0.01fF
C3213 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1747 GND 0.00fF
C3214 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1748 GND 0.00fF
C3215 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1749 GND 0.00fF
C3216 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1750 GND 0.00fF
C3217 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1751 GND 0.01fF
C3218 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1752 GND 0.01fF
C3219 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1753 GND 0.01fF
C3220 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1754 GND 0.53fF
C3221 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN GND 0.45fF
C3222 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1755 GND 1.12fF
C3223 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1756 GND 1.12fF
C3224 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1757 GND 1.12fF
C3225 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1758 GND 1.12fF
C3226 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1759 GND 1.12fF
C3227 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1760 GND 1.12fF
C3228 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE.n1761 GND 1.12fF
C3229 VBIAS.n0 GND 0.01fF
C3230 VBIAS.n1 GND 0.00fF
C3231 VBIAS.n2 GND 0.01fF
C3232 VBIAS.n3 GND 0.01fF
C3233 VBIAS.n4 GND 0.00fF
C3234 VBIAS.n5 GND 0.01fF
C3235 VBIAS.n6 GND 0.01fF
C3236 VBIAS.n7 GND 0.01fF
C3237 VBIAS.n8 GND 0.00fF
C3238 VBIAS.n9 GND 0.01fF
C3239 VBIAS.n10 GND 0.00fF
C3240 VBIAS.n11 GND 0.01fF
C3241 VBIAS.n13 GND 1.34fF
C3242 VBIAS.n14 GND 0.06fF
C3243 VBIAS.n15 GND 0.01fF
C3244 VBIAS.n16 GND 0.00fF
C3245 VBIAS.n17 GND 0.01fF
C3246 VBIAS.n18 GND 0.01fF
C3247 VBIAS.t7 GND 0.17fF $ **FLOATING
C3248 VBIAS.t1 GND 0.17fF $ **FLOATING
C3249 VBIAS.n19 GND 0.51fF
C3250 VBIAS.n20 GND 0.07fF
C3251 VBIAS.n21 GND 0.39fF
C3252 VBIAS.n22 GND 0.01fF
C3253 VBIAS.n23 GND 0.00fF
C3254 VBIAS.n24 GND 0.00fF
C3255 VBIAS.n25 GND 0.01fF
C3256 VBIAS.n26 GND 0.01fF
C3257 VBIAS.n27 GND 0.00fF
C3258 VBIAS.n28 GND 0.00fF
C3259 VBIAS.n29 GND 0.00fF
C3260 VBIAS.n30 GND 0.01fF
C3261 VBIAS.n31 GND 0.01fF
C3262 VBIAS.n32 GND 0.01fF
C3263 VBIAS.n33 GND 0.01fF
C3264 VBIAS.n34 GND 0.01fF
C3265 VBIAS.n35 GND 0.00fF
C3266 VBIAS.n36 GND 0.01fF
C3267 VBIAS.n37 GND 0.00fF
C3268 VBIAS.n38 GND 0.00fF
C3269 VBIAS.n39 GND 0.00fF
C3270 VBIAS.n40 GND 0.00fF
C3271 VBIAS.n41 GND 0.00fF
C3272 VBIAS.n42 GND 0.01fF
C3273 VBIAS.n43 GND 0.01fF
C3274 VBIAS.n44 GND 0.01fF
C3275 VBIAS.n45 GND 0.01fF
C3276 VBIAS.n46 GND 0.01fF
C3277 VBIAS.n47 GND 0.00fF
C3278 VBIAS.n48 GND 0.01fF
C3279 VBIAS.n49 GND 0.00fF
C3280 VBIAS.n50 GND 0.00fF
C3281 VBIAS.n51 GND 0.00fF
C3282 VBIAS.n52 GND 0.00fF
C3283 VBIAS.n53 GND 0.00fF
C3284 VBIAS.n54 GND 0.00fF
C3285 VBIAS.n55 GND 0.01fF
C3286 VBIAS.n56 GND 0.01fF
C3287 VBIAS.n57 GND 0.01fF
C3288 VBIAS.n58 GND 0.06fF
C3289 VBIAS.n59 GND 0.06fF
C3290 VBIAS.n61 GND 0.01fF
C3291 VBIAS.n62 GND 0.01fF
C3292 VBIAS.n63 GND 0.00fF
C3293 VBIAS.n64 GND 0.00fF
C3294 VBIAS.n65 GND 0.02fF
C3295 VBIAS.n66 GND 0.02fF
C3296 VBIAS.n67 GND 0.00fF
C3297 VBIAS.n68 GND 0.00fF
C3298 VBIAS.n70 GND 0.00fF
C3299 VBIAS.n71 GND 0.00fF
C3300 VBIAS.n72 GND 0.00fF
C3301 VBIAS.n73 GND 0.01fF
C3302 VBIAS.n74 GND 0.00fF
C3303 VBIAS.n75 GND 0.01fF
C3304 VBIAS.n76 GND 0.01fF
C3305 VBIAS.n77 GND 0.00fF
C3306 VBIAS.n78 GND 0.01fF
C3307 VBIAS.n79 GND 0.01fF
C3308 VBIAS.n80 GND 0.00fF
C3309 VBIAS.n81 GND 0.01fF
C3310 VBIAS.n82 GND 0.01fF
C3311 VBIAS.n83 GND 0.01fF
C3312 VBIAS.n84 GND 0.00fF
C3313 VBIAS.n85 GND 0.01fF
C3314 VBIAS.n86 GND 0.00fF
C3315 VBIAS.n87 GND 0.01fF
C3316 VBIAS.n89 GND 0.15fF
C3317 VBIAS.n90 GND 0.24fF
C3318 VBIAS.n91 GND 0.27fF
C3319 VBIAS.n92 GND 0.06fF
C3320 VBIAS.n93 GND 0.06fF
C3321 VBIAS.n94 GND 0.06fF
C3322 VBIAS.n95 GND 0.07fF
C3323 VBIAS.n97 GND 0.12fF
C3324 VBIAS.n99 GND 0.12fF
C3325 VBIAS.n101 GND 0.10fF
C3326 VBIAS.n103 GND 0.10fF
C3327 VBIAS.n105 GND 1.06fF
C3328 VBIAS.n107 GND 0.19fF
C3329 VBIAS.n109 GND 0.25fF
C3330 VBIAS.n110 GND 0.06fF
C3331 VBIAS.n111 GND 0.06fF
C3332 VBIAS.n112 GND 0.06fF
C3333 VBIAS.n113 GND 0.07fF
C3334 VBIAS.n115 GND 0.12fF
C3335 VBIAS.n116 GND 0.01fF
C3336 VBIAS.n117 GND 0.01fF
C3337 VBIAS.n118 GND 0.01fF
C3338 VBIAS.n119 GND 0.01fF
C3339 VBIAS.n120 GND 0.03fF
C3340 VBIAS.n121 GND 0.03fF
C3341 VBIAS.n122 GND 0.01fF
C3342 VBIAS.n123 GND 0.04fF
C3343 VBIAS.n124 GND 0.01fF
C3344 VBIAS.n125 GND 0.01fF
C3345 VBIAS.n126 GND 0.01fF
C3346 VBIAS.n127 GND 0.00fF
C3347 VBIAS.n128 GND 0.01fF
C3348 VBIAS.n129 GND 0.00fF
C3349 VBIAS.n130 GND 0.12fF
C3350 VBIAS.n131 GND 0.01fF
C3351 VBIAS.n132 GND 0.01fF
C3352 VBIAS.n133 GND 0.02fF
C3353 VBIAS.n134 GND 0.00fF
C3354 VBIAS.n135 GND 0.01fF
C3355 VBIAS.n136 GND 0.00fF
C3356 VBIAS.n137 GND 0.01fF
C3357 VBIAS.n138 GND 0.01fF
C3358 VBIAS.n139 GND 0.01fF
C3359 VBIAS.n140 GND 0.01fF
C3360 VBIAS.n141 GND 0.01fF
C3361 VBIAS.n142 GND 0.01fF
C3362 VBIAS.n143 GND 0.03fF
C3363 VBIAS.n144 GND 0.12fF
C3364 VBIAS.n145 GND 0.02fF
C3365 VBIAS.n146 GND 0.04fF
C3366 VBIAS.n147 GND 0.01fF
C3367 VBIAS.n148 GND 0.01fF
C3368 VBIAS.n149 GND 0.01fF
C3369 VBIAS.n150 GND 0.01fF
C3370 VBIAS.n151 GND 0.03fF
C3371 VBIAS.n152 GND 0.02fF
C3372 VBIAS.n153 GND 0.01fF
C3373 VBIAS.n154 GND 0.01fF
C3374 VBIAS.n155 GND 0.00fF
C3375 VBIAS.n156 GND 0.00fF
C3376 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE GND 0.00fF
C3377 VBIAS.n157 GND 0.01fF
C3378 VBIAS.n158 GND 0.01fF
C3379 VBIAS.n159 GND 0.01fF
C3380 VBIAS.n160 GND 0.00fF
C3381 VBIAS.n161 GND 0.01fF
C3382 VBIAS.n162 GND 0.04fF
C3383 VBIAS.n163 GND 0.00fF
C3384 VBIAS.n164 GND 0.01fF
C3385 VBIAS.n165 GND 0.01fF
C3386 VBIAS.n166 GND 0.01fF
C3387 VBIAS.n167 GND 0.00fF
C3388 VBIAS.n168 GND 0.00fF
C3389 VBIAS.n169 GND 0.00fF
C3390 VBIAS.n170 GND 0.01fF
C3391 VBIAS.n171 GND 0.01fF
C3392 VBIAS.n172 GND 0.02fF
C3393 VBIAS.n173 GND 0.02fF
C3394 VBIAS.n174 GND 0.01fF
C3395 VBIAS.n175 GND 0.01fF
C3396 VBIAS.n176 GND 0.03fF
C3397 VBIAS.n177 GND 0.12fF
C3398 VBIAS.n178 GND 0.02fF
C3399 VBIAS.n179 GND 0.04fF
C3400 VBIAS.n180 GND 0.01fF
C3401 VBIAS.n181 GND 0.01fF
C3402 VBIAS.n182 GND 0.00fF
C3403 VBIAS.n183 GND 0.01fF
C3404 VBIAS.n184 GND 0.00fF
C3405 VBIAS.n185 GND 0.12fF
C3406 VBIAS.n186 GND 0.01fF
C3407 VBIAS.n187 GND 0.01fF
C3408 VBIAS.n188 GND 0.02fF
C3409 VBIAS.n189 GND 0.00fF
C3410 VBIAS.n190 GND 0.01fF
C3411 VBIAS.n191 GND 0.00fF
C3412 VBIAS.n192 GND 0.01fF
C3413 VBIAS.n193 GND 0.01fF
C3414 VBIAS.n194 GND 0.01fF
C3415 VBIAS.n195 GND 0.01fF
C3416 VBIAS.n196 GND 0.01fF
C3417 VBIAS.n197 GND 0.01fF
C3418 VBIAS.n198 GND 0.01fF
C3419 VBIAS.n199 GND 0.01fF
C3420 VBIAS.n200 GND 0.05fF
C3421 VBIAS.n201 GND 0.10fF
C3422 VBIAS.n202 GND 0.01fF
C3423 VBIAS.n203 GND 0.04fF
C3424 VBIAS.n204 GND 0.04fF
C3425 VBIAS.n205 GND 0.01fF
C3426 VBIAS.n206 GND 0.04fF
C3427 VBIAS.n207 GND 0.03fF
C3428 VBIAS.n208 GND 0.01fF
C3429 VBIAS.n209 GND 0.17fF
C3430 VBIAS.n210 GND 0.01fF
C3431 VBIAS.n211 GND 0.01fF
C3432 VBIAS.n212 GND 0.01fF
C3433 VBIAS.n213 GND 0.03fF
C3434 VBIAS.n214 GND 0.03fF
C3435 VBIAS.n215 GND 0.01fF
C3436 VBIAS.n216 GND 0.04fF
C3437 VBIAS.n217 GND 0.01fF
C3438 VBIAS.n218 GND 0.01fF
C3439 VBIAS.n219 GND 0.01fF
C3440 VBIAS.n220 GND 0.00fF
C3441 VBIAS.n221 GND 0.01fF
C3442 VBIAS.n222 GND 0.00fF
C3443 VBIAS.n223 GND 0.12fF
C3444 VBIAS.n224 GND 0.01fF
C3445 VBIAS.n225 GND 0.01fF
C3446 VBIAS.n226 GND 0.02fF
C3447 VBIAS.n227 GND 0.00fF
C3448 VBIAS.n228 GND 0.01fF
C3449 VBIAS.n229 GND 0.00fF
C3450 VBIAS.n230 GND 0.01fF
C3451 VBIAS.n231 GND 0.01fF
C3452 VBIAS.n232 GND 0.01fF
C3453 VBIAS.n233 GND 0.01fF
C3454 VBIAS.n234 GND 0.01fF
C3455 VBIAS.n235 GND 0.01fF
C3456 VBIAS.n236 GND 0.03fF
C3457 VBIAS.n237 GND 0.12fF
C3458 VBIAS.n238 GND 0.02fF
C3459 VBIAS.n239 GND 0.04fF
C3460 VBIAS.n240 GND 0.01fF
C3461 VBIAS.n241 GND 0.01fF
C3462 VBIAS.n242 GND 0.01fF
C3463 VBIAS.n243 GND 0.01fF
C3464 VBIAS.n244 GND 0.03fF
C3465 VBIAS.n245 GND 0.02fF
C3466 VBIAS.n246 GND 0.01fF
C3467 VBIAS.n247 GND 0.01fF
C3468 VBIAS.n248 GND 0.00fF
C3469 VBIAS.n249 GND 0.00fF
C3470 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE GND 0.00fF
C3471 VBIAS.n250 GND 0.01fF
C3472 VBIAS.n251 GND 0.01fF
C3473 VBIAS.n252 GND 0.01fF
C3474 VBIAS.n253 GND 0.00fF
C3475 VBIAS.n254 GND 0.01fF
C3476 VBIAS.n255 GND 0.04fF
C3477 VBIAS.n256 GND 0.00fF
C3478 VBIAS.n257 GND 0.01fF
C3479 VBIAS.n258 GND 0.01fF
C3480 VBIAS.n259 GND 0.01fF
C3481 VBIAS.n260 GND 0.01fF
C3482 VBIAS.n261 GND 0.00fF
C3483 VBIAS.n262 GND 0.00fF
C3484 VBIAS.n263 GND 0.00fF
C3485 VBIAS.n264 GND 0.01fF
C3486 VBIAS.n265 GND 0.01fF
C3487 VBIAS.n266 GND 0.02fF
C3488 VBIAS.n267 GND 0.02fF
C3489 VBIAS.n268 GND 0.01fF
C3490 VBIAS.n269 GND 0.03fF
C3491 VBIAS.n270 GND 0.12fF
C3492 VBIAS.n271 GND 0.01fF
C3493 VBIAS.n272 GND 0.02fF
C3494 VBIAS.n273 GND 0.04fF
C3495 VBIAS.n274 GND 0.01fF
C3496 VBIAS.n275 GND 0.01fF
C3497 VBIAS.n276 GND 0.00fF
C3498 VBIAS.n277 GND 0.01fF
C3499 VBIAS.n278 GND 0.00fF
C3500 VBIAS.n279 GND 0.12fF
C3501 VBIAS.n280 GND 0.01fF
C3502 VBIAS.n281 GND 0.01fF
C3503 VBIAS.n282 GND 0.02fF
C3504 VBIAS.n283 GND 0.00fF
C3505 VBIAS.n284 GND 0.01fF
C3506 VBIAS.n285 GND 0.00fF
C3507 VBIAS.n286 GND 0.01fF
C3508 VBIAS.n287 GND 0.01fF
C3509 VBIAS.n288 GND 0.01fF
C3510 VBIAS.n289 GND 0.01fF
C3511 VBIAS.n290 GND 0.01fF
C3512 VBIAS.n291 GND 0.01fF
C3513 VBIAS.n292 GND 0.01fF
C3514 VBIAS.n293 GND 0.01fF
C3515 VBIAS.n294 GND 0.05fF
C3516 VBIAS.n295 GND 0.17fF
C3517 VBIAS.n296 GND 0.03fF
C3518 VBIAS.n297 GND 0.03fF
C3519 VBIAS.n298 GND 0.01fF
C3520 VBIAS.n299 GND 0.04fF
C3521 VBIAS.n300 GND 0.04fF
C3522 VBIAS.n301 GND 0.01fF
C3523 VBIAS.n302 GND 0.04fF
C3524 VBIAS.n303 GND 0.03fF
C3525 VBIAS.n304 GND 0.01fF
C3526 VBIAS.n305 GND 0.46fF
C3527 VBIAS.n306 GND 0.01fF
C3528 VBIAS.n307 GND 0.01fF
C3529 VBIAS.n308 GND 0.01fF
C3530 VBIAS.n309 GND 0.03fF
C3531 VBIAS.n310 GND 0.03fF
C3532 VBIAS.n311 GND 0.01fF
C3533 VBIAS.n312 GND 0.04fF
C3534 VBIAS.n313 GND 0.01fF
C3535 VBIAS.n314 GND 0.01fF
C3536 VBIAS.n315 GND 0.01fF
C3537 VBIAS.n316 GND 0.00fF
C3538 VBIAS.n317 GND 0.01fF
C3539 VBIAS.n318 GND 0.00fF
C3540 VBIAS.n319 GND 0.12fF
C3541 VBIAS.n320 GND 0.01fF
C3542 VBIAS.n321 GND 0.01fF
C3543 VBIAS.n322 GND 0.02fF
C3544 VBIAS.n323 GND 0.00fF
C3545 VBIAS.n324 GND 0.01fF
C3546 VBIAS.n325 GND 0.00fF
C3547 VBIAS.n326 GND 0.01fF
C3548 VBIAS.n327 GND 0.01fF
C3549 VBIAS.n328 GND 0.01fF
C3550 VBIAS.n329 GND 0.01fF
C3551 VBIAS.n330 GND 0.01fF
C3552 VBIAS.n331 GND 0.01fF
C3553 VBIAS.n332 GND 0.03fF
C3554 VBIAS.n333 GND 0.12fF
C3555 VBIAS.n334 GND 0.02fF
C3556 VBIAS.n335 GND 0.04fF
C3557 VBIAS.n336 GND 0.01fF
C3558 VBIAS.n337 GND 0.01fF
C3559 VBIAS.n338 GND 0.01fF
C3560 VBIAS.n339 GND 0.01fF
C3561 VBIAS.n340 GND 0.03fF
C3562 VBIAS.n341 GND 0.02fF
C3563 VBIAS.n342 GND 0.01fF
C3564 VBIAS.n343 GND 0.01fF
C3565 VBIAS.n344 GND 0.00fF
C3566 VBIAS.n345 GND 0.00fF
C3567 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE GND 0.00fF
C3568 VBIAS.n346 GND 0.01fF
C3569 VBIAS.n347 GND 0.01fF
C3570 VBIAS.n348 GND 0.01fF
C3571 VBIAS.n349 GND 0.00fF
C3572 VBIAS.n350 GND 0.01fF
C3573 VBIAS.n351 GND 0.04fF
C3574 VBIAS.n352 GND 0.00fF
C3575 VBIAS.n353 GND 0.01fF
C3576 VBIAS.n354 GND 0.01fF
C3577 VBIAS.n355 GND 0.01fF
C3578 VBIAS.n356 GND 0.01fF
C3579 VBIAS.n357 GND 0.00fF
C3580 VBIAS.n358 GND 0.00fF
C3581 VBIAS.n359 GND 0.00fF
C3582 VBIAS.n360 GND 0.01fF
C3583 VBIAS.n361 GND 0.01fF
C3584 VBIAS.n362 GND 0.02fF
C3585 VBIAS.n363 GND 0.02fF
C3586 VBIAS.n364 GND 0.01fF
C3587 VBIAS.n365 GND 0.03fF
C3588 VBIAS.n366 GND 0.12fF
C3589 VBIAS.n367 GND 0.01fF
C3590 VBIAS.n368 GND 0.02fF
C3591 VBIAS.n369 GND 0.04fF
C3592 VBIAS.n370 GND 0.01fF
C3593 VBIAS.n371 GND 0.01fF
C3594 VBIAS.n372 GND 0.00fF
C3595 VBIAS.n373 GND 0.01fF
C3596 VBIAS.n374 GND 0.00fF
C3597 VBIAS.n375 GND 0.12fF
C3598 VBIAS.n376 GND 0.01fF
C3599 VBIAS.n377 GND 0.01fF
C3600 VBIAS.n378 GND 0.02fF
C3601 VBIAS.n379 GND 0.00fF
C3602 VBIAS.n380 GND 0.01fF
C3603 VBIAS.n381 GND 0.00fF
C3604 VBIAS.n382 GND 0.01fF
C3605 VBIAS.n383 GND 0.01fF
C3606 VBIAS.n384 GND 0.01fF
C3607 VBIAS.n385 GND 0.01fF
C3608 VBIAS.n386 GND 0.01fF
C3609 VBIAS.n387 GND 0.01fF
C3610 VBIAS.n388 GND 0.01fF
C3611 VBIAS.n389 GND 0.01fF
C3612 VBIAS.n390 GND 0.05fF
C3613 VBIAS.n391 GND 0.46fF
C3614 VBIAS.n392 GND 0.03fF
C3615 VBIAS.n393 GND 0.03fF
C3616 VBIAS.n394 GND 0.01fF
C3617 VBIAS.n395 GND 0.04fF
C3618 VBIAS.n396 GND 0.04fF
C3619 VBIAS.n397 GND 0.01fF
C3620 VBIAS.n398 GND 0.04fF
C3621 VBIAS.n399 GND 0.03fF
C3622 VBIAS.n400 GND 0.01fF
C3623 VBIAS.n401 GND 0.17fF
C3624 VBIAS.n402 GND 0.01fF
C3625 VBIAS.n403 GND 0.01fF
C3626 VBIAS.n404 GND 0.01fF
C3627 VBIAS.n405 GND 0.03fF
C3628 VBIAS.n406 GND 0.03fF
C3629 VBIAS.n407 GND 0.01fF
C3630 VBIAS.n408 GND 0.04fF
C3631 VBIAS.n409 GND 0.01fF
C3632 VBIAS.n410 GND 0.01fF
C3633 VBIAS.n411 GND 0.01fF
C3634 VBIAS.n412 GND 0.00fF
C3635 VBIAS.n413 GND 0.01fF
C3636 VBIAS.n414 GND 0.00fF
C3637 VBIAS.n415 GND 0.12fF
C3638 VBIAS.n416 GND 0.01fF
C3639 VBIAS.n417 GND 0.01fF
C3640 VBIAS.n418 GND 0.02fF
C3641 VBIAS.n419 GND 0.00fF
C3642 VBIAS.n420 GND 0.01fF
C3643 VBIAS.n421 GND 0.00fF
C3644 VBIAS.n422 GND 0.01fF
C3645 VBIAS.n423 GND 0.01fF
C3646 VBIAS.n424 GND 0.01fF
C3647 VBIAS.n425 GND 0.01fF
C3648 VBIAS.n426 GND 0.01fF
C3649 VBIAS.n427 GND 0.01fF
C3650 VBIAS.n428 GND 0.03fF
C3651 VBIAS.n429 GND 0.12fF
C3652 VBIAS.n430 GND 0.02fF
C3653 VBIAS.n431 GND 0.04fF
C3654 VBIAS.n432 GND 0.01fF
C3655 VBIAS.n433 GND 0.01fF
C3656 VBIAS.n434 GND 0.01fF
C3657 VBIAS.n435 GND 0.01fF
C3658 VBIAS.n436 GND 0.03fF
C3659 VBIAS.n437 GND 0.02fF
C3660 VBIAS.n438 GND 0.01fF
C3661 VBIAS.n439 GND 0.01fF
C3662 VBIAS.n440 GND 0.00fF
C3663 VBIAS.n441 GND 0.00fF
C3664 VBIAS.n442 GND 0.01fF
C3665 VBIAS.n443 GND 0.01fF
C3666 VBIAS.n444 GND 0.01fF
C3667 VBIAS.n445 GND 0.00fF
C3668 VBIAS.n446 GND 0.01fF
C3669 VBIAS.n447 GND 0.04fF
C3670 VBIAS.n448 GND 0.00fF
C3671 VBIAS.n449 GND 0.01fF
C3672 VBIAS.n450 GND 0.01fF
C3673 VBIAS.n451 GND 0.01fF
C3674 VBIAS.n452 GND 0.01fF
C3675 VBIAS.n453 GND 0.00fF
C3676 VBIAS.n454 GND 0.00fF
C3677 VBIAS.n455 GND 0.00fF
C3678 VBIAS.n456 GND 0.01fF
C3679 VBIAS.n457 GND 0.01fF
C3680 VBIAS.n458 GND 0.02fF
C3681 VBIAS.n459 GND 0.02fF
C3682 VBIAS.n460 GND 0.01fF
C3683 VBIAS.n461 GND 0.03fF
C3684 VBIAS.n462 GND 0.12fF
C3685 VBIAS.n463 GND 0.01fF
C3686 VBIAS.n464 GND 0.02fF
C3687 VBIAS.n465 GND 0.04fF
C3688 VBIAS.n466 GND 0.01fF
C3689 VBIAS.n467 GND 0.01fF
C3690 VBIAS.n468 GND 0.00fF
C3691 VBIAS.n469 GND 0.01fF
C3692 VBIAS.n470 GND 0.00fF
C3693 VBIAS.n471 GND 0.12fF
C3694 VBIAS.n472 GND 0.01fF
C3695 VBIAS.n473 GND 0.01fF
C3696 VBIAS.n474 GND 0.02fF
C3697 VBIAS.n475 GND 0.00fF
C3698 VBIAS.n476 GND 0.01fF
C3699 VBIAS.n477 GND 0.00fF
C3700 VBIAS.n478 GND 0.01fF
C3701 VBIAS.n479 GND 0.01fF
C3702 VBIAS.n480 GND 0.01fF
C3703 VBIAS.n481 GND 0.01fF
C3704 VBIAS.n482 GND 0.01fF
C3705 VBIAS.n483 GND 0.01fF
C3706 VBIAS.n484 GND 0.01fF
C3707 VBIAS.n485 GND 0.01fF
C3708 VBIAS.n486 GND 0.05fF
C3709 VBIAS.n487 GND 0.17fF
C3710 VBIAS.n488 GND 0.03fF
C3711 VBIAS.n489 GND 0.03fF
C3712 VBIAS.n490 GND 0.01fF
C3713 VBIAS.n491 GND 0.04fF
C3714 VBIAS.n492 GND 0.04fF
C3715 VBIAS.n493 GND 0.01fF
C3716 VBIAS.n494 GND 0.04fF
C3717 VBIAS.n495 GND 0.03fF
C3718 VBIAS.n496 GND 0.01fF
C3719 VBIAS.n497 GND 0.51fF
C3720 VBIAS.n498 GND 0.00fF
C3721 VBIAS.n499 GND 0.03fF
C3722 VBIAS.t9 GND 0.20fF $ **FLOATING
C3723 VBIAS.n500 GND 0.12fF
C3724 VBIAS.n501 GND 0.01fF
C3725 VBIAS.n502 GND 0.02fF
C3726 VBIAS.n503 GND 0.05fF
C3727 VBIAS.n504 GND 0.01fF
C3728 VBIAS.n505 GND 0.01fF
C3729 VBIAS.n506 GND 0.01fF
C3730 VBIAS.n507 GND 0.02fF
C3731 VBIAS.n508 GND 0.01fF
C3732 VBIAS.n509 GND 0.02fF
C3733 VBIAS.n510 GND 0.00fF
C3734 VBIAS.n511 GND 0.01fF
C3735 VBIAS.n512 GND 0.00fF
C3736 VBIAS.n513 GND 0.00fF
C3737 VBIAS.n514 GND 0.00fF
C3738 VBIAS.t31 GND 0.20fF $ **FLOATING
C3739 VBIAS.n515 GND 0.12fF
C3740 VBIAS.n516 GND 0.01fF
C3741 VBIAS.n517 GND 0.01fF
C3742 VBIAS.n518 GND 0.02fF
C3743 VBIAS.n519 GND 0.00fF
C3744 VBIAS.n520 GND 0.01fF
C3745 VBIAS.n521 GND 0.01fF
C3746 VBIAS.n522 GND 0.00fF
C3747 VBIAS.n523 GND 0.02fF
C3748 VBIAS.n524 GND 0.01fF
C3749 VBIAS.n525 GND 0.03fF
C3750 VBIAS.n526 GND 0.03fF
C3751 VBIAS.n527 GND 0.01fF
C3752 VBIAS.n528 GND 0.00fF
C3753 VBIAS.n529 GND 0.04fF
C3754 VBIAS.n530 GND 0.01fF
C3755 VBIAS.n531 GND 0.01fF
C3756 VBIAS.n532 GND 0.01fF
C3757 VBIAS.n533 GND 0.01fF
C3758 VBIAS.n534 GND 0.03fF
C3759 VBIAS.n535 GND 0.02fF
C3760 VBIAS.n536 GND 0.01fF
C3761 VBIAS.n537 GND 0.01fF
C3762 VBIAS.n538 GND 0.00fF
C3763 VBIAS.n539 GND 0.01fF
C3764 VBIAS.n540 GND 0.00fF
C3765 VBIAS.n541 GND 0.01fF
C3766 VBIAS.n542 GND 0.01fF
C3767 VBIAS.n543 GND 0.02fF
C3768 VBIAS.n544 GND 0.01fF
C3769 VBIAS.n545 GND 0.00fF
C3770 VBIAS.n546 GND 0.04fF
C3771 VBIAS.n547 GND 0.00fF
C3772 VBIAS.n548 GND 0.01fF
C3773 VBIAS.n549 GND 0.01fF
C3774 VBIAS.n550 GND 0.02fF
C3775 VBIAS.n551 GND 0.01fF
C3776 VBIAS.n552 GND 0.00fF
C3777 VBIAS.n553 GND 0.01fF
C3778 VBIAS.n554 GND 0.00fF
C3779 VBIAS.n555 GND 0.01fF
C3780 VBIAS.n556 GND 0.01fF
C3781 VBIAS.n557 GND 0.02fF
C3782 VBIAS.n558 GND 0.02fF
C3783 VBIAS.n559 GND 0.01fF
C3784 VBIAS.n560 GND 0.01fF
C3785 VBIAS.n561 GND 0.01fF
C3786 VBIAS.t17 GND 0.20fF $ **FLOATING
C3787 VBIAS.n562 GND 0.03fF
C3788 VBIAS.n563 GND 0.12fF
C3789 VBIAS.n564 GND 0.02fF
C3790 VBIAS.n565 GND 0.06fF
C3791 VBIAS.n566 GND 0.01fF
C3792 VBIAS.n567 GND 0.00fF
C3793 VBIAS.n568 GND 0.02fF
C3794 VBIAS.n569 GND 0.00fF
C3795 VBIAS.t32 GND 0.20fF $ **FLOATING
C3796 VBIAS.n570 GND 0.12fF
C3797 VBIAS.n571 GND 0.01fF
C3798 VBIAS.n572 GND 0.01fF
C3799 VBIAS.n573 GND 0.02fF
C3800 VBIAS.n574 GND 0.00fF
C3801 VBIAS.n575 GND 0.01fF
C3802 VBIAS.n576 GND 0.00fF
C3803 VBIAS.n577 GND 0.00fF
C3804 VBIAS.n578 GND 0.00fF
C3805 VBIAS.n579 GND 0.01fF
C3806 VBIAS.n580 GND 0.01fF
C3807 VBIAS.n581 GND 0.01fF
C3808 VBIAS.n582 GND 0.01fF
C3809 VBIAS.n583 GND 0.01fF
C3810 VBIAS.n584 GND 0.01fF
C3811 VBIAS.n585 GND 0.01fF
C3812 VBIAS.n586 GND 0.01fF
C3813 VBIAS.n587 GND 0.05fF
C3814 VBIAS.n588 GND 0.10fF
C3815 VBIAS.n589 GND 0.01fF
C3816 VBIAS.n590 GND 0.04fF
C3817 VBIAS.n591 GND 0.04fF
C3818 VBIAS.n592 GND 0.01fF
C3819 VBIAS.n593 GND 0.04fF
C3820 VBIAS.n594 GND 0.03fF
C3821 VBIAS.n595 GND 0.01fF
C3822 VBIAS.n596 GND 0.17fF
C3823 VBIAS.n597 GND 0.01fF
C3824 VBIAS.n598 GND 0.01fF
C3825 VBIAS.t10 GND 0.20fF $ **FLOATING
C3826 VBIAS.n599 GND 0.03fF
C3827 VBIAS.n600 GND 0.12fF
C3828 VBIAS.n601 GND 0.02fF
C3829 VBIAS.n602 GND 0.06fF
C3830 VBIAS.n603 GND 0.01fF
C3831 VBIAS.n604 GND 0.01fF
C3832 VBIAS.n605 GND 0.01fF
C3833 VBIAS.t11 GND 0.20fF $ **FLOATING
C3834 VBIAS.n606 GND 0.03fF
C3835 VBIAS.n607 GND 0.12fF
C3836 VBIAS.n608 GND 0.02fF
C3837 VBIAS.n609 GND 0.05fF
C3838 VBIAS.n610 GND 0.01fF
C3839 VBIAS.n611 GND 0.01fF
C3840 VBIAS.n612 GND 0.01fF
C3841 VBIAS.n613 GND 0.02fF
C3842 VBIAS.n614 GND 0.01fF
C3843 VBIAS.n615 GND 0.02fF
C3844 VBIAS.n616 GND 0.00fF
C3845 VBIAS.n617 GND 0.01fF
C3846 VBIAS.n618 GND 0.00fF
C3847 VBIAS.n619 GND 0.00fF
C3848 VBIAS.n620 GND 0.00fF
C3849 VBIAS.t28 GND 0.20fF $ **FLOATING
C3850 VBIAS.n621 GND 0.12fF
C3851 VBIAS.n622 GND 0.01fF
C3852 VBIAS.n623 GND 0.01fF
C3853 VBIAS.n624 GND 0.02fF
C3854 VBIAS.n625 GND 0.00fF
C3855 VBIAS.n626 GND 0.01fF
C3856 VBIAS.n627 GND 0.01fF
C3857 VBIAS.n628 GND 0.00fF
C3858 VBIAS.n629 GND 0.02fF
C3859 VBIAS.n630 GND 0.01fF
C3860 VBIAS.n631 GND 0.02fF
C3861 VBIAS.n632 GND 0.02fF
C3862 VBIAS.n633 GND 0.01fF
C3863 VBIAS.n634 GND 0.01fF
C3864 VBIAS.n635 GND 0.00fF
C3865 VBIAS.n636 GND 0.00fF
C3866 VBIAS.n637 GND 0.01fF
C3867 VBIAS.n638 GND 0.03fF
C3868 VBIAS.n639 GND 0.03fF
C3869 VBIAS.n640 GND 0.01fF
C3870 VBIAS.n641 GND 0.00fF
C3871 VBIAS.n642 GND 0.04fF
C3872 VBIAS.n643 GND 0.01fF
C3873 VBIAS.n644 GND 0.01fF
C3874 VBIAS.n645 GND 0.01fF
C3875 VBIAS.n646 GND 0.01fF
C3876 VBIAS.n647 GND 0.03fF
C3877 VBIAS.n648 GND 0.02fF
C3878 VBIAS.n649 GND 0.01fF
C3879 VBIAS.n650 GND 0.01fF
C3880 VBIAS.n651 GND 0.00fF
C3881 VBIAS.n652 GND 0.01fF
C3882 VBIAS.n653 GND 0.00fF
C3883 VBIAS.n654 GND 0.01fF
C3884 VBIAS.n655 GND 0.02fF
C3885 VBIAS.n656 GND 0.01fF
C3886 VBIAS.n657 GND 0.04fF
C3887 VBIAS.n658 GND 0.00fF
C3888 VBIAS.n659 GND 0.00fF
C3889 VBIAS.n660 GND 0.01fF
C3890 VBIAS.n661 GND 0.02fF
C3891 VBIAS.n662 GND 0.01fF
C3892 VBIAS.n663 GND 0.00fF
C3893 VBIAS.n664 GND 0.01fF
C3894 VBIAS.n665 GND 0.01fF
C3895 VBIAS.n666 GND 0.00fF
C3896 VBIAS.n667 GND 0.02fF
C3897 VBIAS.n668 GND 0.00fF
C3898 VBIAS.t35 GND 0.20fF $ **FLOATING
C3899 VBIAS.n669 GND 0.12fF
C3900 VBIAS.n670 GND 0.01fF
C3901 VBIAS.n671 GND 0.01fF
C3902 VBIAS.n672 GND 0.02fF
C3903 VBIAS.n673 GND 0.00fF
C3904 VBIAS.n674 GND 0.01fF
C3905 VBIAS.n675 GND 0.00fF
C3906 VBIAS.n676 GND 0.00fF
C3907 VBIAS.n677 GND 0.00fF
C3908 VBIAS.n678 GND 0.01fF
C3909 VBIAS.n679 GND 0.01fF
C3910 VBIAS.n680 GND 0.01fF
C3911 VBIAS.n681 GND 0.01fF
C3912 VBIAS.n682 GND 0.01fF
C3913 VBIAS.n683 GND 0.01fF
C3914 VBIAS.n684 GND 0.01fF
C3915 VBIAS.n685 GND 0.01fF
C3916 VBIAS.n686 GND 0.05fF
C3917 VBIAS.n687 GND 0.17fF
C3918 VBIAS.n688 GND 0.03fF
C3919 VBIAS.n689 GND 0.03fF
C3920 VBIAS.n690 GND 0.01fF
C3921 VBIAS.n691 GND 0.04fF
C3922 VBIAS.n692 GND 0.04fF
C3923 VBIAS.n693 GND 0.01fF
C3924 VBIAS.n694 GND 0.04fF
C3925 VBIAS.n695 GND 0.03fF
C3926 VBIAS.n696 GND 0.01fF
C3927 VBIAS.n697 GND 0.46fF
C3928 VBIAS.n698 GND 0.01fF
C3929 VBIAS.n699 GND 0.01fF
C3930 VBIAS.t15 GND 0.20fF $ **FLOATING
C3931 VBIAS.n700 GND 0.03fF
C3932 VBIAS.n701 GND 0.12fF
C3933 VBIAS.n702 GND 0.02fF
C3934 VBIAS.n703 GND 0.06fF
C3935 VBIAS.n704 GND 0.01fF
C3936 VBIAS.n705 GND 0.01fF
C3937 VBIAS.n706 GND 0.01fF
C3938 VBIAS.t18 GND 0.20fF $ **FLOATING
C3939 VBIAS.n707 GND 0.03fF
C3940 VBIAS.n708 GND 0.12fF
C3941 VBIAS.n709 GND 0.02fF
C3942 VBIAS.n710 GND 0.05fF
C3943 VBIAS.n711 GND 0.01fF
C3944 VBIAS.n712 GND 0.01fF
C3945 VBIAS.n713 GND 0.01fF
C3946 VBIAS.n714 GND 0.02fF
C3947 VBIAS.n715 GND 0.01fF
C3948 VBIAS.n716 GND 0.02fF
C3949 VBIAS.n717 GND 0.00fF
C3950 VBIAS.n718 GND 0.01fF
C3951 VBIAS.n719 GND 0.00fF
C3952 VBIAS.n720 GND 0.00fF
C3953 VBIAS.n721 GND 0.00fF
C3954 VBIAS.t19 GND 0.20fF $ **FLOATING
C3955 VBIAS.n722 GND 0.12fF
C3956 VBIAS.n723 GND 0.01fF
C3957 VBIAS.n724 GND 0.01fF
C3958 VBIAS.n725 GND 0.02fF
C3959 VBIAS.n726 GND 0.00fF
C3960 VBIAS.n727 GND 0.01fF
C3961 VBIAS.n728 GND 0.01fF
C3962 VBIAS.n729 GND 0.00fF
C3963 VBIAS.n730 GND 0.02fF
C3964 VBIAS.n731 GND 0.01fF
C3965 VBIAS.n732 GND 0.02fF
C3966 VBIAS.n733 GND 0.02fF
C3967 VBIAS.n734 GND 0.01fF
C3968 VBIAS.n735 GND 0.01fF
C3969 VBIAS.n736 GND 0.00fF
C3970 VBIAS.n737 GND 0.00fF
C3971 VBIAS.n738 GND 0.01fF
C3972 VBIAS.n739 GND 0.03fF
C3973 VBIAS.n740 GND 0.03fF
C3974 VBIAS.n741 GND 0.01fF
C3975 VBIAS.n742 GND 0.00fF
C3976 VBIAS.n743 GND 0.04fF
C3977 VBIAS.n744 GND 0.01fF
C3978 VBIAS.n745 GND 0.01fF
C3979 VBIAS.n746 GND 0.01fF
C3980 VBIAS.n747 GND 0.01fF
C3981 VBIAS.n748 GND 0.03fF
C3982 VBIAS.n749 GND 0.02fF
C3983 VBIAS.n750 GND 0.01fF
C3984 VBIAS.n751 GND 0.01fF
C3985 VBIAS.n752 GND 0.00fF
C3986 VBIAS.n753 GND 0.01fF
C3987 VBIAS.n754 GND 0.00fF
C3988 VBIAS.n755 GND 0.01fF
C3989 VBIAS.n756 GND 0.02fF
C3990 VBIAS.n757 GND 0.01fF
C3991 VBIAS.n758 GND 0.04fF
C3992 VBIAS.n759 GND 0.00fF
C3993 VBIAS.n760 GND 0.00fF
C3994 VBIAS.n761 GND 0.01fF
C3995 VBIAS.n762 GND 0.02fF
C3996 VBIAS.n763 GND 0.01fF
C3997 VBIAS.n764 GND 0.00fF
C3998 VBIAS.n765 GND 0.01fF
C3999 VBIAS.n766 GND 0.01fF
C4000 VBIAS.n767 GND 0.00fF
C4001 VBIAS.n768 GND 0.02fF
C4002 VBIAS.n769 GND 0.00fF
C4003 VBIAS.t30 GND 0.20fF $ **FLOATING
C4004 VBIAS.n770 GND 0.12fF
C4005 VBIAS.n771 GND 0.01fF
C4006 VBIAS.n772 GND 0.01fF
C4007 VBIAS.n773 GND 0.02fF
C4008 VBIAS.n774 GND 0.00fF
C4009 VBIAS.n775 GND 0.01fF
C4010 VBIAS.n776 GND 0.00fF
C4011 VBIAS.n777 GND 0.00fF
C4012 VBIAS.n778 GND 0.00fF
C4013 VBIAS.n779 GND 0.01fF
C4014 VBIAS.n780 GND 0.01fF
C4015 VBIAS.n781 GND 0.01fF
C4016 VBIAS.n782 GND 0.01fF
C4017 VBIAS.n783 GND 0.01fF
C4018 VBIAS.n784 GND 0.01fF
C4019 VBIAS.n785 GND 0.01fF
C4020 VBIAS.n786 GND 0.01fF
C4021 VBIAS.n787 GND 0.05fF
C4022 VBIAS.n788 GND 0.46fF
C4023 VBIAS.n789 GND 0.03fF
C4024 VBIAS.n790 GND 0.03fF
C4025 VBIAS.n791 GND 0.01fF
C4026 VBIAS.n792 GND 0.04fF
C4027 VBIAS.n793 GND 0.04fF
C4028 VBIAS.n794 GND 0.01fF
C4029 VBIAS.n795 GND 0.04fF
C4030 VBIAS.n796 GND 0.03fF
C4031 VBIAS.n797 GND 0.01fF
C4032 VBIAS.n798 GND 0.17fF
C4033 VBIAS.n799 GND 0.01fF
C4034 VBIAS.n800 GND 0.01fF
C4035 VBIAS.t8 GND 0.20fF $ **FLOATING
C4036 VBIAS.n801 GND 0.03fF
C4037 VBIAS.n802 GND 0.12fF
C4038 VBIAS.n803 GND 0.02fF
C4039 VBIAS.n804 GND 0.06fF
C4040 VBIAS.n805 GND 0.01fF
C4041 VBIAS.n806 GND 0.01fF
C4042 VBIAS.n807 GND 0.01fF
C4043 VBIAS.t20 GND 0.20fF $ **FLOATING
C4044 VBIAS.n808 GND 0.03fF
C4045 VBIAS.n809 GND 0.12fF
C4046 VBIAS.n810 GND 0.02fF
C4047 VBIAS.n811 GND 0.05fF
C4048 VBIAS.n812 GND 0.01fF
C4049 VBIAS.n813 GND 0.01fF
C4050 VBIAS.n814 GND 0.01fF
C4051 VBIAS.n815 GND 0.02fF
C4052 VBIAS.n816 GND 0.01fF
C4053 VBIAS.n817 GND 0.02fF
C4054 VBIAS.n818 GND 0.00fF
C4055 VBIAS.n819 GND 0.01fF
C4056 VBIAS.n820 GND 0.00fF
C4057 VBIAS.n821 GND 0.00fF
C4058 VBIAS.n822 GND 0.00fF
C4059 VBIAS.t21 GND 0.20fF $ **FLOATING
C4060 VBIAS.n823 GND 0.12fF
C4061 VBIAS.n824 GND 0.01fF
C4062 VBIAS.n825 GND 0.01fF
C4063 VBIAS.n826 GND 0.02fF
C4064 VBIAS.n827 GND 0.00fF
C4065 VBIAS.n828 GND 0.01fF
C4066 VBIAS.n829 GND 0.01fF
C4067 VBIAS.n830 GND 0.00fF
C4068 VBIAS.n831 GND 0.02fF
C4069 VBIAS.n832 GND 0.01fF
C4070 VBIAS.n833 GND 0.02fF
C4071 VBIAS.n834 GND 0.02fF
C4072 VBIAS.n835 GND 0.01fF
C4073 VBIAS.n836 GND 0.01fF
C4074 VBIAS.n837 GND 0.00fF
C4075 VBIAS.n838 GND 0.00fF
C4076 VBIAS.n839 GND 0.01fF
C4077 VBIAS.n840 GND 0.03fF
C4078 VBIAS.n841 GND 0.03fF
C4079 VBIAS.n842 GND 0.01fF
C4080 VBIAS.n843 GND 0.00fF
C4081 VBIAS.n844 GND 0.04fF
C4082 VBIAS.n845 GND 0.01fF
C4083 VBIAS.n846 GND 0.01fF
C4084 VBIAS.n847 GND 0.01fF
C4085 VBIAS.n848 GND 0.01fF
C4086 VBIAS.n849 GND 0.03fF
C4087 VBIAS.n850 GND 0.02fF
C4088 VBIAS.n851 GND 0.01fF
C4089 VBIAS.n852 GND 0.01fF
C4090 VBIAS.n853 GND 0.00fF
C4091 VBIAS.n854 GND 0.01fF
C4092 VBIAS.n855 GND 0.00fF
C4093 VBIAS.n856 GND 0.01fF
C4094 VBIAS.n857 GND 0.02fF
C4095 VBIAS.n858 GND 0.01fF
C4096 VBIAS.n859 GND 0.04fF
C4097 VBIAS.n860 GND 0.00fF
C4098 VBIAS.n861 GND 0.00fF
C4099 VBIAS.n862 GND 0.01fF
C4100 VBIAS.n863 GND 0.02fF
C4101 VBIAS.n864 GND 0.01fF
C4102 VBIAS.n865 GND 0.00fF
C4103 VBIAS.n866 GND 0.01fF
C4104 VBIAS.n867 GND 0.01fF
C4105 VBIAS.n868 GND 0.00fF
C4106 VBIAS.n869 GND 0.02fF
C4107 VBIAS.n870 GND 0.00fF
C4108 VBIAS.t33 GND 0.20fF $ **FLOATING
C4109 VBIAS.n871 GND 0.12fF
C4110 VBIAS.n872 GND 0.01fF
C4111 VBIAS.n873 GND 0.01fF
C4112 VBIAS.n874 GND 0.02fF
C4113 VBIAS.n875 GND 0.00fF
C4114 VBIAS.n876 GND 0.01fF
C4115 VBIAS.n877 GND 0.00fF
C4116 VBIAS.n878 GND 0.00fF
C4117 VBIAS.n879 GND 0.00fF
C4118 VBIAS.n880 GND 0.01fF
C4119 VBIAS.n881 GND 0.01fF
C4120 VBIAS.n882 GND 0.01fF
C4121 VBIAS.n883 GND 0.01fF
C4122 VBIAS.n884 GND 0.01fF
C4123 VBIAS.n885 GND 0.01fF
C4124 VBIAS.n886 GND 0.01fF
C4125 VBIAS.n887 GND 0.01fF
C4126 VBIAS.n888 GND 0.05fF
C4127 VBIAS.n889 GND 0.17fF
C4128 VBIAS.n890 GND 0.03fF
C4129 VBIAS.n891 GND 0.03fF
C4130 VBIAS.n892 GND 0.01fF
C4131 VBIAS.n893 GND 0.04fF
C4132 VBIAS.n894 GND 0.04fF
C4133 VBIAS.n895 GND 0.01fF
C4134 VBIAS.n896 GND 0.04fF
C4135 VBIAS.n897 GND 0.03fF
C4136 VBIAS.n898 GND 0.01fF
C4137 VBIAS.n899 GND 0.26fF
C4138 VBIAS.n900 GND 0.91fF
C4139 VBIAS.n901 GND 0.01fF
C4140 VBIAS.n902 GND 0.01fF
C4141 VBIAS.n903 GND 0.03fF
C4142 VBIAS.n904 GND 0.12fF
C4143 VBIAS.n905 GND 0.02fF
C4144 VBIAS.n906 GND 0.05fF
C4145 VBIAS.n907 GND 0.01fF
C4146 VBIAS.n908 GND 0.03fF
C4147 VBIAS.n909 GND 0.12fF
C4148 VBIAS.n910 GND 0.02fF
C4149 VBIAS.n911 GND 0.05fF
C4150 VBIAS.n912 GND 0.01fF
C4151 VBIAS.n913 GND 0.01fF
C4152 VBIAS.n914 GND 0.01fF
C4153 VBIAS.n915 GND 0.02fF
C4154 VBIAS.n916 GND 0.01fF
C4155 VBIAS.n917 GND 0.02fF
C4156 VBIAS.n918 GND 0.00fF
C4157 VBIAS.n919 GND 0.01fF
C4158 VBIAS.n920 GND 0.00fF
C4159 VBIAS.n921 GND 0.00fF
C4160 VBIAS.n922 GND 0.00fF
C4161 VBIAS.n923 GND 0.12fF
C4162 VBIAS.n924 GND 0.01fF
C4163 VBIAS.n925 GND 0.01fF
C4164 VBIAS.n926 GND 0.02fF
C4165 VBIAS.n927 GND 0.00fF
C4166 VBIAS.n928 GND 0.01fF
C4167 VBIAS.n929 GND 0.01fF
C4168 VBIAS.n930 GND 0.00fF
C4169 VBIAS.n931 GND 0.02fF
C4170 VBIAS.n932 GND 0.01fF
C4171 VBIAS.n933 GND 0.01fF
C4172 VBIAS.n934 GND 0.02fF
C4173 VBIAS.n935 GND 0.02fF
C4174 VBIAS.n936 GND 0.01fF
C4175 VBIAS.n937 GND 0.01fF
C4176 VBIAS.n938 GND 0.00fF
C4177 VBIAS.n939 GND 0.00fF
C4178 VBIAS.n940 GND 0.01fF
C4179 VBIAS.n941 GND 0.03fF
C4180 VBIAS.n942 GND 0.03fF
C4181 VBIAS.n943 GND 0.01fF
C4182 VBIAS.n944 GND 0.04fF
C4183 VBIAS.n945 GND 0.01fF
C4184 VBIAS.n946 GND 0.01fF
C4185 VBIAS.n947 GND 0.01fF
C4186 VBIAS.n948 GND 0.01fF
C4187 VBIAS.n949 GND 0.03fF
C4188 VBIAS.n950 GND 0.02fF
C4189 VBIAS.n951 GND 0.01fF
C4190 VBIAS.n952 GND 0.01fF
C4191 VBIAS.n953 GND 0.00fF
C4192 VBIAS.n954 GND 0.00fF
C4193 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE GND 0.01fF
C4194 VBIAS.n955 GND 0.01fF
C4195 VBIAS.n956 GND 0.01fF
C4196 VBIAS.n957 GND 0.02fF
C4197 VBIAS.n958 GND 0.01fF
C4198 VBIAS.n959 GND 0.00fF
C4199 VBIAS.n960 GND 0.04fF
C4200 VBIAS.n961 GND 0.00fF
C4201 VBIAS.n962 GND 0.01fF
C4202 VBIAS.n963 GND 0.01fF
C4203 VBIAS.n964 GND 0.02fF
C4204 VBIAS.n965 GND 0.01fF
C4205 VBIAS.n966 GND 0.00fF
C4206 VBIAS.n967 GND 0.01fF
C4207 VBIAS.n968 GND 0.01fF
C4208 VBIAS.n969 GND 0.00fF
C4209 VBIAS.n970 GND 0.02fF
C4210 VBIAS.n971 GND 0.00fF
C4211 VBIAS.n972 GND 0.12fF
C4212 VBIAS.n973 GND 0.01fF
C4213 VBIAS.n974 GND 0.01fF
C4214 VBIAS.n975 GND 0.02fF
C4215 VBIAS.n976 GND 0.00fF
C4216 VBIAS.n977 GND 0.01fF
C4217 VBIAS.n978 GND 0.00fF
C4218 VBIAS.n979 GND 0.00fF
C4219 VBIAS.n980 GND 0.00fF
C4220 VBIAS.n981 GND 0.01fF
C4221 VBIAS.n982 GND 0.01fF
C4222 VBIAS.n983 GND 0.01fF
C4223 VBIAS.n984 GND 0.01fF
C4224 VBIAS.n985 GND 0.01fF
C4225 VBIAS.n986 GND 0.01fF
C4226 VBIAS.n987 GND 0.01fF
C4227 VBIAS.n988 GND 0.01fF
C4228 VBIAS.n989 GND 0.05fF
C4229 VBIAS.n990 GND 0.10fF
C4230 VBIAS.n991 GND 0.01fF
C4231 VBIAS.n992 GND 0.04fF
C4232 VBIAS.n993 GND 0.04fF
C4233 VBIAS.n994 GND 0.01fF
C4234 VBIAS.n995 GND 0.04fF
C4235 VBIAS.n996 GND 0.03fF
C4236 VBIAS.n997 GND 0.01fF
C4237 VBIAS.n998 GND 0.17fF
C4238 VBIAS.n999 GND 0.01fF
C4239 VBIAS.n1000 GND 0.01fF
C4240 VBIAS.n1001 GND 0.03fF
C4241 VBIAS.n1002 GND 0.12fF
C4242 VBIAS.n1003 GND 0.02fF
C4243 VBIAS.n1004 GND 0.05fF
C4244 VBIAS.n1005 GND 0.03fF
C4245 VBIAS.n1006 GND 0.12fF
C4246 VBIAS.n1007 GND 0.01fF
C4247 VBIAS.n1008 GND 0.02fF
C4248 VBIAS.n1009 GND 0.05fF
C4249 VBIAS.n1010 GND 0.01fF
C4250 VBIAS.n1011 GND 0.01fF
C4251 VBIAS.n1012 GND 0.01fF
C4252 VBIAS.n1013 GND 0.02fF
C4253 VBIAS.n1014 GND 0.01fF
C4254 VBIAS.n1015 GND 0.02fF
C4255 VBIAS.n1016 GND 0.00fF
C4256 VBIAS.n1017 GND 0.01fF
C4257 VBIAS.n1018 GND 0.00fF
C4258 VBIAS.n1019 GND 0.00fF
C4259 VBIAS.n1020 GND 0.00fF
C4260 VBIAS.n1021 GND 0.12fF
C4261 VBIAS.n1022 GND 0.01fF
C4262 VBIAS.n1023 GND 0.01fF
C4263 VBIAS.n1024 GND 0.02fF
C4264 VBIAS.n1025 GND 0.00fF
C4265 VBIAS.n1026 GND 0.01fF
C4266 VBIAS.n1027 GND 0.01fF
C4267 VBIAS.n1028 GND 0.00fF
C4268 VBIAS.n1029 GND 0.02fF
C4269 VBIAS.n1030 GND 0.01fF
C4270 VBIAS.n1031 GND 0.01fF
C4271 VBIAS.n1032 GND 0.02fF
C4272 VBIAS.n1033 GND 0.02fF
C4273 VBIAS.n1034 GND 0.01fF
C4274 VBIAS.n1035 GND 0.01fF
C4275 VBIAS.n1036 GND 0.00fF
C4276 VBIAS.n1037 GND 0.00fF
C4277 VBIAS.n1038 GND 0.01fF
C4278 VBIAS.n1039 GND 0.03fF
C4279 VBIAS.n1040 GND 0.03fF
C4280 VBIAS.n1041 GND 0.01fF
C4281 VBIAS.n1042 GND 0.04fF
C4282 VBIAS.n1043 GND 0.01fF
C4283 VBIAS.n1044 GND 0.01fF
C4284 VBIAS.n1045 GND 0.01fF
C4285 VBIAS.n1046 GND 0.01fF
C4286 VBIAS.n1047 GND 0.03fF
C4287 VBIAS.n1048 GND 0.02fF
C4288 VBIAS.n1049 GND 0.01fF
C4289 VBIAS.n1050 GND 0.01fF
C4290 VBIAS.n1051 GND 0.00fF
C4291 VBIAS.n1052 GND 0.00fF
C4292 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE GND 0.01fF
C4293 VBIAS.n1053 GND 0.01fF
C4294 VBIAS.n1054 GND 0.01fF
C4295 VBIAS.n1055 GND 0.02fF
C4296 VBIAS.n1056 GND 0.01fF
C4297 VBIAS.n1057 GND 0.00fF
C4298 VBIAS.n1058 GND 0.04fF
C4299 VBIAS.n1059 GND 0.00fF
C4300 VBIAS.n1060 GND 0.01fF
C4301 VBIAS.n1061 GND 0.01fF
C4302 VBIAS.n1062 GND 0.02fF
C4303 VBIAS.n1063 GND 0.01fF
C4304 VBIAS.n1064 GND 0.00fF
C4305 VBIAS.n1065 GND 0.01fF
C4306 VBIAS.n1066 GND 0.01fF
C4307 VBIAS.n1067 GND 0.00fF
C4308 VBIAS.n1068 GND 0.02fF
C4309 VBIAS.n1069 GND 0.00fF
C4310 VBIAS.n1070 GND 0.12fF
C4311 VBIAS.n1071 GND 0.01fF
C4312 VBIAS.n1072 GND 0.01fF
C4313 VBIAS.n1073 GND 0.02fF
C4314 VBIAS.n1074 GND 0.00fF
C4315 VBIAS.n1075 GND 0.01fF
C4316 VBIAS.n1076 GND 0.00fF
C4317 VBIAS.n1077 GND 0.00fF
C4318 VBIAS.n1078 GND 0.00fF
C4319 VBIAS.n1079 GND 0.01fF
C4320 VBIAS.n1080 GND 0.01fF
C4321 VBIAS.n1081 GND 0.01fF
C4322 VBIAS.n1082 GND 0.01fF
C4323 VBIAS.n1083 GND 0.01fF
C4324 VBIAS.n1084 GND 0.01fF
C4325 VBIAS.n1085 GND 0.01fF
C4326 VBIAS.n1086 GND 0.01fF
C4327 VBIAS.n1087 GND 0.05fF
C4328 VBIAS.n1088 GND 0.16fF
C4329 VBIAS.n1089 GND 0.03fF
C4330 VBIAS.n1090 GND 0.03fF
C4331 VBIAS.n1091 GND 0.01fF
C4332 VBIAS.n1092 GND 0.04fF
C4333 VBIAS.n1093 GND 0.04fF
C4334 VBIAS.n1094 GND 0.01fF
C4335 VBIAS.n1095 GND 0.04fF
C4336 VBIAS.n1096 GND 0.03fF
C4337 VBIAS.n1097 GND 0.01fF
C4338 VBIAS.n1098 GND 0.17fF
C4339 VBIAS.n1099 GND 0.01fF
C4340 VBIAS.n1100 GND 0.03fF
C4341 VBIAS.n1101 GND 0.12fF
C4342 VBIAS.n1102 GND 0.01fF
C4343 VBIAS.n1103 GND 0.02fF
C4344 VBIAS.n1104 GND 0.05fF
C4345 VBIAS.n1105 GND 0.01fF
C4346 VBIAS.n1106 GND 0.03fF
C4347 VBIAS.n1107 GND 0.12fF
C4348 VBIAS.n1108 GND 0.02fF
C4349 VBIAS.n1109 GND 0.05fF
C4350 VBIAS.n1110 GND 0.01fF
C4351 VBIAS.n1111 GND 0.01fF
C4352 VBIAS.n1112 GND 0.01fF
C4353 VBIAS.n1113 GND 0.02fF
C4354 VBIAS.n1114 GND 0.01fF
C4355 VBIAS.n1115 GND 0.02fF
C4356 VBIAS.n1116 GND 0.00fF
C4357 VBIAS.n1117 GND 0.01fF
C4358 VBIAS.n1118 GND 0.00fF
C4359 VBIAS.n1119 GND 0.00fF
C4360 VBIAS.n1120 GND 0.00fF
C4361 VBIAS.n1121 GND 0.12fF
C4362 VBIAS.n1122 GND 0.01fF
C4363 VBIAS.n1123 GND 0.01fF
C4364 VBIAS.n1124 GND 0.02fF
C4365 VBIAS.n1125 GND 0.00fF
C4366 VBIAS.n1126 GND 0.01fF
C4367 VBIAS.n1127 GND 0.01fF
C4368 VBIAS.n1128 GND 0.00fF
C4369 VBIAS.n1129 GND 0.02fF
C4370 VBIAS.n1130 GND 0.01fF
C4371 VBIAS.n1131 GND 0.01fF
C4372 VBIAS.n1132 GND 0.02fF
C4373 VBIAS.n1133 GND 0.02fF
C4374 VBIAS.n1134 GND 0.01fF
C4375 VBIAS.n1135 GND 0.01fF
C4376 VBIAS.n1136 GND 0.00fF
C4377 VBIAS.n1137 GND 0.00fF
C4378 VBIAS.n1138 GND 0.01fF
C4379 VBIAS.n1139 GND 0.03fF
C4380 VBIAS.n1140 GND 0.03fF
C4381 VBIAS.n1141 GND 0.01fF
C4382 VBIAS.n1142 GND 0.04fF
C4383 VBIAS.n1143 GND 0.01fF
C4384 VBIAS.n1144 GND 0.01fF
C4385 VBIAS.n1145 GND 0.01fF
C4386 VBIAS.n1146 GND 0.01fF
C4387 VBIAS.n1147 GND 0.03fF
C4388 VBIAS.n1148 GND 0.02fF
C4389 VBIAS.n1149 GND 0.01fF
C4390 VBIAS.n1150 GND 0.01fF
C4391 VBIAS.n1151 GND 0.00fF
C4392 VBIAS.n1152 GND 0.00fF
C4393 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE GND 0.01fF
C4394 VBIAS.n1153 GND 0.01fF
C4395 VBIAS.n1154 GND 0.01fF
C4396 VBIAS.n1155 GND 0.02fF
C4397 VBIAS.n1156 GND 0.01fF
C4398 VBIAS.n1157 GND 0.00fF
C4399 VBIAS.n1158 GND 0.04fF
C4400 VBIAS.n1159 GND 0.00fF
C4401 VBIAS.n1160 GND 0.01fF
C4402 VBIAS.n1161 GND 0.01fF
C4403 VBIAS.n1162 GND 0.02fF
C4404 VBIAS.n1163 GND 0.01fF
C4405 VBIAS.n1164 GND 0.00fF
C4406 VBIAS.n1165 GND 0.01fF
C4407 VBIAS.n1166 GND 0.01fF
C4408 VBIAS.n1167 GND 0.00fF
C4409 VBIAS.n1168 GND 0.02fF
C4410 VBIAS.n1169 GND 0.00fF
C4411 VBIAS.n1170 GND 0.12fF
C4412 VBIAS.n1171 GND 0.01fF
C4413 VBIAS.n1172 GND 0.01fF
C4414 VBIAS.n1173 GND 0.02fF
C4415 VBIAS.n1174 GND 0.00fF
C4416 VBIAS.n1175 GND 0.01fF
C4417 VBIAS.n1176 GND 0.00fF
C4418 VBIAS.n1177 GND 0.00fF
C4419 VBIAS.n1178 GND 0.00fF
C4420 VBIAS.n1179 GND 0.01fF
C4421 VBIAS.n1180 GND 0.01fF
C4422 VBIAS.n1181 GND 0.01fF
C4423 VBIAS.n1182 GND 0.01fF
C4424 VBIAS.n1183 GND 0.01fF
C4425 VBIAS.n1184 GND 0.01fF
C4426 VBIAS.n1185 GND 0.01fF
C4427 VBIAS.n1186 GND 0.01fF
C4428 VBIAS.n1187 GND 0.05fF
C4429 VBIAS.n1188 GND 0.16fF
C4430 VBIAS.n1189 GND 0.03fF
C4431 VBIAS.n1190 GND 0.03fF
C4432 VBIAS.n1191 GND 0.01fF
C4433 VBIAS.n1192 GND 0.04fF
C4434 VBIAS.n1193 GND 0.04fF
C4435 VBIAS.n1194 GND 0.01fF
C4436 VBIAS.n1195 GND 0.04fF
C4437 VBIAS.n1196 GND 0.03fF
C4438 VBIAS.n1197 GND 0.01fF
C4439 VBIAS.n1198 GND 0.17fF
C4440 VBIAS.n1199 GND 0.01fF
C4441 VBIAS.n1200 GND 0.01fF
C4442 VBIAS.n1201 GND 0.03fF
C4443 VBIAS.n1202 GND 0.12fF
C4444 VBIAS.n1203 GND 0.02fF
C4445 VBIAS.n1204 GND 0.05fF
C4446 VBIAS.n1205 GND 0.03fF
C4447 VBIAS.n1206 GND 0.12fF
C4448 VBIAS.n1207 GND 0.01fF
C4449 VBIAS.n1208 GND 0.02fF
C4450 VBIAS.n1209 GND 0.05fF
C4451 VBIAS.n1210 GND 0.01fF
C4452 VBIAS.n1211 GND 0.01fF
C4453 VBIAS.n1212 GND 0.01fF
C4454 VBIAS.n1213 GND 0.02fF
C4455 VBIAS.n1214 GND 0.01fF
C4456 VBIAS.n1215 GND 0.02fF
C4457 VBIAS.n1216 GND 0.00fF
C4458 VBIAS.n1217 GND 0.01fF
C4459 VBIAS.n1218 GND 0.00fF
C4460 VBIAS.n1219 GND 0.00fF
C4461 VBIAS.n1220 GND 0.00fF
C4462 VBIAS.n1221 GND 0.12fF
C4463 VBIAS.n1222 GND 0.01fF
C4464 VBIAS.n1223 GND 0.01fF
C4465 VBIAS.n1224 GND 0.02fF
C4466 VBIAS.n1225 GND 0.00fF
C4467 VBIAS.n1226 GND 0.01fF
C4468 VBIAS.n1227 GND 0.01fF
C4469 VBIAS.n1228 GND 0.00fF
C4470 VBIAS.n1229 GND 0.02fF
C4471 VBIAS.n1230 GND 0.01fF
C4472 VBIAS.n1231 GND 0.01fF
C4473 VBIAS.n1232 GND 0.02fF
C4474 VBIAS.n1233 GND 0.02fF
C4475 VBIAS.n1234 GND 0.01fF
C4476 VBIAS.n1235 GND 0.01fF
C4477 VBIAS.n1236 GND 0.00fF
C4478 VBIAS.n1237 GND 0.00fF
C4479 VBIAS.n1238 GND 0.01fF
C4480 VBIAS.n1239 GND 0.03fF
C4481 VBIAS.n1240 GND 0.03fF
C4482 VBIAS.n1241 GND 0.01fF
C4483 VBIAS.n1242 GND 0.04fF
C4484 VBIAS.n1243 GND 0.01fF
C4485 VBIAS.n1244 GND 0.01fF
C4486 VBIAS.n1245 GND 0.01fF
C4487 VBIAS.n1246 GND 0.01fF
C4488 VBIAS.n1247 GND 0.03fF
C4489 VBIAS.n1248 GND 0.02fF
C4490 VBIAS.n1249 GND 0.01fF
C4491 VBIAS.n1250 GND 0.01fF
C4492 VBIAS.n1251 GND 0.00fF
C4493 VBIAS.n1252 GND 0.00fF
C4494 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE GND 0.01fF
C4495 VBIAS.n1253 GND 0.01fF
C4496 VBIAS.n1254 GND 0.01fF
C4497 VBIAS.n1255 GND 0.02fF
C4498 VBIAS.n1256 GND 0.01fF
C4499 VBIAS.n1257 GND 0.00fF
C4500 VBIAS.n1258 GND 0.04fF
C4501 VBIAS.n1259 GND 0.00fF
C4502 VBIAS.n1260 GND 0.01fF
C4503 VBIAS.n1261 GND 0.01fF
C4504 VBIAS.n1262 GND 0.02fF
C4505 VBIAS.n1263 GND 0.01fF
C4506 VBIAS.n1264 GND 0.00fF
C4507 VBIAS.n1265 GND 0.01fF
C4508 VBIAS.n1266 GND 0.01fF
C4509 VBIAS.n1267 GND 0.00fF
C4510 VBIAS.n1268 GND 0.02fF
C4511 VBIAS.n1269 GND 0.00fF
C4512 VBIAS.n1270 GND 0.12fF
C4513 VBIAS.n1271 GND 0.01fF
C4514 VBIAS.n1272 GND 0.01fF
C4515 VBIAS.n1273 GND 0.02fF
C4516 VBIAS.n1274 GND 0.00fF
C4517 VBIAS.n1275 GND 0.01fF
C4518 VBIAS.n1276 GND 0.00fF
C4519 VBIAS.n1277 GND 0.00fF
C4520 VBIAS.n1278 GND 0.00fF
C4521 VBIAS.n1279 GND 0.01fF
C4522 VBIAS.n1280 GND 0.01fF
C4523 VBIAS.n1281 GND 0.01fF
C4524 VBIAS.n1282 GND 0.01fF
C4525 VBIAS.n1283 GND 0.01fF
C4526 VBIAS.n1284 GND 0.01fF
C4527 VBIAS.n1285 GND 0.01fF
C4528 VBIAS.n1286 GND 0.01fF
C4529 VBIAS.n1287 GND 0.05fF
C4530 VBIAS.n1288 GND 0.16fF
C4531 VBIAS.n1289 GND 0.03fF
C4532 VBIAS.n1290 GND 0.03fF
C4533 VBIAS.n1291 GND 0.01fF
C4534 VBIAS.n1292 GND 0.04fF
C4535 VBIAS.n1293 GND 0.04fF
C4536 VBIAS.n1294 GND 0.01fF
C4537 VBIAS.n1295 GND 0.04fF
C4538 VBIAS.n1296 GND 0.03fF
C4539 VBIAS.n1297 GND 0.01fF
C4540 VBIAS.n1298 GND 0.17fF
C4541 VBIAS.n1299 GND 0.01fF
C4542 VBIAS.n1300 GND 0.01fF
C4543 VBIAS.n1301 GND 0.03fF
C4544 VBIAS.n1302 GND 0.12fF
C4545 VBIAS.n1303 GND 0.02fF
C4546 VBIAS.n1304 GND 0.05fF
C4547 VBIAS.n1305 GND 0.03fF
C4548 VBIAS.n1306 GND 0.12fF
C4549 VBIAS.n1307 GND 0.01fF
C4550 VBIAS.n1308 GND 0.02fF
C4551 VBIAS.n1309 GND 0.05fF
C4552 VBIAS.n1310 GND 0.01fF
C4553 VBIAS.n1311 GND 0.01fF
C4554 VBIAS.n1312 GND 0.01fF
C4555 VBIAS.n1313 GND 0.02fF
C4556 VBIAS.n1314 GND 0.01fF
C4557 VBIAS.n1315 GND 0.02fF
C4558 VBIAS.n1316 GND 0.00fF
C4559 VBIAS.n1317 GND 0.01fF
C4560 VBIAS.n1318 GND 0.00fF
C4561 VBIAS.n1319 GND 0.00fF
C4562 VBIAS.n1320 GND 0.00fF
C4563 VBIAS.n1321 GND 0.12fF
C4564 VBIAS.n1322 GND 0.01fF
C4565 VBIAS.n1323 GND 0.01fF
C4566 VBIAS.n1324 GND 0.02fF
C4567 VBIAS.n1325 GND 0.00fF
C4568 VBIAS.n1326 GND 0.01fF
C4569 VBIAS.n1327 GND 0.01fF
C4570 VBIAS.n1328 GND 0.00fF
C4571 VBIAS.n1329 GND 0.02fF
C4572 VBIAS.n1330 GND 0.01fF
C4573 VBIAS.n1331 GND 0.01fF
C4574 VBIAS.n1332 GND 0.02fF
C4575 VBIAS.n1333 GND 0.02fF
C4576 VBIAS.n1334 GND 0.01fF
C4577 VBIAS.n1335 GND 0.01fF
C4578 VBIAS.n1336 GND 0.00fF
C4579 VBIAS.n1337 GND 0.00fF
C4580 VBIAS.n1338 GND 0.01fF
C4581 VBIAS.n1339 GND 0.03fF
C4582 VBIAS.n1340 GND 0.03fF
C4583 VBIAS.n1341 GND 0.01fF
C4584 VBIAS.n1342 GND 0.04fF
C4585 VBIAS.n1343 GND 0.01fF
C4586 VBIAS.n1344 GND 0.01fF
C4587 VBIAS.n1345 GND 0.01fF
C4588 VBIAS.n1346 GND 0.01fF
C4589 VBIAS.n1347 GND 0.03fF
C4590 VBIAS.n1348 GND 0.02fF
C4591 VBIAS.n1349 GND 0.01fF
C4592 VBIAS.n1350 GND 0.01fF
C4593 VBIAS.n1351 GND 0.00fF
C4594 VBIAS.n1352 GND 0.00fF
C4595 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE GND 0.01fF
C4596 VBIAS.n1353 GND 0.01fF
C4597 VBIAS.n1354 GND 0.01fF
C4598 VBIAS.n1355 GND 0.02fF
C4599 VBIAS.n1356 GND 0.01fF
C4600 VBIAS.n1357 GND 0.00fF
C4601 VBIAS.n1358 GND 0.04fF
C4602 VBIAS.n1359 GND 0.00fF
C4603 VBIAS.n1360 GND 0.01fF
C4604 VBIAS.n1361 GND 0.01fF
C4605 VBIAS.n1362 GND 0.02fF
C4606 VBIAS.n1363 GND 0.01fF
C4607 VBIAS.n1364 GND 0.00fF
C4608 VBIAS.n1365 GND 0.01fF
C4609 VBIAS.n1366 GND 0.01fF
C4610 VBIAS.n1367 GND 0.00fF
C4611 VBIAS.n1368 GND 0.02fF
C4612 VBIAS.n1369 GND 0.00fF
C4613 VBIAS.n1370 GND 0.12fF
C4614 VBIAS.n1371 GND 0.01fF
C4615 VBIAS.n1372 GND 0.01fF
C4616 VBIAS.n1373 GND 0.02fF
C4617 VBIAS.n1374 GND 0.00fF
C4618 VBIAS.n1375 GND 0.01fF
C4619 VBIAS.n1376 GND 0.00fF
C4620 VBIAS.n1377 GND 0.00fF
C4621 VBIAS.n1378 GND 0.00fF
C4622 VBIAS.n1379 GND 0.01fF
C4623 VBIAS.n1380 GND 0.01fF
C4624 VBIAS.n1381 GND 0.01fF
C4625 VBIAS.n1382 GND 0.01fF
C4626 VBIAS.n1383 GND 0.01fF
C4627 VBIAS.n1384 GND 0.01fF
C4628 VBIAS.n1385 GND 0.01fF
C4629 VBIAS.n1386 GND 0.01fF
C4630 VBIAS.n1387 GND 0.05fF
C4631 VBIAS.n1388 GND 0.16fF
C4632 VBIAS.n1389 GND 0.03fF
C4633 VBIAS.n1390 GND 0.03fF
C4634 VBIAS.n1391 GND 0.01fF
C4635 VBIAS.n1392 GND 0.04fF
C4636 VBIAS.n1393 GND 0.04fF
C4637 VBIAS.n1394 GND 0.01fF
C4638 VBIAS.n1395 GND 0.04fF
C4639 VBIAS.n1396 GND 0.03fF
C4640 VBIAS.n1397 GND 0.01fF
C4641 VBIAS.n1398 GND 0.25fF
C4642 VBIAS.n1399 GND 0.63fF
C4643 VBIAS.n1400 GND 0.04fF
C4644 VBIAS.n1401 GND 0.01fF
C4645 VBIAS.n1402 GND 0.02fF
C4646 VBIAS.n1403 GND 0.02fF
C4647 VBIAS.n1404 GND 0.01fF
C4648 VBIAS.n1405 GND 0.01fF
C4649 VBIAS.n1406 GND 0.01fF
C4650 VBIAS.t13 GND 0.20fF $ **FLOATING
C4651 VBIAS.n1407 GND 0.03fF
C4652 VBIAS.n1408 GND 0.12fF
C4653 VBIAS.n1409 GND 0.02fF
C4654 VBIAS.n1410 GND 0.04fF
C4655 VBIAS.n1411 GND 0.01fF
C4656 VBIAS.n1412 GND 0.01fF
C4657 VBIAS.n1413 GND 0.01fF
C4658 VBIAS.n1414 GND 0.01fF
C4659 VBIAS.n1415 GND 0.01fF
C4660 VBIAS.n1416 GND 0.01fF
C4661 VBIAS.n1417 GND 0.00fF
C4662 VBIAS.n1418 GND 0.01fF
C4663 VBIAS.n1419 GND 0.00fF
C4664 VBIAS.t38 GND 0.20fF $ **FLOATING
C4665 VBIAS.n1420 GND 0.12fF
C4666 VBIAS.n1421 GND 0.01fF
C4667 VBIAS.n1422 GND 0.01fF
C4668 VBIAS.n1423 GND 0.02fF
C4669 VBIAS.n1424 GND 0.00fF
C4670 VBIAS.n1425 GND 0.01fF
C4671 VBIAS.n1426 GND 0.01fF
C4672 VBIAS.n1427 GND 0.00fF
C4673 VBIAS.n1428 GND 0.01fF
C4674 VBIAS.n1429 GND 0.01fF
C4675 VBIAS.n1430 GND 0.01fF
C4676 VBIAS.n1431 GND 0.02fF
C4677 VBIAS.n1432 GND 0.02fF
C4678 VBIAS.n1433 GND 0.01fF
C4679 VBIAS.n1434 GND 0.04fF
C4680 VBIAS.n1435 GND 0.01fF
C4681 VBIAS.n1436 GND 0.02fF
C4682 VBIAS.n1437 GND 0.02fF
C4683 VBIAS.n1438 GND 0.01fF
C4684 VBIAS.n1439 GND 0.01fF
C4685 VBIAS.n1440 GND 0.01fF
C4686 VBIAS.t22 GND 0.20fF $ **FLOATING
C4687 VBIAS.n1441 GND 0.03fF
C4688 VBIAS.n1442 GND 0.12fF
C4689 VBIAS.n1443 GND 0.02fF
C4690 VBIAS.n1444 GND 0.04fF
C4691 VBIAS.n1445 GND 0.01fF
C4692 VBIAS.n1446 GND 0.01fF
C4693 VBIAS.n1447 GND 0.01fF
C4694 VBIAS.n1448 GND 0.01fF
C4695 VBIAS.n1449 GND 0.01fF
C4696 VBIAS.n1450 GND 0.01fF
C4697 VBIAS.n1451 GND 0.00fF
C4698 VBIAS.n1452 GND 0.01fF
C4699 VBIAS.n1453 GND 0.00fF
C4700 VBIAS.t34 GND 0.20fF $ **FLOATING
C4701 VBIAS.n1454 GND 0.12fF
C4702 VBIAS.n1455 GND 0.01fF
C4703 VBIAS.n1456 GND 0.01fF
C4704 VBIAS.n1457 GND 0.02fF
C4705 VBIAS.n1458 GND 0.00fF
C4706 VBIAS.n1459 GND 0.01fF
C4707 VBIAS.n1460 GND 0.01fF
C4708 VBIAS.n1461 GND 0.00fF
C4709 VBIAS.n1462 GND 0.01fF
C4710 VBIAS.n1463 GND 0.01fF
C4711 VBIAS.n1464 GND 0.01fF
C4712 VBIAS.n1465 GND 0.02fF
C4713 VBIAS.n1466 GND 0.02fF
C4714 VBIAS.n1467 GND 0.01fF
C4715 VBIAS.n1468 GND 0.01fF
C4716 VBIAS.n1469 GND 0.01fF
C4717 VBIAS.n1470 GND 0.01fF
C4718 VBIAS.n1471 GND 0.01fF
C4719 VBIAS.n1472 GND 0.01fF
C4720 VBIAS.n1473 GND 0.00fF
C4721 VBIAS.n1474 GND 0.01fF
C4722 VBIAS.n1475 GND 0.00fF
C4723 VBIAS.t36 GND 0.20fF $ **FLOATING
C4724 VBIAS.n1476 GND 0.12fF
C4725 VBIAS.n1477 GND 0.01fF
C4726 VBIAS.n1478 GND 0.01fF
C4727 VBIAS.n1479 GND 0.02fF
C4728 VBIAS.n1480 GND 0.00fF
C4729 VBIAS.n1481 GND 0.01fF
C4730 VBIAS.n1482 GND 0.01fF
C4731 VBIAS.n1483 GND 0.00fF
C4732 VBIAS.n1484 GND 0.01fF
C4733 VBIAS.n1485 GND 0.01fF
C4734 VBIAS.n1486 GND 0.03fF
C4735 VBIAS.n1487 GND 0.03fF
C4736 VBIAS.n1488 GND 0.01fF
C4737 VBIAS.n1489 GND 0.04fF
C4738 VBIAS.n1490 GND 0.01fF
C4739 VBIAS.n1491 GND 0.01fF
C4740 VBIAS.n1492 GND 0.01fF
C4741 VBIAS.n1493 GND 0.01fF
C4742 VBIAS.n1494 GND 0.03fF
C4743 VBIAS.t12 GND 0.20fF $ **FLOATING
C4744 VBIAS.n1495 GND 0.12fF
C4745 VBIAS.n1496 GND 0.02fF
C4746 VBIAS.n1497 GND 0.04fF
C4747 VBIAS.n1498 GND 0.01fF
C4748 VBIAS.n1499 GND 0.01fF
C4749 VBIAS.n1500 GND 0.01fF
C4750 VBIAS.n1501 GND 0.01fF
C4751 VBIAS.n1502 GND 0.03fF
C4752 VBIAS.n1503 GND 0.02fF
C4753 VBIAS.n1504 GND 0.01fF
C4754 VBIAS.n1505 GND 0.01fF
C4755 VBIAS.n1506 GND 0.00fF
C4756 VBIAS.n1507 GND 0.00fF
C4757 VBIAS.n1508 GND 0.00fF
C4758 VBIAS.n1509 GND 0.01fF
C4759 VBIAS.n1510 GND 0.01fF
C4760 VBIAS.n1511 GND 0.01fF
C4761 VBIAS.n1512 GND 0.00fF
C4762 VBIAS.n1513 GND 0.01fF
C4763 VBIAS.n1514 GND 0.04fF
C4764 VBIAS.n1515 GND 0.00fF
C4765 VBIAS.n1516 GND 0.01fF
C4766 VBIAS.n1517 GND 0.01fF
C4767 VBIAS.n1518 GND 0.01fF
C4768 VBIAS.n1519 GND 0.01fF
C4769 VBIAS.n1520 GND 0.00fF
C4770 VBIAS.n1521 GND 0.00fF
C4771 VBIAS.n1522 GND 0.00fF
C4772 VBIAS.n1523 GND 0.01fF
C4773 VBIAS.n1524 GND 0.01fF
C4774 VBIAS.n1525 GND 0.02fF
C4775 VBIAS.n1526 GND 0.02fF
C4776 VBIAS.n1527 GND 0.01fF
C4777 VBIAS.n1528 GND 0.01fF
C4778 VBIAS.t24 GND 0.20fF $ **FLOATING
C4779 VBIAS.n1529 GND 0.03fF
C4780 VBIAS.n1530 GND 0.12fF
C4781 VBIAS.n1531 GND 0.02fF
C4782 VBIAS.n1532 GND 0.04fF
C4783 VBIAS.n1533 GND 0.01fF
C4784 VBIAS.n1534 GND 0.01fF
C4785 VBIAS.n1535 GND 0.00fF
C4786 VBIAS.n1536 GND 0.01fF
C4787 VBIAS.n1537 GND 0.00fF
C4788 VBIAS.t37 GND 0.20fF $ **FLOATING
C4789 VBIAS.n1538 GND 0.12fF
C4790 VBIAS.n1539 GND 0.01fF
C4791 VBIAS.n1540 GND 0.01fF
C4792 VBIAS.n1541 GND 0.02fF
C4793 VBIAS.n1542 GND 0.00fF
C4794 VBIAS.n1543 GND 0.01fF
C4795 VBIAS.n1544 GND 0.00fF
C4796 VBIAS.n1545 GND 0.01fF
C4797 VBIAS.n1546 GND 0.01fF
C4798 VBIAS.n1547 GND 0.01fF
C4799 VBIAS.n1548 GND 0.01fF
C4800 VBIAS.n1549 GND 0.01fF
C4801 VBIAS.n1550 GND 0.01fF
C4802 VBIAS.n1551 GND 0.01fF
C4803 VBIAS.n1552 GND 0.01fF
C4804 VBIAS.n1553 GND 0.05fF
C4805 VBIAS.n1554 GND 0.10fF
C4806 VBIAS.n1555 GND 0.01fF
C4807 VBIAS.n1556 GND 0.04fF
C4808 VBIAS.n1557 GND 0.04fF
C4809 VBIAS.n1558 GND 0.01fF
C4810 VBIAS.n1559 GND 0.04fF
C4811 VBIAS.n1560 GND 0.03fF
C4812 VBIAS.n1561 GND 0.01fF
C4813 VBIAS.n1562 GND 0.17fF
C4814 VBIAS.n1563 GND 0.01fF
C4815 VBIAS.n1564 GND 0.01fF
C4816 VBIAS.n1565 GND 0.01fF
C4817 VBIAS.n1566 GND 0.01fF
C4818 VBIAS.n1567 GND 0.01fF
C4819 VBIAS.n1568 GND 0.00fF
C4820 VBIAS.n1569 GND 0.01fF
C4821 VBIAS.n1570 GND 0.00fF
C4822 VBIAS.t29 GND 0.20fF $ **FLOATING
C4823 VBIAS.n1571 GND 0.12fF
C4824 VBIAS.n1572 GND 0.01fF
C4825 VBIAS.n1573 GND 0.01fF
C4826 VBIAS.n1574 GND 0.02fF
C4827 VBIAS.n1575 GND 0.00fF
C4828 VBIAS.n1576 GND 0.01fF
C4829 VBIAS.n1577 GND 0.01fF
C4830 VBIAS.n1578 GND 0.00fF
C4831 VBIAS.n1579 GND 0.01fF
C4832 VBIAS.n1580 GND 0.01fF
C4833 VBIAS.n1581 GND 0.03fF
C4834 VBIAS.n1582 GND 0.03fF
C4835 VBIAS.n1583 GND 0.01fF
C4836 VBIAS.n1584 GND 0.04fF
C4837 VBIAS.n1585 GND 0.01fF
C4838 VBIAS.n1586 GND 0.01fF
C4839 VBIAS.n1587 GND 0.01fF
C4840 VBIAS.n1588 GND 0.01fF
C4841 VBIAS.t16 GND 0.20fF $ **FLOATING
C4842 VBIAS.n1589 GND 0.03fF
C4843 VBIAS.n1590 GND 0.12fF
C4844 VBIAS.n1591 GND 0.02fF
C4845 VBIAS.n1592 GND 0.04fF
C4846 VBIAS.n1593 GND 0.01fF
C4847 VBIAS.n1594 GND 0.01fF
C4848 VBIAS.n1595 GND 0.01fF
C4849 VBIAS.n1596 GND 0.01fF
C4850 VBIAS.n1597 GND 0.03fF
C4851 VBIAS.n1598 GND 0.02fF
C4852 VBIAS.n1599 GND 0.01fF
C4853 VBIAS.n1600 GND 0.01fF
C4854 VBIAS.n1601 GND 0.00fF
C4855 VBIAS.n1602 GND 0.00fF
C4856 VBIAS.n1603 GND 0.00fF
C4857 VBIAS.n1604 GND 0.01fF
C4858 VBIAS.n1605 GND 0.01fF
C4859 VBIAS.n1606 GND 0.01fF
C4860 VBIAS.n1607 GND 0.00fF
C4861 VBIAS.n1608 GND 0.01fF
C4862 VBIAS.n1609 GND 0.04fF
C4863 VBIAS.n1610 GND 0.00fF
C4864 VBIAS.n1611 GND 0.01fF
C4865 VBIAS.n1612 GND 0.01fF
C4866 VBIAS.n1613 GND 0.01fF
C4867 VBIAS.n1614 GND 0.01fF
C4868 VBIAS.n1615 GND 0.00fF
C4869 VBIAS.n1616 GND 0.00fF
C4870 VBIAS.n1617 GND 0.00fF
C4871 VBIAS.n1618 GND 0.01fF
C4872 VBIAS.n1619 GND 0.01fF
C4873 VBIAS.n1620 GND 0.02fF
C4874 VBIAS.n1621 GND 0.02fF
C4875 VBIAS.n1622 GND 0.01fF
C4876 VBIAS.n1623 GND 0.01fF
C4877 VBIAS.t14 GND 0.20fF $ **FLOATING
C4878 VBIAS.n1624 GND 0.03fF
C4879 VBIAS.n1625 GND 0.12fF
C4880 VBIAS.n1626 GND 0.02fF
C4881 VBIAS.n1627 GND 0.04fF
C4882 VBIAS.n1628 GND 0.01fF
C4883 VBIAS.n1629 GND 0.01fF
C4884 VBIAS.n1630 GND 0.00fF
C4885 VBIAS.n1631 GND 0.01fF
C4886 VBIAS.n1632 GND 0.00fF
C4887 VBIAS.t39 GND 0.20fF $ **FLOATING
C4888 VBIAS.n1633 GND 0.12fF
C4889 VBIAS.n1634 GND 0.01fF
C4890 VBIAS.n1635 GND 0.01fF
C4891 VBIAS.n1636 GND 0.02fF
C4892 VBIAS.n1637 GND 0.00fF
C4893 VBIAS.n1638 GND 0.01fF
C4894 VBIAS.n1639 GND 0.00fF
C4895 VBIAS.n1640 GND 0.01fF
C4896 VBIAS.n1641 GND 0.01fF
C4897 VBIAS.n1642 GND 0.01fF
C4898 VBIAS.n1643 GND 0.01fF
C4899 VBIAS.n1644 GND 0.01fF
C4900 VBIAS.n1645 GND 0.01fF
C4901 VBIAS.n1646 GND 0.01fF
C4902 VBIAS.n1647 GND 0.01fF
C4903 VBIAS.n1648 GND 0.05fF
C4904 VBIAS.n1649 GND 0.17fF
C4905 VBIAS.n1650 GND 0.03fF
C4906 VBIAS.n1651 GND 0.03fF
C4907 VBIAS.n1652 GND 0.01fF
C4908 VBIAS.n1653 GND 0.04fF
C4909 VBIAS.n1654 GND 0.04fF
C4910 VBIAS.n1655 GND 0.01fF
C4911 VBIAS.n1656 GND 0.04fF
C4912 VBIAS.n1657 GND 0.03fF
C4913 VBIAS.n1658 GND 0.01fF
C4914 VBIAS.n1659 GND 0.17fF
C4915 VBIAS.n1660 GND 0.01fF
C4916 VBIAS.n1661 GND 0.01fF
C4917 VBIAS.n1662 GND 0.01fF
C4918 VBIAS.n1663 GND 0.01fF
C4919 VBIAS.n1664 GND 0.01fF
C4920 VBIAS.n1665 GND 0.00fF
C4921 VBIAS.n1666 GND 0.01fF
C4922 VBIAS.n1667 GND 0.00fF
C4923 VBIAS.t2 GND 0.20fF $ **FLOATING
C4924 VBIAS.n1668 GND 0.12fF
C4925 VBIAS.n1669 GND 0.01fF
C4926 VBIAS.n1670 GND 0.01fF
C4927 VBIAS.n1671 GND 0.02fF
C4928 VBIAS.n1672 GND 0.00fF
C4929 VBIAS.n1673 GND 0.01fF
C4930 VBIAS.n1674 GND 0.01fF
C4931 VBIAS.n1675 GND 0.00fF
C4932 VBIAS.n1676 GND 0.01fF
C4933 VBIAS.n1677 GND 0.01fF
C4934 VBIAS.n1678 GND 0.03fF
C4935 VBIAS.n1679 GND 0.03fF
C4936 VBIAS.n1680 GND 0.01fF
C4937 VBIAS.n1681 GND 0.04fF
C4938 VBIAS.n1682 GND 0.01fF
C4939 VBIAS.n1683 GND 0.01fF
C4940 VBIAS.n1684 GND 0.01fF
C4941 VBIAS.n1685 GND 0.01fF
C4942 VBIAS.t4 GND 0.20fF $ **FLOATING
C4943 VBIAS.n1686 GND 0.03fF
C4944 VBIAS.n1687 GND 0.12fF
C4945 VBIAS.n1688 GND 0.02fF
C4946 VBIAS.n1689 GND 0.04fF
C4947 VBIAS.n1690 GND 0.01fF
C4948 VBIAS.n1691 GND 0.01fF
C4949 VBIAS.n1692 GND 0.01fF
C4950 VBIAS.n1693 GND 0.01fF
C4951 VBIAS.n1694 GND 0.03fF
C4952 VBIAS.n1695 GND 0.02fF
C4953 VBIAS.n1696 GND 0.01fF
C4954 VBIAS.n1697 GND 0.01fF
C4955 VBIAS.n1698 GND 0.00fF
C4956 VBIAS.n1699 GND 0.00fF
C4957 VBIAS.n1700 GND 0.00fF
C4958 VBIAS.n1701 GND 0.01fF
C4959 VBIAS.n1702 GND 0.01fF
C4960 VBIAS.n1703 GND 0.01fF
C4961 VBIAS.n1704 GND 0.00fF
C4962 VBIAS.n1705 GND 0.01fF
C4963 VBIAS.n1706 GND 0.04fF
C4964 VBIAS.n1707 GND 0.00fF
C4965 VBIAS.n1708 GND 0.01fF
C4966 VBIAS.n1709 GND 0.01fF
C4967 VBIAS.n1710 GND 0.01fF
C4968 VBIAS.n1711 GND 0.01fF
C4969 VBIAS.n1712 GND 0.00fF
C4970 VBIAS.n1713 GND 0.00fF
C4971 VBIAS.n1714 GND 0.00fF
C4972 VBIAS.n1715 GND 0.01fF
C4973 VBIAS.n1716 GND 0.01fF
C4974 VBIAS.n1717 GND 0.02fF
C4975 VBIAS.n1718 GND 0.02fF
C4976 VBIAS.n1719 GND 0.01fF
C4977 VBIAS.n1720 GND 0.01fF
C4978 VBIAS.t6 GND 0.20fF $ **FLOATING
C4979 VBIAS.n1721 GND 0.03fF
C4980 VBIAS.n1722 GND 0.12fF
C4981 VBIAS.n1723 GND 0.02fF
C4982 VBIAS.n1724 GND 0.04fF
C4983 VBIAS.n1725 GND 0.01fF
C4984 VBIAS.n1726 GND 0.01fF
C4985 VBIAS.n1727 GND 0.00fF
C4986 VBIAS.n1728 GND 0.01fF
C4987 VBIAS.n1729 GND 0.00fF
C4988 VBIAS.t0 GND 0.20fF $ **FLOATING
C4989 VBIAS.n1730 GND 0.12fF
C4990 VBIAS.n1731 GND 0.01fF
C4991 VBIAS.n1732 GND 0.01fF
C4992 VBIAS.n1733 GND 0.02fF
C4993 VBIAS.n1734 GND 0.00fF
C4994 VBIAS.n1735 GND 0.01fF
C4995 VBIAS.n1736 GND 0.00fF
C4996 VBIAS.n1737 GND 0.01fF
C4997 VBIAS.n1738 GND 0.01fF
C4998 VBIAS.n1739 GND 0.01fF
C4999 VBIAS.n1740 GND 0.01fF
C5000 VBIAS.n1741 GND 0.01fF
C5001 VBIAS.n1742 GND 0.01fF
C5002 VBIAS.n1743 GND 0.01fF
C5003 VBIAS.n1744 GND 0.01fF
C5004 VBIAS.n1745 GND 0.05fF
C5005 VBIAS.n1746 GND 0.17fF
C5006 VBIAS.n1747 GND 0.03fF
C5007 VBIAS.n1748 GND 0.03fF
C5008 VBIAS.n1749 GND 0.01fF
C5009 VBIAS.n1750 GND 0.04fF
C5010 VBIAS.n1751 GND 0.04fF
C5011 VBIAS.n1752 GND 0.01fF
C5012 VBIAS.n1753 GND 0.04fF
C5013 VBIAS.n1754 GND 0.03fF
C5014 VBIAS.n1755 GND 0.01fF
C5015 VBIAS.n1756 GND 0.17fF
C5016 VBIAS.n1757 GND 0.17fF
C5017 VBIAS.n1758 GND 0.04fF
C5018 VBIAS.n1759 GND 0.01fF
C5019 VBIAS.n1760 GND 0.01fF
C5020 VBIAS.n1761 GND 0.01fF
C5021 VBIAS.n1762 GND 0.01fF
C5022 VBIAS.n1763 GND 0.03fF
C5023 VBIAS.n1764 GND 0.03fF
C5024 VBIAS.n1765 GND 0.04fF
C5025 VBIAS.n1766 GND 0.01fF
C5026 VBIAS.n1767 GND 0.01fF
C5027 VBIAS.n1768 GND 0.00fF
C5028 VBIAS.n1769 GND 0.01fF
C5029 VBIAS.n1770 GND 0.01fF
C5030 VBIAS.n1771 GND 0.01fF
C5031 VBIAS.n1772 GND 0.01fF
C5032 VBIAS.n1773 GND 0.01fF
C5033 VBIAS.n1774 GND 0.04fF
C5034 VBIAS.n1775 GND 0.00fF
C5035 VBIAS.n1776 GND 0.01fF
C5036 VBIAS.n1777 GND 0.00fF
C5037 VBIAS.n1778 GND 0.01fF
C5038 VBIAS.n1779 GND 0.01fF
C5039 VBIAS.n1780 GND 0.01fF
C5040 VBIAS.n1781 GND 0.01fF
C5041 VBIAS.n1782 GND 0.01fF
C5042 VBIAS.n1783 GND 0.01fF
C5043 VBIAS.n1784 GND 0.00fF
C5044 VBIAS.n1785 GND 0.01fF
C5045 VBIAS.n1786 GND 0.01fF
C5046 VBIAS.n1787 GND 0.00fF
C5047 VBIAS.n1788 GND 0.00fF
C5048 VBIAS.n1789 GND 0.00fF
C5049 VBIAS.n1790 GND 0.01fF
C5050 VBIAS.n1791 GND 0.01fF
C5051 VBIAS.n1792 GND 0.01fF
C5052 VBIAS.n1793 GND 0.04fF
C5053 VBIAS.n1794 GND 0.03fF
C5054 VBIAS.n1795 GND 0.03fF
C5055 VBIAS.n1796 GND 0.02fF
C5056 VBIAS.n1797 GND 0.01fF
C5057 VBIAS.n1798 GND 0.00fF
C5058 VBIAS.t27 GND 0.20fF $ **FLOATING
C5059 VBIAS.n1799 GND 0.12fF
C5060 VBIAS.n1800 GND 0.01fF
C5061 VBIAS.n1801 GND 0.01fF
C5062 VBIAS.n1802 GND 0.02fF
C5063 VBIAS.n1803 GND 0.00fF
C5064 VBIAS.n1804 GND 0.01fF
C5065 VBIAS.n1805 GND 0.00fF
C5066 VBIAS.n1806 GND 0.01fF
C5067 VBIAS.n1807 GND 0.01fF
C5068 VBIAS.n1808 GND 0.01fF
C5069 VBIAS.n1809 GND 0.01fF
C5070 VBIAS.n1810 GND 0.01fF
C5071 VBIAS.n1811 GND 0.01fF
C5072 VBIAS.t23 GND 0.20fF $ **FLOATING
C5073 VBIAS.n1812 GND 0.03fF
C5074 VBIAS.n1813 GND 0.12fF
C5075 VBIAS.n1814 GND 0.02fF
C5076 VBIAS.n1815 GND 0.04fF
C5077 VBIAS.n1816 GND 0.01fF
C5078 VBIAS.n1817 GND 0.01fF
C5079 VBIAS.n1818 GND 0.01fF
C5080 VBIAS.n1819 GND 0.01fF
C5081 VBIAS.n1820 GND 0.04fF
C5082 VBIAS.n1821 GND 0.01fF
C5083 VBIAS.n1822 GND 0.01fF
C5084 VBIAS.n1823 GND 0.17fF
C5085 VBIAS.n1824 GND 0.17fF
C5086 VBIAS.n1825 GND 0.04fF
C5087 VBIAS.n1826 GND 0.01fF
C5088 VBIAS.n1827 GND 0.01fF
C5089 VBIAS.n1828 GND 0.01fF
C5090 VBIAS.n1829 GND 0.01fF
C5091 VBIAS.n1830 GND 0.03fF
C5092 VBIAS.n1831 GND 0.03fF
C5093 VBIAS.n1832 GND 0.04fF
C5094 VBIAS.n1833 GND 0.01fF
C5095 VBIAS.n1834 GND 0.01fF
C5096 VBIAS.n1835 GND 0.00fF
C5097 VBIAS.n1836 GND 0.01fF
C5098 VBIAS.n1837 GND 0.01fF
C5099 VBIAS.n1838 GND 0.01fF
C5100 VBIAS.n1839 GND 0.01fF
C5101 VBIAS.n1840 GND 0.01fF
C5102 VBIAS.n1841 GND 0.04fF
C5103 VBIAS.n1842 GND 0.00fF
C5104 VBIAS.n1843 GND 0.01fF
C5105 VBIAS.n1844 GND 0.00fF
C5106 VBIAS.n1845 GND 0.01fF
C5107 VBIAS.n1846 GND 0.01fF
C5108 VBIAS.n1847 GND 0.01fF
C5109 VBIAS.n1848 GND 0.01fF
C5110 VBIAS.n1849 GND 0.01fF
C5111 VBIAS.n1850 GND 0.01fF
C5112 VBIAS.n1851 GND 0.00fF
C5113 VBIAS.n1852 GND 0.01fF
C5114 VBIAS.n1853 GND 0.01fF
C5115 VBIAS.n1854 GND 0.00fF
C5116 VBIAS.n1855 GND 0.00fF
C5117 VBIAS.n1856 GND 0.00fF
C5118 VBIAS.n1857 GND 0.01fF
C5119 VBIAS.n1858 GND 0.01fF
C5120 VBIAS.n1859 GND 0.01fF
C5121 VBIAS.n1860 GND 0.04fF
C5122 VBIAS.n1861 GND 0.03fF
C5123 VBIAS.n1862 GND 0.03fF
C5124 VBIAS.n1863 GND 0.02fF
C5125 VBIAS.n1864 GND 0.01fF
C5126 VBIAS.n1865 GND 0.00fF
C5127 VBIAS.t26 GND 0.20fF $ **FLOATING
C5128 VBIAS.n1866 GND 0.12fF
C5129 VBIAS.n1867 GND 0.01fF
C5130 VBIAS.n1868 GND 0.01fF
C5131 VBIAS.n1869 GND 0.02fF
C5132 VBIAS.n1870 GND 0.00fF
C5133 VBIAS.n1871 GND 0.01fF
C5134 VBIAS.n1872 GND 0.00fF
C5135 VBIAS.n1873 GND 0.01fF
C5136 VBIAS.n1874 GND 0.01fF
C5137 VBIAS.n1875 GND 0.01fF
C5138 VBIAS.n1876 GND 0.01fF
C5139 VBIAS.n1877 GND 0.01fF
C5140 VBIAS.n1878 GND 0.01fF
C5141 VBIAS.t25 GND 0.20fF $ **FLOATING
C5142 VBIAS.n1879 GND 0.03fF
C5143 VBIAS.n1880 GND 0.12fF
C5144 VBIAS.n1881 GND 0.02fF
C5145 VBIAS.n1882 GND 0.04fF
C5146 VBIAS.n1883 GND 0.01fF
C5147 VBIAS.n1884 GND 0.01fF
C5148 VBIAS.n1885 GND 0.01fF
C5149 VBIAS.n1886 GND 0.01fF
C5150 VBIAS.n1887 GND 0.04fF
C5151 VBIAS.n1888 GND 0.01fF
C5152 VBIAS.n1889 GND 0.01fF
C5153 VBIAS.n1890 GND 0.26fF
C5154 VBIAS.n1891 GND 1.45fF
C5155 VBIAS.n1892 GND 7.96fF
C5156 VBIAS.n1893 GND 5.76fF
C5157 VBIAS.n1895 GND 0.16fF
C5158 VBIAS.n1897 GND 0.19fF
C5159 VBIAS.n1899 GND 0.16fF
C5160 VBIAS.n1901 GND 0.16fF
C5161 VBIAS.n1903 GND 0.16fF
C5162 VBIAS.n1905 GND 0.19fF
C5163 VBIAS.n1907 GND 0.16fF
C5164 VBIAS.n1909 GND 0.16fF
C5165 VBIAS.n1911 GND 0.19fF
C5166 VBIAS.n1913 GND 0.12fF
C5167 VBIAS.n1914 GND 0.33fF
C5168 VBIAS.n1915 GND 0.01fF
C5169 VBIAS.n1916 GND 0.01fF
C5170 VBIAS.n1917 GND 0.00fF
C5171 VBIAS.n1918 GND 0.00fF
C5172 VBIAS.n1919 GND 0.02fF
C5173 VBIAS.n1920 GND 0.02fF
C5174 VBIAS.n1921 GND 0.00fF
C5175 VBIAS.n1922 GND 0.00fF
C5176 VBIAS.n1924 GND 0.13fF
C5177 VBIAS.n1925 GND 0.00fF
C5178 VBIAS.n1926 GND 0.01fF
C5179 VBIAS.n1927 GND 0.00fF
C5180 VBIAS.n1928 GND 0.01fF
C5181 VBIAS.n1929 GND 0.00fF
C5182 VBIAS.n1930 GND 0.00fF
C5183 VBIAS.n1931 GND 0.00fF
C5184 VBIAS.n1932 GND 0.00fF
C5185 VBIAS.n1933 GND 0.01fF
C5186 VBIAS.n1934 GND 0.01fF
C5187 VBIAS.n1935 GND 0.01fF
C5188 VBIAS.n1936 GND 0.00fF
C5189 VBIAS.n1938 GND 0.06fF
C5190 VBIAS.n1939 GND 0.01fF
C5191 VBIAS.n1940 GND 0.00fF
C5192 VBIAS.n1941 GND 0.01fF
C5193 VBIAS.n1942 GND 0.01fF
C5194 VBIAS.t3 GND 0.17fF $ **FLOATING
C5195 VBIAS.t5 GND 0.17fF $ **FLOATING
C5196 VBIAS.n1943 GND 0.51fF
C5197 VBIAS.n1944 GND 0.07fF
C5198 VBIAS.n1945 GND 0.39fF
C5199 VBIAS.n1946 GND 0.01fF
C5200 VBIAS.n1947 GND 0.00fF
C5201 VBIAS.n1948 GND 0.00fF
C5202 VBIAS.n1949 GND 0.01fF
C5203 VBIAS.n1950 GND 0.01fF
C5204 VBIAS.n1951 GND 0.01fF
C5205 VBIAS.n1952 GND 0.01fF
C5206 VBIAS.n1953 GND 0.00fF
C5207 VBIAS.n1954 GND 0.01fF
C5208 VBIAS.n1955 GND 0.00fF
C5209 VBIAS.n1956 GND 0.00fF
C5210 VBIAS.n1957 GND 0.00fF
C5211 VBIAS.n1958 GND 0.00fF
C5212 VBIAS.n1959 GND 0.00fF
C5213 VBIAS.n1960 GND 0.01fF
C5214 VBIAS.n1961 GND 0.01fF
C5215 VBIAS.n1962 GND 0.01fF
C5216 VBIAS.n1963 GND 0.01fF
C5217 VBIAS.n1964 GND 0.01fF
C5218 VBIAS.n1965 GND 0.00fF
C5219 VBIAS.n1966 GND 0.01fF
C5220 VBIAS.n1967 GND 0.00fF
C5221 VBIAS.n1968 GND 0.00fF
C5222 VBIAS.n1969 GND 0.00fF
C5223 VBIAS.n1970 GND 0.00fF
C5224 VBIAS.n1971 GND 0.00fF
C5225 VBIAS.n1972 GND 0.00fF
C5226 VBIAS.n1973 GND 0.01fF
C5227 VBIAS.n1974 GND 0.01fF
C5228 VBIAS.n1975 GND 0.01fF
C5229 VBIAS.n1976 GND 0.06fF
C5230 VBIAS.n1977 GND 0.06fF
C5231 VBIAS.n1978 GND 0.05fF
C5232 VBIAS.n1979 GND 0.06fF
C5233 VBIAS.n1980 GND 0.62fF
C5234 buffer_mirror_0/buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_10/DRAIN GND 0.62fF
.ends



**** end user architecture code
**.ends
** flattened .save nodes
.end
