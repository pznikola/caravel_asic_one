* NGSPICE file created from buffer.ext - technology: sky130B

.subckt rf_nfet_01v8_lvt_aM04W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
X0 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8_lvt ad=4.242e+12p pd=3.198e+07u as=2.828e+12p ps=2.132e+07u w=5.05e+06u l=150000u
X1 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends

.subckt buffer_input_base m5_566_1418# rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_1/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SOURCE
+ VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_0 rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_1 rf_nfet_01v8_lvt_aM04W5p00L0p15_1/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_2 rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_3 rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_4 rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_5 rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_6 rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_7 rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
.ends

.subckt buffer_input GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE
+ a_n330_n214# buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN
Xbuffer_input_base_0 buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE
+ buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE
+ GATE GATE GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE GATE
+ buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN
+ buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE GATE GATE GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN
+ GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN GATE GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE
+ buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE
+ GATE GATE buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE buffer_input_base
.ends

.subckt sky130_fd_pr__res_generic_po_TC8HWG a_n350_n423# a_n350_350#
R0 a_n350_n423# a_n350_350# sky130_fd_pr__res_generic_po w=3.5e+06u l=3.5e+06u
.ends

.subckt buffer_mirror_base rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_9/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_12/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_1/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_13/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_10/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_11/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_9/DRAIN
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_12/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_13/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SOURCE rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_11/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SOURCE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SOURCE
+ VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_0 rf_nfet_01v8_lvt_aM04W5p00L0p15_0/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_0/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_0/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_1 rf_nfet_01v8_lvt_aM04W5p00L0p15_1/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_1/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_1/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_2 rf_nfet_01v8_lvt_aM04W5p00L0p15_2/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_2/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_2/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_3 rf_nfet_01v8_lvt_aM04W5p00L0p15_3/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_3/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_3/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_4 rf_nfet_01v8_lvt_aM04W5p00L0p15_4/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_4/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_4/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_5 rf_nfet_01v8_lvt_aM04W5p00L0p15_5/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_5/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_5/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_6 rf_nfet_01v8_lvt_aM04W5p00L0p15_6/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_6/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_8 rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_8/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_7 rf_nfet_01v8_lvt_aM04W5p00L0p15_7/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_7/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_7/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_10 rf_nfet_01v8_lvt_aM04W5p00L0p15_10/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_10/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_10/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_11 rf_nfet_01v8_lvt_aM04W5p00L0p15_11/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_11/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_11/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_9 rf_nfet_01v8_lvt_aM04W5p00L0p15_9/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_9/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_9/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_12 rf_nfet_01v8_lvt_aM04W5p00L0p15_12/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_12/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_12/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
Xrf_nfet_01v8_lvt_aM04W5p00L0p15_13 rf_nfet_01v8_lvt_aM04W5p00L0p15_13/DRAIN rf_nfet_01v8_lvt_aM04W5p00L0p15_13/GATE
+ rf_nfet_01v8_lvt_aM04W5p00L0p15_13/SOURCE VSUBS rf_nfet_01v8_lvt_aM04W5p00L0p15
.ends

.subckt buffer_mirror buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN
+ buffer_mirror_base_0/VSUBS
Xbuffer_mirror_base_0 buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN buffer_mirror_base_0/VSUBS
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN buffer_mirror_base_0/VSUBS
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/DRAIN buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS
+ buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE buffer_mirror_base_0/VSUBS
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_8/GATE
+ buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS buffer_mirror_base_0/VSUBS
+ buffer_mirror_base
.ends

.subckt buffer VBIAS VDD GND OUT_P OUT_N IN_P IN_N
Xbuffer_input_0 buffer_input_0/GATE buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE
+ buffer_input_0/GATE OUT_N OUT_P buffer_input
Xsky130_fd_pr__res_generic_po_TC8HWG_0 VDD OUT_P sky130_fd_pr__res_generic_po_TC8HWG
Xsky130_fd_pr__res_generic_po_TC8HWG_1 OUT_N VDD sky130_fd_pr__res_generic_po_TC8HWG
Xbuffer_mirror_0 buffer_input_0/buffer_input_base_0/rf_nfet_01v8_lvt_aM04W5p00L0p15_6/SOURCE
+ buffer_input_0/GATE buffer_mirror
.ends

