magic
tech sky130B
magscale 1 2
timestamp 1654612318
<< pwell >>
rect 70 -194 106 -190
rect 0 -1030 70 -218
rect 1826 -1030 1896 -128
<< psubdiff >>
rect 0 -198 1896 -128
rect 0 -960 70 -198
rect 1826 -260 1896 -198
rect 1860 -898 1896 -260
rect 1826 -960 1896 -898
rect 0 -1030 1896 -960
<< psubdiffcont >>
rect 1826 -898 1860 -260
<< locali >>
rect 1826 -238 1860 -164
rect 1826 -260 1832 -238
rect 1826 -912 1832 -898
rect 1826 -994 1860 -912
<< viali >>
rect 70 -192 104 -158
rect 150 -192 184 -158
rect 230 -192 264 -158
rect 310 -192 344 -158
rect 390 -192 424 -158
rect 470 -192 504 -158
rect 550 -192 584 -158
rect 630 -192 664 -158
rect 710 -192 744 -158
rect 790 -192 824 -158
rect 870 -192 904 -158
rect 950 -192 984 -158
rect 1030 -192 1064 -158
rect 1110 -192 1144 -158
rect 1190 -192 1224 -158
rect 1270 -192 1304 -158
rect 1350 -192 1384 -158
rect 1430 -192 1464 -158
rect 1510 -192 1544 -158
rect 1590 -192 1624 -158
rect 1670 -192 1704 -158
rect 1750 -192 1784 -158
rect 30 -272 64 -238
rect 1832 -260 1866 -238
rect 1832 -272 1860 -260
rect 1860 -272 1866 -260
rect 30 -352 64 -318
rect 1832 -352 1860 -318
rect 1860 -352 1866 -318
rect 30 -432 64 -398
rect 1832 -432 1860 -398
rect 1860 -432 1866 -398
rect 30 -512 64 -478
rect 1832 -512 1860 -478
rect 1860 -512 1866 -478
rect 30 -592 64 -558
rect 1832 -592 1860 -558
rect 1860 -592 1866 -558
rect 30 -672 64 -638
rect 1832 -672 1860 -638
rect 1860 -672 1866 -638
rect 30 -752 64 -718
rect 1832 -752 1860 -718
rect 1860 -752 1866 -718
rect 30 -832 64 -798
rect 1832 -832 1860 -798
rect 1860 -832 1866 -798
rect 30 -912 64 -878
rect 1832 -898 1860 -878
rect 1860 -898 1866 -878
rect 1832 -912 1866 -898
rect 70 -1000 104 -966
rect 150 -1000 184 -966
rect 230 -1000 264 -966
rect 310 -1000 344 -966
rect 390 -1000 424 -966
rect 470 -1000 504 -966
rect 550 -1000 584 -966
rect 630 -1000 664 -966
rect 710 -1000 744 -966
rect 790 -1000 824 -966
rect 870 -1000 904 -966
rect 950 -1000 984 -966
rect 1030 -1000 1064 -966
rect 1110 -1000 1144 -966
rect 1190 -1000 1224 -966
rect 1270 -1000 1304 -966
rect 1350 -1000 1384 -966
rect 1430 -1000 1464 -966
rect 1510 -1000 1544 -966
rect 1590 -1000 1624 -966
rect 1670 -1000 1704 -966
rect 1750 -1000 1784 -966
<< metal1 >>
rect 172 2514 250 2550
rect 172 2462 184 2514
rect 238 2462 250 2514
rect 172 2434 250 2462
rect 172 2382 184 2434
rect 238 2382 250 2434
rect 172 2354 250 2382
rect 172 2302 184 2354
rect 238 2302 250 2354
rect 172 2274 250 2302
rect 172 2222 184 2274
rect 238 2222 250 2274
rect 172 2194 250 2222
rect 172 2142 184 2194
rect 238 2142 250 2194
rect 172 2114 250 2142
rect 172 2062 184 2114
rect 238 2062 250 2114
rect 172 2034 250 2062
rect 172 1982 184 2034
rect 238 1982 250 2034
rect 172 1950 250 1982
rect 1402 2514 1480 2550
rect 1402 2462 1414 2514
rect 1468 2462 1480 2514
rect 1402 2434 1480 2462
rect 1402 2382 1414 2434
rect 1468 2382 1480 2434
rect 1402 2354 1480 2382
rect 1402 2302 1414 2354
rect 1468 2302 1480 2354
rect 1402 2274 1480 2302
rect 1402 2222 1414 2274
rect 1468 2222 1480 2274
rect 1402 2194 1480 2222
rect 1402 2142 1414 2194
rect 1468 2142 1480 2194
rect 1402 2114 1480 2142
rect 1402 2062 1414 2114
rect 1468 2062 1480 2114
rect 1402 2034 1480 2062
rect 1402 1982 1414 2034
rect 1468 1982 1480 2034
rect 1402 1950 1480 1982
rect 2632 2514 2710 2550
rect 2632 2462 2644 2514
rect 2698 2462 2710 2514
rect 2632 2434 2710 2462
rect 2632 2382 2644 2434
rect 2698 2382 2710 2434
rect 2632 2354 2710 2382
rect 2632 2302 2644 2354
rect 2698 2302 2710 2354
rect 2632 2274 2710 2302
rect 2632 2222 2644 2274
rect 2698 2222 2710 2274
rect 2632 2194 2710 2222
rect 2632 2142 2644 2194
rect 2698 2142 2710 2194
rect 2632 2114 2710 2142
rect 2632 2062 2644 2114
rect 2698 2062 2710 2114
rect 2632 2034 2710 2062
rect 2632 1982 2644 2034
rect 2698 1982 2710 2034
rect 2632 1950 2710 1982
rect 554 1860 758 1864
rect 554 1850 594 1860
rect 646 1850 674 1860
rect 554 1798 590 1850
rect 646 1808 670 1850
rect 726 1808 758 1860
rect 642 1798 670 1808
rect 722 1798 758 1808
rect 948 1860 1152 1864
rect 948 1850 988 1860
rect 1040 1850 1068 1860
rect 948 1798 984 1850
rect 1040 1808 1064 1850
rect 1120 1808 1152 1860
rect 1036 1798 1064 1808
rect 1116 1798 1152 1808
rect 1736 1860 1940 1864
rect 1736 1850 1776 1860
rect 1828 1850 1856 1860
rect 1736 1798 1772 1850
rect 1828 1808 1852 1850
rect 1908 1808 1940 1860
rect 1824 1798 1852 1808
rect 1904 1798 1940 1808
rect 554 1072 590 1124
rect 642 1114 670 1124
rect 722 1114 758 1124
rect 646 1072 670 1114
rect 554 1062 594 1072
rect 646 1062 674 1072
rect 726 1062 758 1114
rect 554 1058 758 1062
rect 948 1072 984 1124
rect 1036 1114 1064 1124
rect 1116 1114 1152 1124
rect 1040 1072 1064 1114
rect 948 1062 988 1072
rect 1040 1062 1068 1072
rect 1120 1062 1152 1114
rect 948 1058 1152 1062
rect 1736 1072 1772 1124
rect 1824 1114 1852 1124
rect 1904 1114 1940 1124
rect 1828 1072 1852 1114
rect 1736 1062 1776 1072
rect 1828 1062 1856 1072
rect 1908 1062 1940 1114
rect 1736 1058 1940 1062
rect 558 1052 758 1058
rect 952 1052 1152 1058
rect 1740 1052 1940 1058
rect 558 928 758 934
rect 952 928 1152 934
rect 1346 928 1546 934
rect 1740 928 1940 934
rect 554 924 758 928
rect 554 914 594 924
rect 646 914 674 924
rect 554 862 590 914
rect 646 872 670 914
rect 726 872 758 924
rect 642 862 670 872
rect 722 862 758 872
rect 948 924 1152 928
rect 948 914 988 924
rect 1040 914 1068 924
rect 948 862 984 914
rect 1040 872 1064 914
rect 1120 872 1152 924
rect 1036 862 1064 872
rect 1116 862 1152 872
rect 1342 924 1546 928
rect 1342 914 1382 924
rect 1434 914 1462 924
rect 1342 862 1378 914
rect 1434 872 1458 914
rect 1514 872 1546 924
rect 1430 862 1458 872
rect 1510 862 1546 872
rect 1736 924 1940 928
rect 1736 914 1776 924
rect 1828 914 1856 924
rect 1736 862 1772 914
rect 1828 872 1852 914
rect 1908 872 1940 924
rect 1824 862 1852 872
rect 1904 862 1940 872
rect 558 174 758 184
rect 952 174 1152 184
rect 554 122 590 174
rect 646 122 670 174
rect 726 122 758 174
rect 948 122 984 174
rect 1040 122 1064 174
rect 1120 122 1152 174
rect 1330 180 1558 188
rect 1330 128 1378 180
rect 1430 128 1458 180
rect 1510 128 1558 180
rect 1740 174 1940 184
rect 1330 122 1558 128
rect 1736 122 1772 174
rect 1828 122 1852 174
rect 1908 122 1940 174
rect 2130 122 2166 174
rect 2218 122 2246 174
rect 2298 122 2334 174
rect 0 -158 1896 -128
rect 0 -192 70 -158
rect 104 -192 150 -158
rect 184 -192 230 -158
rect 264 -192 310 -158
rect 344 -192 390 -158
rect 424 -192 470 -158
rect 504 -192 550 -158
rect 584 -192 630 -158
rect 664 -192 710 -158
rect 744 -192 790 -158
rect 824 -192 870 -158
rect 904 -192 950 -158
rect 984 -192 1030 -158
rect 1064 -192 1110 -158
rect 1144 -192 1190 -158
rect 1224 -192 1270 -158
rect 1304 -192 1350 -158
rect 1384 -192 1430 -158
rect 1464 -192 1510 -158
rect 1544 -192 1590 -158
rect 1624 -192 1670 -158
rect 1704 -192 1750 -158
rect 1784 -192 1896 -158
rect 0 -198 1896 -192
rect 0 -238 70 -198
rect 0 -272 30 -238
rect 64 -272 70 -238
rect 0 -318 70 -272
rect 1826 -238 1896 -198
rect 1826 -272 1832 -238
rect 1866 -272 1896 -238
rect 0 -352 30 -318
rect 64 -352 70 -318
rect 0 -398 70 -352
rect 0 -432 30 -398
rect 64 -432 70 -398
rect 0 -478 70 -432
rect 0 -512 30 -478
rect 64 -512 70 -478
rect 0 -558 70 -512
rect 0 -592 30 -558
rect 64 -592 70 -558
rect 0 -638 70 -592
rect 0 -672 30 -638
rect 64 -672 70 -638
rect 0 -718 70 -672
rect 0 -752 30 -718
rect 64 -752 70 -718
rect 0 -798 70 -752
rect 0 -832 30 -798
rect 64 -832 70 -798
rect 0 -878 70 -832
rect 166 -298 598 -294
rect 166 -350 196 -298
rect 248 -350 260 -298
rect 312 -350 324 -298
rect 376 -350 388 -298
rect 440 -350 452 -298
rect 504 -350 516 -298
rect 568 -350 598 -298
rect 166 -362 598 -350
rect 166 -414 196 -362
rect 248 -414 260 -362
rect 312 -414 324 -362
rect 376 -414 388 -362
rect 440 -414 452 -362
rect 504 -414 516 -362
rect 568 -414 598 -362
rect 166 -426 598 -414
rect 166 -478 196 -426
rect 248 -478 260 -426
rect 312 -478 324 -426
rect 376 -478 388 -426
rect 440 -478 452 -426
rect 504 -478 516 -426
rect 568 -478 598 -426
rect 166 -490 598 -478
rect 166 -542 196 -490
rect 248 -542 260 -490
rect 312 -542 324 -490
rect 376 -542 388 -490
rect 440 -542 452 -490
rect 504 -542 516 -490
rect 568 -542 598 -490
rect 166 -554 598 -542
rect 166 -606 196 -554
rect 248 -606 260 -554
rect 312 -606 324 -554
rect 376 -606 388 -554
rect 440 -606 452 -554
rect 504 -606 516 -554
rect 568 -606 598 -554
rect 166 -618 598 -606
rect 166 -670 196 -618
rect 248 -670 260 -618
rect 312 -670 324 -618
rect 376 -670 388 -618
rect 440 -670 452 -618
rect 504 -670 516 -618
rect 568 -670 598 -618
rect 166 -682 598 -670
rect 166 -734 196 -682
rect 248 -734 260 -682
rect 312 -734 324 -682
rect 376 -734 388 -682
rect 440 -734 452 -682
rect 504 -734 516 -682
rect 568 -734 598 -682
rect 166 -746 598 -734
rect 166 -798 196 -746
rect 248 -798 260 -746
rect 312 -798 324 -746
rect 376 -798 388 -746
rect 440 -798 452 -746
rect 504 -798 516 -746
rect 568 -798 598 -746
rect 166 -810 598 -798
rect 166 -862 196 -810
rect 248 -862 260 -810
rect 312 -862 324 -810
rect 376 -862 388 -810
rect 440 -862 452 -810
rect 504 -862 516 -810
rect 568 -862 598 -810
rect 166 -864 598 -862
rect 1298 -298 1730 -294
rect 1298 -350 1328 -298
rect 1380 -350 1392 -298
rect 1444 -350 1456 -298
rect 1508 -350 1520 -298
rect 1572 -350 1584 -298
rect 1636 -350 1648 -298
rect 1700 -350 1730 -298
rect 1298 -362 1730 -350
rect 1298 -414 1328 -362
rect 1380 -414 1392 -362
rect 1444 -414 1456 -362
rect 1508 -414 1520 -362
rect 1572 -414 1584 -362
rect 1636 -414 1648 -362
rect 1700 -414 1730 -362
rect 1298 -426 1730 -414
rect 1298 -478 1328 -426
rect 1380 -478 1392 -426
rect 1444 -478 1456 -426
rect 1508 -478 1520 -426
rect 1572 -478 1584 -426
rect 1636 -478 1648 -426
rect 1700 -478 1730 -426
rect 1298 -490 1730 -478
rect 1298 -542 1328 -490
rect 1380 -542 1392 -490
rect 1444 -542 1456 -490
rect 1508 -542 1520 -490
rect 1572 -542 1584 -490
rect 1636 -542 1648 -490
rect 1700 -542 1730 -490
rect 1298 -554 1730 -542
rect 1298 -606 1328 -554
rect 1380 -606 1392 -554
rect 1444 -606 1456 -554
rect 1508 -606 1520 -554
rect 1572 -606 1584 -554
rect 1636 -606 1648 -554
rect 1700 -606 1730 -554
rect 1298 -618 1730 -606
rect 1298 -670 1328 -618
rect 1380 -670 1392 -618
rect 1444 -670 1456 -618
rect 1508 -670 1520 -618
rect 1572 -670 1584 -618
rect 1636 -670 1648 -618
rect 1700 -670 1730 -618
rect 1298 -682 1730 -670
rect 1298 -734 1328 -682
rect 1380 -734 1392 -682
rect 1444 -734 1456 -682
rect 1508 -734 1520 -682
rect 1572 -734 1584 -682
rect 1636 -734 1648 -682
rect 1700 -734 1730 -682
rect 1298 -746 1730 -734
rect 1298 -798 1328 -746
rect 1380 -798 1392 -746
rect 1444 -798 1456 -746
rect 1508 -798 1520 -746
rect 1572 -798 1584 -746
rect 1636 -798 1648 -746
rect 1700 -798 1730 -746
rect 1298 -810 1730 -798
rect 1298 -862 1328 -810
rect 1380 -862 1392 -810
rect 1444 -862 1456 -810
rect 1508 -862 1520 -810
rect 1572 -862 1584 -810
rect 1636 -862 1648 -810
rect 1700 -862 1730 -810
rect 1298 -864 1730 -862
rect 1826 -318 1896 -272
rect 1826 -352 1832 -318
rect 1866 -352 1896 -318
rect 1826 -398 1896 -352
rect 1826 -432 1832 -398
rect 1866 -432 1896 -398
rect 1826 -478 1896 -432
rect 1826 -512 1832 -478
rect 1866 -512 1896 -478
rect 1826 -558 1896 -512
rect 1826 -592 1832 -558
rect 1866 -592 1896 -558
rect 1826 -638 1896 -592
rect 1826 -672 1832 -638
rect 1866 -672 1896 -638
rect 1826 -718 1896 -672
rect 1826 -752 1832 -718
rect 1866 -752 1896 -718
rect 1826 -798 1896 -752
rect 1826 -832 1832 -798
rect 1866 -832 1896 -798
rect 0 -912 30 -878
rect 64 -912 70 -878
rect 0 -960 70 -912
rect 1826 -878 1896 -832
rect 1826 -912 1832 -878
rect 1866 -912 1896 -878
rect 1826 -960 1896 -912
rect 0 -966 1896 -960
rect 0 -1000 70 -966
rect 104 -1000 150 -966
rect 184 -1000 230 -966
rect 264 -1000 310 -966
rect 344 -1000 390 -966
rect 424 -1000 470 -966
rect 504 -1000 550 -966
rect 584 -1000 630 -966
rect 664 -1000 710 -966
rect 744 -1000 790 -966
rect 824 -1000 870 -966
rect 904 -1000 950 -966
rect 984 -1000 1030 -966
rect 1064 -1000 1110 -966
rect 1144 -1000 1190 -966
rect 1224 -1000 1270 -966
rect 1304 -1000 1350 -966
rect 1384 -1000 1430 -966
rect 1464 -1000 1510 -966
rect 1544 -1000 1590 -966
rect 1624 -1000 1670 -966
rect 1704 -1000 1750 -966
rect 1784 -1000 1896 -966
rect 0 -1030 1896 -1000
<< via1 >>
rect 184 2462 238 2514
rect 184 2382 238 2434
rect 184 2302 238 2354
rect 184 2222 238 2274
rect 184 2142 238 2194
rect 184 2062 238 2114
rect 184 1982 238 2034
rect 1414 2462 1468 2514
rect 1414 2382 1468 2434
rect 1414 2302 1468 2354
rect 1414 2222 1468 2274
rect 1414 2142 1468 2194
rect 1414 2062 1468 2114
rect 1414 1982 1468 2034
rect 2644 2462 2698 2514
rect 2644 2382 2698 2434
rect 2644 2302 2698 2354
rect 2644 2222 2698 2274
rect 2644 2142 2698 2194
rect 2644 2062 2698 2114
rect 2644 1982 2698 2034
rect 594 1850 646 1860
rect 674 1850 726 1860
rect 590 1808 646 1850
rect 670 1808 726 1850
rect 590 1798 642 1808
rect 670 1798 722 1808
rect 988 1850 1040 1860
rect 1068 1850 1120 1860
rect 984 1808 1040 1850
rect 1064 1808 1120 1850
rect 984 1798 1036 1808
rect 1064 1798 1116 1808
rect 1776 1850 1828 1860
rect 1856 1850 1908 1860
rect 1772 1808 1828 1850
rect 1852 1808 1908 1850
rect 1772 1798 1824 1808
rect 1852 1798 1904 1808
rect 2166 1798 2218 1850
rect 2246 1798 2298 1850
rect 590 1114 642 1124
rect 670 1114 722 1124
rect 590 1072 646 1114
rect 670 1072 726 1114
rect 594 1062 646 1072
rect 674 1062 726 1072
rect 984 1114 1036 1124
rect 1064 1114 1116 1124
rect 984 1072 1040 1114
rect 1064 1072 1120 1114
rect 988 1062 1040 1072
rect 1068 1062 1120 1072
rect 1772 1114 1824 1124
rect 1852 1114 1904 1124
rect 1772 1072 1828 1114
rect 1852 1072 1908 1114
rect 1776 1062 1828 1072
rect 1856 1062 1908 1072
rect 2166 1072 2218 1124
rect 2246 1072 2298 1124
rect 594 914 646 924
rect 674 914 726 924
rect 590 872 646 914
rect 670 872 726 914
rect 590 862 642 872
rect 670 862 722 872
rect 988 914 1040 924
rect 1068 914 1120 924
rect 984 872 1040 914
rect 1064 872 1120 914
rect 984 862 1036 872
rect 1064 862 1116 872
rect 1382 914 1434 924
rect 1462 914 1514 924
rect 1378 872 1434 914
rect 1458 872 1514 914
rect 1378 862 1430 872
rect 1458 862 1510 872
rect 1776 914 1828 924
rect 1856 914 1908 924
rect 1772 872 1828 914
rect 1852 872 1908 914
rect 1772 862 1824 872
rect 1852 862 1904 872
rect 2166 862 2218 914
rect 2246 862 2298 914
rect 590 122 646 174
rect 670 122 726 174
rect 984 122 1040 174
rect 1064 122 1120 174
rect 1378 128 1430 180
rect 1458 128 1510 180
rect 1772 122 1828 174
rect 1852 122 1908 174
rect 2166 122 2218 180
rect 2246 122 2298 180
rect 196 -350 248 -298
rect 260 -350 312 -298
rect 324 -350 376 -298
rect 388 -350 440 -298
rect 452 -350 504 -298
rect 516 -350 568 -298
rect 196 -414 248 -362
rect 260 -414 312 -362
rect 324 -414 376 -362
rect 388 -414 440 -362
rect 452 -414 504 -362
rect 516 -414 568 -362
rect 196 -478 248 -426
rect 260 -478 312 -426
rect 324 -478 376 -426
rect 388 -478 440 -426
rect 452 -478 504 -426
rect 516 -478 568 -426
rect 196 -542 248 -490
rect 260 -542 312 -490
rect 324 -542 376 -490
rect 388 -542 440 -490
rect 452 -542 504 -490
rect 516 -542 568 -490
rect 196 -606 248 -554
rect 260 -606 312 -554
rect 324 -606 376 -554
rect 388 -606 440 -554
rect 452 -606 504 -554
rect 516 -606 568 -554
rect 196 -670 248 -618
rect 260 -670 312 -618
rect 324 -670 376 -618
rect 388 -670 440 -618
rect 452 -670 504 -618
rect 516 -670 568 -618
rect 196 -734 248 -682
rect 260 -734 312 -682
rect 324 -734 376 -682
rect 388 -734 440 -682
rect 452 -734 504 -682
rect 516 -734 568 -682
rect 196 -798 248 -746
rect 260 -798 312 -746
rect 324 -798 376 -746
rect 388 -798 440 -746
rect 452 -798 504 -746
rect 516 -798 568 -746
rect 196 -862 248 -810
rect 260 -862 312 -810
rect 324 -862 376 -810
rect 388 -862 440 -810
rect 452 -862 504 -810
rect 516 -862 568 -810
rect 1328 -350 1380 -298
rect 1392 -350 1444 -298
rect 1456 -350 1508 -298
rect 1520 -350 1572 -298
rect 1584 -350 1636 -298
rect 1648 -350 1700 -298
rect 1328 -414 1380 -362
rect 1392 -414 1444 -362
rect 1456 -414 1508 -362
rect 1520 -414 1572 -362
rect 1584 -414 1636 -362
rect 1648 -414 1700 -362
rect 1328 -478 1380 -426
rect 1392 -478 1444 -426
rect 1456 -478 1508 -426
rect 1520 -478 1572 -426
rect 1584 -478 1636 -426
rect 1648 -478 1700 -426
rect 1328 -542 1380 -490
rect 1392 -542 1444 -490
rect 1456 -542 1508 -490
rect 1520 -542 1572 -490
rect 1584 -542 1636 -490
rect 1648 -542 1700 -490
rect 1328 -606 1380 -554
rect 1392 -606 1444 -554
rect 1456 -606 1508 -554
rect 1520 -606 1572 -554
rect 1584 -606 1636 -554
rect 1648 -606 1700 -554
rect 1328 -670 1380 -618
rect 1392 -670 1444 -618
rect 1456 -670 1508 -618
rect 1520 -670 1572 -618
rect 1584 -670 1636 -618
rect 1648 -670 1700 -618
rect 1328 -734 1380 -682
rect 1392 -734 1444 -682
rect 1456 -734 1508 -682
rect 1520 -734 1572 -682
rect 1584 -734 1636 -682
rect 1648 -734 1700 -682
rect 1328 -798 1380 -746
rect 1392 -798 1444 -746
rect 1456 -798 1508 -746
rect 1520 -798 1572 -746
rect 1584 -798 1636 -746
rect 1648 -798 1700 -746
rect 1328 -862 1380 -810
rect 1392 -862 1444 -810
rect 1456 -862 1508 -810
rect 1520 -862 1572 -810
rect 1584 -862 1636 -810
rect 1648 -862 1700 -810
<< metal2 >>
rect 172 2516 250 2550
rect 172 2460 182 2516
rect 240 2460 250 2516
rect 172 2436 250 2460
rect 172 2380 182 2436
rect 240 2380 250 2436
rect 172 2356 250 2380
rect 172 2300 182 2356
rect 240 2300 250 2356
rect 172 2276 250 2300
rect 172 2220 182 2276
rect 240 2220 250 2276
rect 172 2196 250 2220
rect 172 2140 182 2196
rect 240 2140 250 2196
rect 172 2116 250 2140
rect 172 2060 182 2116
rect 240 2060 250 2116
rect 172 2036 250 2060
rect 172 1980 182 2036
rect 240 1980 250 2036
rect 172 1950 250 1980
rect 1402 2516 1480 2550
rect 1402 2460 1412 2516
rect 1470 2460 1480 2516
rect 1402 2436 1480 2460
rect 1402 2380 1412 2436
rect 1470 2380 1480 2436
rect 1402 2356 1480 2380
rect 1402 2300 1412 2356
rect 1470 2300 1480 2356
rect 1402 2276 1480 2300
rect 1402 2220 1412 2276
rect 1470 2220 1480 2276
rect 1402 2196 1480 2220
rect 1402 2140 1412 2196
rect 1470 2140 1480 2196
rect 1402 2116 1480 2140
rect 1402 2060 1412 2116
rect 1470 2060 1480 2116
rect 1402 2036 1480 2060
rect 1402 1980 1412 2036
rect 1470 1980 1480 2036
rect 1402 1950 1480 1980
rect 2632 2516 2710 2550
rect 2632 2460 2642 2516
rect 2700 2460 2710 2516
rect 2632 2436 2710 2460
rect 2632 2380 2642 2436
rect 2700 2380 2710 2436
rect 2632 2356 2710 2380
rect 2632 2300 2642 2356
rect 2700 2300 2710 2356
rect 2632 2276 2710 2300
rect 2632 2220 2642 2276
rect 2700 2220 2710 2276
rect 2632 2196 2710 2220
rect 2632 2140 2642 2196
rect 2700 2140 2710 2196
rect 2632 2116 2710 2140
rect 2632 2060 2642 2116
rect 2700 2060 2710 2116
rect 2632 2036 2710 2060
rect 2632 1980 2642 2036
rect 2700 1980 2710 2036
rect 2632 1950 2710 1980
rect 558 1864 758 1870
rect 952 1864 1152 1870
rect 1740 1864 1940 1870
rect 554 1862 758 1864
rect 554 1850 592 1862
rect 554 1798 590 1850
rect 648 1850 672 1862
rect 648 1806 670 1850
rect 728 1806 758 1862
rect 642 1798 670 1806
rect 722 1798 758 1806
rect 948 1862 1152 1864
rect 948 1850 986 1862
rect 948 1798 984 1850
rect 1042 1850 1066 1862
rect 1042 1806 1064 1850
rect 1122 1806 1152 1862
rect 1036 1798 1064 1806
rect 1116 1798 1152 1806
rect 1736 1862 1940 1864
rect 1736 1850 1774 1862
rect 1736 1798 1772 1850
rect 1830 1850 1854 1862
rect 1830 1806 1852 1850
rect 1910 1806 1940 1862
rect 1824 1798 1852 1806
rect 1904 1798 1940 1806
rect 2130 1862 2462 1870
rect 2130 1806 2152 1862
rect 2208 1850 2236 1862
rect 2292 1850 2316 1862
rect 2218 1806 2236 1850
rect 2298 1806 2316 1850
rect 2372 1806 2396 1862
rect 2452 1806 2462 1862
rect 2130 1798 2166 1806
rect 2218 1798 2246 1806
rect 2298 1798 2462 1806
rect 542 1722 770 1736
rect 542 1666 548 1722
rect 604 1666 628 1722
rect 684 1666 708 1722
rect 764 1666 770 1722
rect 542 1642 770 1666
rect 542 1586 548 1642
rect 604 1586 628 1642
rect 684 1586 708 1642
rect 764 1586 770 1642
rect 542 1562 770 1586
rect 542 1506 548 1562
rect 604 1506 628 1562
rect 684 1506 708 1562
rect 764 1506 770 1562
rect 542 1492 770 1506
rect 936 1722 1164 1736
rect 936 1666 942 1722
rect 998 1666 1022 1722
rect 1078 1666 1102 1722
rect 1158 1666 1164 1722
rect 936 1642 1164 1666
rect 936 1586 942 1642
rect 998 1586 1022 1642
rect 1078 1586 1102 1642
rect 1158 1586 1164 1642
rect 936 1562 1164 1586
rect 936 1506 942 1562
rect 998 1506 1022 1562
rect 1078 1506 1102 1562
rect 1158 1506 1164 1562
rect 936 1492 1164 1506
rect 1724 1722 1952 1736
rect 1724 1666 1730 1722
rect 1786 1666 1810 1722
rect 1866 1666 1890 1722
rect 1946 1666 1952 1722
rect 1724 1642 1952 1666
rect 1724 1586 1730 1642
rect 1786 1586 1810 1642
rect 1866 1586 1890 1642
rect 1946 1586 1952 1642
rect 1724 1562 1952 1586
rect 1724 1506 1730 1562
rect 1786 1506 1810 1562
rect 1866 1506 1890 1562
rect 1946 1506 1952 1562
rect 1724 1492 1952 1506
rect 2118 1722 2346 1736
rect 2118 1666 2124 1722
rect 2180 1666 2204 1722
rect 2260 1666 2284 1722
rect 2340 1666 2346 1722
rect 2118 1642 2346 1666
rect 2118 1586 2124 1642
rect 2180 1586 2204 1642
rect 2260 1586 2284 1642
rect 2340 1586 2346 1642
rect 2118 1562 2346 1586
rect 2118 1506 2124 1562
rect 2180 1506 2204 1562
rect 2260 1506 2284 1562
rect 2340 1506 2346 1562
rect 2118 1492 2346 1506
rect 542 1416 770 1430
rect 542 1360 548 1416
rect 604 1360 628 1416
rect 684 1360 708 1416
rect 764 1360 770 1416
rect 542 1336 770 1360
rect 542 1280 548 1336
rect 604 1280 628 1336
rect 684 1280 708 1336
rect 764 1280 770 1336
rect 542 1256 770 1280
rect 542 1200 548 1256
rect 604 1200 628 1256
rect 684 1200 708 1256
rect 764 1200 770 1256
rect 542 1186 770 1200
rect 936 1416 1164 1430
rect 936 1360 942 1416
rect 998 1360 1022 1416
rect 1078 1360 1102 1416
rect 1158 1360 1164 1416
rect 936 1336 1164 1360
rect 936 1280 942 1336
rect 998 1280 1022 1336
rect 1078 1280 1102 1336
rect 1158 1280 1164 1336
rect 936 1256 1164 1280
rect 936 1200 942 1256
rect 998 1200 1022 1256
rect 1078 1200 1102 1256
rect 1158 1200 1164 1256
rect 936 1186 1164 1200
rect 1724 1416 1952 1430
rect 1724 1360 1730 1416
rect 1786 1360 1810 1416
rect 1866 1360 1890 1416
rect 1946 1360 1952 1416
rect 1724 1336 1952 1360
rect 1724 1280 1730 1336
rect 1786 1280 1810 1336
rect 1866 1280 1890 1336
rect 1946 1280 1952 1336
rect 1724 1256 1952 1280
rect 1724 1200 1730 1256
rect 1786 1200 1810 1256
rect 1866 1200 1890 1256
rect 1946 1200 1952 1256
rect 1724 1186 1952 1200
rect 2118 1416 2346 1430
rect 2118 1360 2124 1416
rect 2180 1360 2204 1416
rect 2260 1360 2284 1416
rect 2340 1360 2346 1416
rect 2118 1336 2346 1360
rect 2118 1280 2124 1336
rect 2180 1280 2204 1336
rect 2260 1280 2284 1336
rect 2340 1280 2346 1336
rect 2118 1256 2346 1280
rect 2118 1200 2124 1256
rect 2180 1200 2204 1256
rect 2260 1200 2284 1256
rect 2340 1200 2346 1256
rect 2118 1186 2346 1200
rect 2396 1124 2462 1798
rect 554 1072 590 1124
rect 642 1116 670 1124
rect 722 1116 758 1124
rect 554 1060 592 1072
rect 648 1072 670 1116
rect 648 1060 672 1072
rect 728 1060 758 1116
rect 554 1058 758 1060
rect 948 1072 984 1124
rect 1036 1116 1064 1124
rect 1116 1116 1152 1124
rect 948 1060 986 1072
rect 1042 1072 1064 1116
rect 1042 1060 1066 1072
rect 1122 1060 1152 1116
rect 948 1058 1152 1060
rect 1736 1072 1772 1124
rect 1824 1116 1852 1124
rect 1904 1116 1940 1124
rect 1736 1060 1774 1072
rect 1830 1072 1852 1116
rect 1830 1060 1854 1072
rect 1910 1060 1940 1116
rect 1736 1058 1940 1060
rect 558 1052 758 1058
rect 952 1052 1152 1058
rect 1740 1052 1940 1058
rect 2130 1116 2166 1124
rect 2218 1116 2246 1124
rect 2298 1116 2462 1124
rect 2130 1060 2152 1116
rect 2218 1072 2236 1116
rect 2298 1072 2316 1116
rect 2208 1060 2236 1072
rect 2292 1060 2316 1072
rect 2372 1060 2396 1116
rect 2452 1060 2462 1116
rect 2130 1052 2462 1060
rect 2396 934 2462 1052
rect 558 928 758 934
rect 952 928 1152 934
rect 1346 928 1546 934
rect 1740 928 1940 934
rect 554 926 758 928
rect 554 914 592 926
rect 554 862 590 914
rect 648 914 672 926
rect 648 870 670 914
rect 728 870 758 926
rect 642 862 670 870
rect 722 862 758 870
rect 948 926 1152 928
rect 948 914 986 926
rect 948 862 984 914
rect 1042 914 1066 926
rect 1042 870 1064 914
rect 1122 870 1152 926
rect 1036 862 1064 870
rect 1116 862 1152 870
rect 1342 926 1546 928
rect 1342 914 1380 926
rect 1342 862 1378 914
rect 1436 914 1460 926
rect 1436 870 1458 914
rect 1516 870 1546 926
rect 1430 862 1458 870
rect 1510 862 1546 870
rect 1736 926 1940 928
rect 1736 914 1774 926
rect 1736 862 1772 914
rect 1830 914 1854 926
rect 1830 870 1852 914
rect 1910 870 1940 926
rect 1824 862 1852 870
rect 1904 862 1940 870
rect 2130 926 2462 934
rect 2130 870 2152 926
rect 2208 914 2236 926
rect 2292 914 2316 926
rect 2218 870 2236 914
rect 2298 870 2316 914
rect 2372 870 2396 926
rect 2452 870 2462 926
rect 2130 862 2166 870
rect 2218 862 2246 870
rect 2298 862 2462 870
rect 542 786 770 800
rect 542 730 548 786
rect 604 730 628 786
rect 684 730 708 786
rect 764 730 770 786
rect 542 706 770 730
rect 542 650 548 706
rect 604 650 628 706
rect 684 650 708 706
rect 764 650 770 706
rect 542 626 770 650
rect 542 570 548 626
rect 604 570 628 626
rect 684 570 708 626
rect 764 570 770 626
rect 542 556 770 570
rect 936 786 1164 800
rect 936 730 942 786
rect 998 730 1022 786
rect 1078 730 1102 786
rect 1158 730 1164 786
rect 936 706 1164 730
rect 936 650 942 706
rect 998 650 1022 706
rect 1078 650 1102 706
rect 1158 650 1164 706
rect 936 626 1164 650
rect 936 570 942 626
rect 998 570 1022 626
rect 1078 570 1102 626
rect 1158 570 1164 626
rect 936 556 1164 570
rect 1330 786 1558 800
rect 1330 730 1336 786
rect 1392 730 1416 786
rect 1472 730 1496 786
rect 1552 730 1558 786
rect 1330 706 1558 730
rect 1330 650 1336 706
rect 1392 650 1416 706
rect 1472 650 1496 706
rect 1552 650 1558 706
rect 1330 626 1558 650
rect 1330 570 1336 626
rect 1392 570 1416 626
rect 1472 570 1496 626
rect 1552 570 1558 626
rect 1330 556 1558 570
rect 1724 786 1952 800
rect 1724 730 1730 786
rect 1786 730 1810 786
rect 1866 730 1890 786
rect 1946 730 1952 786
rect 1724 706 1952 730
rect 1724 650 1730 706
rect 1786 650 1810 706
rect 1866 650 1890 706
rect 1946 650 1952 706
rect 1724 626 1952 650
rect 1724 570 1730 626
rect 1786 570 1810 626
rect 1866 570 1890 626
rect 1946 570 1952 626
rect 1724 556 1952 570
rect 2118 786 2346 800
rect 2118 730 2124 786
rect 2180 730 2204 786
rect 2260 730 2284 786
rect 2340 730 2346 786
rect 2118 706 2346 730
rect 2118 650 2124 706
rect 2180 650 2204 706
rect 2260 650 2284 706
rect 2340 650 2346 706
rect 2118 626 2346 650
rect 2118 570 2124 626
rect 2180 570 2204 626
rect 2260 570 2284 626
rect 2340 570 2346 626
rect 2118 556 2346 570
rect 542 474 770 488
rect 542 418 548 474
rect 604 418 628 474
rect 684 418 708 474
rect 764 418 770 474
rect 542 394 770 418
rect 542 338 548 394
rect 604 338 628 394
rect 684 338 708 394
rect 764 338 770 394
rect 542 314 770 338
rect 542 258 548 314
rect 604 258 628 314
rect 684 258 708 314
rect 764 258 770 314
rect 542 244 770 258
rect 936 474 1164 488
rect 936 418 942 474
rect 998 418 1022 474
rect 1078 418 1102 474
rect 1158 418 1164 474
rect 936 394 1164 418
rect 936 338 942 394
rect 998 338 1022 394
rect 1078 338 1102 394
rect 1158 338 1164 394
rect 936 314 1164 338
rect 936 258 942 314
rect 998 258 1022 314
rect 1078 258 1102 314
rect 1158 258 1164 314
rect 936 244 1164 258
rect 558 176 758 184
rect 558 174 592 176
rect 648 174 672 176
rect 554 122 590 174
rect 648 122 670 174
rect 558 120 592 122
rect 648 120 672 122
rect 728 120 758 176
rect 952 176 1152 184
rect 952 174 986 176
rect 1042 174 1066 176
rect 948 122 984 174
rect 1042 122 1064 174
rect 558 112 758 120
rect 952 120 986 122
rect 1042 120 1066 122
rect 1122 120 1152 176
rect 952 112 1152 120
rect 1330 180 1558 500
rect 1724 474 1952 488
rect 1724 418 1730 474
rect 1786 418 1810 474
rect 1866 418 1890 474
rect 1946 418 1952 474
rect 1724 394 1952 418
rect 1724 338 1730 394
rect 1786 338 1810 394
rect 1866 338 1890 394
rect 1946 338 1952 394
rect 1724 314 1952 338
rect 1724 258 1730 314
rect 1786 258 1810 314
rect 1866 258 1890 314
rect 1946 258 1952 314
rect 1724 244 1952 258
rect 2118 474 2346 488
rect 2118 418 2124 474
rect 2180 418 2204 474
rect 2260 418 2284 474
rect 2340 418 2346 474
rect 2118 394 2346 418
rect 2118 338 2124 394
rect 2180 338 2204 394
rect 2260 338 2284 394
rect 2340 338 2346 394
rect 2118 314 2346 338
rect 2118 258 2124 314
rect 2180 258 2204 314
rect 2260 258 2284 314
rect 2340 258 2346 314
rect 2118 246 2346 258
rect 2118 244 2166 246
rect 2218 244 2246 246
rect 2298 244 2346 246
rect 2396 184 2462 862
rect 1330 128 1378 180
rect 1430 128 1458 180
rect 1510 128 1558 180
rect 1740 176 1940 184
rect 1740 174 1774 176
rect 1830 174 1854 176
rect 1330 34 1558 128
rect 1736 122 1772 174
rect 1830 122 1852 174
rect 1740 120 1774 122
rect 1830 120 1854 122
rect 1910 120 1940 176
rect 1740 112 1940 120
rect 2130 180 2462 184
rect 2130 176 2166 180
rect 2218 176 2246 180
rect 2298 176 2462 180
rect 2130 120 2152 176
rect 2218 122 2236 176
rect 2298 122 2316 176
rect 2208 120 2236 122
rect 2292 120 2316 122
rect 2372 120 2396 176
rect 2452 120 2462 176
rect 2130 112 2462 120
rect 2396 42 2462 112
rect 1330 -22 1336 34
rect 1392 -22 1416 34
rect 1472 -22 1496 34
rect 1552 -22 1558 34
rect 1330 -46 1558 -22
rect 1330 -102 1336 -46
rect 1392 -102 1416 -46
rect 1472 -102 1496 -46
rect 1552 -102 1558 -46
rect 1330 -126 1558 -102
rect 1330 -182 1336 -126
rect 1392 -182 1416 -126
rect 1472 -182 1496 -126
rect 1552 -182 1558 -126
rect 1330 -192 1558 -182
rect 2388 34 2468 42
rect 2388 -22 2400 34
rect 2456 -22 2468 34
rect 2388 -46 2468 -22
rect 2388 -102 2400 -46
rect 2456 -102 2468 -46
rect 2388 -126 2468 -102
rect 2388 -182 2400 -126
rect 2456 -182 2468 -126
rect 2388 -192 2468 -182
rect 166 -298 598 -294
rect 166 -310 196 -298
rect 248 -310 260 -298
rect 312 -310 324 -298
rect 376 -310 388 -298
rect 440 -310 452 -298
rect 504 -310 516 -298
rect 568 -310 598 -298
rect 166 -366 194 -310
rect 250 -350 260 -310
rect 504 -350 514 -310
rect 250 -362 274 -350
rect 330 -362 354 -350
rect 410 -362 434 -350
rect 490 -362 514 -350
rect 250 -366 260 -362
rect 504 -366 514 -362
rect 570 -366 598 -310
rect 166 -390 196 -366
rect 248 -390 260 -366
rect 312 -390 324 -366
rect 376 -390 388 -366
rect 440 -390 452 -366
rect 504 -390 516 -366
rect 568 -390 598 -366
rect 166 -446 194 -390
rect 250 -414 260 -390
rect 504 -414 514 -390
rect 250 -426 274 -414
rect 330 -426 354 -414
rect 410 -426 434 -414
rect 490 -426 514 -414
rect 250 -446 260 -426
rect 504 -446 514 -426
rect 570 -446 598 -390
rect 166 -470 196 -446
rect 248 -470 260 -446
rect 312 -470 324 -446
rect 376 -470 388 -446
rect 440 -470 452 -446
rect 504 -470 516 -446
rect 568 -470 598 -446
rect 166 -526 194 -470
rect 250 -478 260 -470
rect 504 -478 514 -470
rect 250 -490 274 -478
rect 330 -490 354 -478
rect 410 -490 434 -478
rect 490 -490 514 -478
rect 250 -526 260 -490
rect 504 -526 514 -490
rect 570 -526 598 -470
rect 166 -542 196 -526
rect 248 -542 260 -526
rect 312 -542 324 -526
rect 376 -542 388 -526
rect 440 -542 452 -526
rect 504 -542 516 -526
rect 568 -542 598 -526
rect 166 -550 598 -542
rect 166 -606 194 -550
rect 250 -554 274 -550
rect 330 -554 354 -550
rect 410 -554 434 -550
rect 490 -554 514 -550
rect 250 -606 260 -554
rect 504 -606 514 -554
rect 570 -606 598 -550
rect 166 -618 598 -606
rect 166 -630 196 -618
rect 248 -630 260 -618
rect 312 -630 324 -618
rect 376 -630 388 -618
rect 440 -630 452 -618
rect 504 -630 516 -618
rect 568 -630 598 -618
rect 166 -686 194 -630
rect 250 -670 260 -630
rect 504 -670 514 -630
rect 250 -682 274 -670
rect 330 -682 354 -670
rect 410 -682 434 -670
rect 490 -682 514 -670
rect 250 -686 260 -682
rect 504 -686 514 -682
rect 570 -686 598 -630
rect 166 -710 196 -686
rect 248 -710 260 -686
rect 312 -710 324 -686
rect 376 -710 388 -686
rect 440 -710 452 -686
rect 504 -710 516 -686
rect 568 -710 598 -686
rect 166 -766 194 -710
rect 250 -734 260 -710
rect 504 -734 514 -710
rect 250 -746 274 -734
rect 330 -746 354 -734
rect 410 -746 434 -734
rect 490 -746 514 -734
rect 250 -766 260 -746
rect 504 -766 514 -746
rect 570 -766 598 -710
rect 166 -790 196 -766
rect 248 -790 260 -766
rect 312 -790 324 -766
rect 376 -790 388 -766
rect 440 -790 452 -766
rect 504 -790 516 -766
rect 568 -790 598 -766
rect 166 -846 194 -790
rect 250 -798 260 -790
rect 504 -798 514 -790
rect 250 -810 274 -798
rect 330 -810 354 -798
rect 410 -810 434 -798
rect 490 -810 514 -798
rect 250 -846 260 -810
rect 504 -846 514 -810
rect 570 -846 598 -790
rect 166 -862 196 -846
rect 248 -862 260 -846
rect 312 -862 324 -846
rect 376 -862 388 -846
rect 440 -862 452 -846
rect 504 -862 516 -846
rect 568 -862 598 -846
rect 166 -864 598 -862
rect 1298 -298 1730 -294
rect 1298 -310 1328 -298
rect 1380 -310 1392 -298
rect 1444 -310 1456 -298
rect 1508 -310 1520 -298
rect 1572 -310 1584 -298
rect 1636 -310 1648 -298
rect 1700 -310 1730 -298
rect 1298 -366 1326 -310
rect 1382 -350 1392 -310
rect 1636 -350 1646 -310
rect 1382 -362 1406 -350
rect 1462 -362 1486 -350
rect 1542 -362 1566 -350
rect 1622 -362 1646 -350
rect 1382 -366 1392 -362
rect 1636 -366 1646 -362
rect 1702 -366 1730 -310
rect 1298 -390 1328 -366
rect 1380 -390 1392 -366
rect 1444 -390 1456 -366
rect 1508 -390 1520 -366
rect 1572 -390 1584 -366
rect 1636 -390 1648 -366
rect 1700 -390 1730 -366
rect 1298 -446 1326 -390
rect 1382 -414 1392 -390
rect 1636 -414 1646 -390
rect 1382 -426 1406 -414
rect 1462 -426 1486 -414
rect 1542 -426 1566 -414
rect 1622 -426 1646 -414
rect 1382 -446 1392 -426
rect 1636 -446 1646 -426
rect 1702 -446 1730 -390
rect 1298 -470 1328 -446
rect 1380 -470 1392 -446
rect 1444 -470 1456 -446
rect 1508 -470 1520 -446
rect 1572 -470 1584 -446
rect 1636 -470 1648 -446
rect 1700 -470 1730 -446
rect 1298 -526 1326 -470
rect 1382 -478 1392 -470
rect 1636 -478 1646 -470
rect 1382 -490 1406 -478
rect 1462 -490 1486 -478
rect 1542 -490 1566 -478
rect 1622 -490 1646 -478
rect 1382 -526 1392 -490
rect 1636 -526 1646 -490
rect 1702 -526 1730 -470
rect 1298 -542 1328 -526
rect 1380 -542 1392 -526
rect 1444 -542 1456 -526
rect 1508 -542 1520 -526
rect 1572 -542 1584 -526
rect 1636 -542 1648 -526
rect 1700 -542 1730 -526
rect 1298 -550 1730 -542
rect 1298 -606 1326 -550
rect 1382 -554 1406 -550
rect 1462 -554 1486 -550
rect 1542 -554 1566 -550
rect 1622 -554 1646 -550
rect 1382 -606 1392 -554
rect 1636 -606 1646 -554
rect 1702 -606 1730 -550
rect 1298 -618 1730 -606
rect 1298 -630 1328 -618
rect 1380 -630 1392 -618
rect 1444 -630 1456 -618
rect 1508 -630 1520 -618
rect 1572 -630 1584 -618
rect 1636 -630 1648 -618
rect 1700 -630 1730 -618
rect 1298 -686 1326 -630
rect 1382 -670 1392 -630
rect 1636 -670 1646 -630
rect 1382 -682 1406 -670
rect 1462 -682 1486 -670
rect 1542 -682 1566 -670
rect 1622 -682 1646 -670
rect 1382 -686 1392 -682
rect 1636 -686 1646 -682
rect 1702 -686 1730 -630
rect 1298 -710 1328 -686
rect 1380 -710 1392 -686
rect 1444 -710 1456 -686
rect 1508 -710 1520 -686
rect 1572 -710 1584 -686
rect 1636 -710 1648 -686
rect 1700 -710 1730 -686
rect 1298 -766 1326 -710
rect 1382 -734 1392 -710
rect 1636 -734 1646 -710
rect 1382 -746 1406 -734
rect 1462 -746 1486 -734
rect 1542 -746 1566 -734
rect 1622 -746 1646 -734
rect 1382 -766 1392 -746
rect 1636 -766 1646 -746
rect 1702 -766 1730 -710
rect 1298 -790 1328 -766
rect 1380 -790 1392 -766
rect 1444 -790 1456 -766
rect 1508 -790 1520 -766
rect 1572 -790 1584 -766
rect 1636 -790 1648 -766
rect 1700 -790 1730 -766
rect 1298 -846 1326 -790
rect 1382 -798 1392 -790
rect 1636 -798 1646 -790
rect 1382 -810 1406 -798
rect 1462 -810 1486 -798
rect 1542 -810 1566 -798
rect 1622 -810 1646 -798
rect 1382 -846 1392 -810
rect 1636 -846 1646 -810
rect 1702 -846 1730 -790
rect 1298 -862 1328 -846
rect 1380 -862 1392 -846
rect 1444 -862 1456 -846
rect 1508 -862 1520 -846
rect 1572 -862 1584 -846
rect 1636 -862 1648 -846
rect 1700 -862 1730 -846
rect 1298 -864 1730 -862
<< via2 >>
rect 182 2514 240 2516
rect 182 2462 184 2514
rect 184 2462 238 2514
rect 238 2462 240 2514
rect 182 2460 240 2462
rect 182 2434 240 2436
rect 182 2382 184 2434
rect 184 2382 238 2434
rect 238 2382 240 2434
rect 182 2380 240 2382
rect 182 2354 240 2356
rect 182 2302 184 2354
rect 184 2302 238 2354
rect 238 2302 240 2354
rect 182 2300 240 2302
rect 182 2274 240 2276
rect 182 2222 184 2274
rect 184 2222 238 2274
rect 238 2222 240 2274
rect 182 2220 240 2222
rect 182 2194 240 2196
rect 182 2142 184 2194
rect 184 2142 238 2194
rect 238 2142 240 2194
rect 182 2140 240 2142
rect 182 2114 240 2116
rect 182 2062 184 2114
rect 184 2062 238 2114
rect 238 2062 240 2114
rect 182 2060 240 2062
rect 182 2034 240 2036
rect 182 1982 184 2034
rect 184 1982 238 2034
rect 238 1982 240 2034
rect 182 1980 240 1982
rect 1412 2514 1470 2516
rect 1412 2462 1414 2514
rect 1414 2462 1468 2514
rect 1468 2462 1470 2514
rect 1412 2460 1470 2462
rect 1412 2434 1470 2436
rect 1412 2382 1414 2434
rect 1414 2382 1468 2434
rect 1468 2382 1470 2434
rect 1412 2380 1470 2382
rect 1412 2354 1470 2356
rect 1412 2302 1414 2354
rect 1414 2302 1468 2354
rect 1468 2302 1470 2354
rect 1412 2300 1470 2302
rect 1412 2274 1470 2276
rect 1412 2222 1414 2274
rect 1414 2222 1468 2274
rect 1468 2222 1470 2274
rect 1412 2220 1470 2222
rect 1412 2194 1470 2196
rect 1412 2142 1414 2194
rect 1414 2142 1468 2194
rect 1468 2142 1470 2194
rect 1412 2140 1470 2142
rect 1412 2114 1470 2116
rect 1412 2062 1414 2114
rect 1414 2062 1468 2114
rect 1468 2062 1470 2114
rect 1412 2060 1470 2062
rect 1412 2034 1470 2036
rect 1412 1982 1414 2034
rect 1414 1982 1468 2034
rect 1468 1982 1470 2034
rect 1412 1980 1470 1982
rect 2642 2514 2700 2516
rect 2642 2462 2644 2514
rect 2644 2462 2698 2514
rect 2698 2462 2700 2514
rect 2642 2460 2700 2462
rect 2642 2434 2700 2436
rect 2642 2382 2644 2434
rect 2644 2382 2698 2434
rect 2698 2382 2700 2434
rect 2642 2380 2700 2382
rect 2642 2354 2700 2356
rect 2642 2302 2644 2354
rect 2644 2302 2698 2354
rect 2698 2302 2700 2354
rect 2642 2300 2700 2302
rect 2642 2274 2700 2276
rect 2642 2222 2644 2274
rect 2644 2222 2698 2274
rect 2698 2222 2700 2274
rect 2642 2220 2700 2222
rect 2642 2194 2700 2196
rect 2642 2142 2644 2194
rect 2644 2142 2698 2194
rect 2698 2142 2700 2194
rect 2642 2140 2700 2142
rect 2642 2114 2700 2116
rect 2642 2062 2644 2114
rect 2644 2062 2698 2114
rect 2698 2062 2700 2114
rect 2642 2060 2700 2062
rect 2642 2034 2700 2036
rect 2642 1982 2644 2034
rect 2644 1982 2698 2034
rect 2698 1982 2700 2034
rect 2642 1980 2700 1982
rect 592 1860 648 1862
rect 592 1850 594 1860
rect 594 1850 646 1860
rect 592 1808 646 1850
rect 646 1808 648 1860
rect 672 1860 728 1862
rect 672 1850 674 1860
rect 674 1850 726 1860
rect 592 1806 642 1808
rect 642 1806 648 1808
rect 672 1808 726 1850
rect 726 1808 728 1860
rect 672 1806 722 1808
rect 722 1806 728 1808
rect 986 1860 1042 1862
rect 986 1850 988 1860
rect 988 1850 1040 1860
rect 986 1808 1040 1850
rect 1040 1808 1042 1860
rect 1066 1860 1122 1862
rect 1066 1850 1068 1860
rect 1068 1850 1120 1860
rect 986 1806 1036 1808
rect 1036 1806 1042 1808
rect 1066 1808 1120 1850
rect 1120 1808 1122 1860
rect 1066 1806 1116 1808
rect 1116 1806 1122 1808
rect 1774 1860 1830 1862
rect 1774 1850 1776 1860
rect 1776 1850 1828 1860
rect 1774 1808 1828 1850
rect 1828 1808 1830 1860
rect 1854 1860 1910 1862
rect 1854 1850 1856 1860
rect 1856 1850 1908 1860
rect 1774 1806 1824 1808
rect 1824 1806 1830 1808
rect 1854 1808 1908 1850
rect 1908 1808 1910 1860
rect 1854 1806 1904 1808
rect 1904 1806 1910 1808
rect 2152 1850 2208 1862
rect 2236 1850 2292 1862
rect 2152 1806 2166 1850
rect 2166 1806 2208 1850
rect 2236 1806 2246 1850
rect 2246 1806 2292 1850
rect 2316 1806 2372 1862
rect 2396 1806 2452 1862
rect 548 1666 604 1722
rect 628 1666 684 1722
rect 708 1666 764 1722
rect 548 1586 604 1642
rect 628 1586 684 1642
rect 708 1586 764 1642
rect 548 1506 604 1562
rect 628 1506 684 1562
rect 708 1506 764 1562
rect 942 1666 998 1722
rect 1022 1666 1078 1722
rect 1102 1666 1158 1722
rect 942 1586 998 1642
rect 1022 1586 1078 1642
rect 1102 1586 1158 1642
rect 942 1506 998 1562
rect 1022 1506 1078 1562
rect 1102 1506 1158 1562
rect 1730 1666 1786 1722
rect 1810 1666 1866 1722
rect 1890 1666 1946 1722
rect 1730 1586 1786 1642
rect 1810 1586 1866 1642
rect 1890 1586 1946 1642
rect 1730 1506 1786 1562
rect 1810 1506 1866 1562
rect 1890 1506 1946 1562
rect 2124 1666 2180 1722
rect 2204 1666 2260 1722
rect 2284 1666 2340 1722
rect 2124 1586 2180 1642
rect 2204 1586 2260 1642
rect 2284 1586 2340 1642
rect 2124 1506 2180 1562
rect 2204 1506 2260 1562
rect 2284 1506 2340 1562
rect 548 1360 604 1416
rect 628 1360 684 1416
rect 708 1360 764 1416
rect 548 1280 604 1336
rect 628 1280 684 1336
rect 708 1280 764 1336
rect 548 1200 604 1256
rect 628 1200 684 1256
rect 708 1200 764 1256
rect 942 1360 998 1416
rect 1022 1360 1078 1416
rect 1102 1360 1158 1416
rect 942 1280 998 1336
rect 1022 1280 1078 1336
rect 1102 1280 1158 1336
rect 942 1200 998 1256
rect 1022 1200 1078 1256
rect 1102 1200 1158 1256
rect 1730 1360 1786 1416
rect 1810 1360 1866 1416
rect 1890 1360 1946 1416
rect 1730 1280 1786 1336
rect 1810 1280 1866 1336
rect 1890 1280 1946 1336
rect 1730 1200 1786 1256
rect 1810 1200 1866 1256
rect 1890 1200 1946 1256
rect 2124 1360 2180 1416
rect 2204 1360 2260 1416
rect 2284 1360 2340 1416
rect 2124 1280 2180 1336
rect 2204 1280 2260 1336
rect 2284 1280 2340 1336
rect 2124 1200 2180 1256
rect 2204 1200 2260 1256
rect 2284 1200 2340 1256
rect 592 1114 642 1116
rect 642 1114 648 1116
rect 592 1072 646 1114
rect 592 1062 594 1072
rect 594 1062 646 1072
rect 646 1062 648 1114
rect 672 1114 722 1116
rect 722 1114 728 1116
rect 672 1072 726 1114
rect 592 1060 648 1062
rect 672 1062 674 1072
rect 674 1062 726 1072
rect 726 1062 728 1114
rect 672 1060 728 1062
rect 986 1114 1036 1116
rect 1036 1114 1042 1116
rect 986 1072 1040 1114
rect 986 1062 988 1072
rect 988 1062 1040 1072
rect 1040 1062 1042 1114
rect 1066 1114 1116 1116
rect 1116 1114 1122 1116
rect 1066 1072 1120 1114
rect 986 1060 1042 1062
rect 1066 1062 1068 1072
rect 1068 1062 1120 1072
rect 1120 1062 1122 1114
rect 1066 1060 1122 1062
rect 1774 1114 1824 1116
rect 1824 1114 1830 1116
rect 1774 1072 1828 1114
rect 1774 1062 1776 1072
rect 1776 1062 1828 1072
rect 1828 1062 1830 1114
rect 1854 1114 1904 1116
rect 1904 1114 1910 1116
rect 1854 1072 1908 1114
rect 1774 1060 1830 1062
rect 1854 1062 1856 1072
rect 1856 1062 1908 1072
rect 1908 1062 1910 1114
rect 1854 1060 1910 1062
rect 2152 1072 2166 1116
rect 2166 1072 2208 1116
rect 2236 1072 2246 1116
rect 2246 1072 2292 1116
rect 2152 1060 2208 1072
rect 2236 1060 2292 1072
rect 2316 1060 2372 1116
rect 2396 1060 2452 1116
rect 592 924 648 926
rect 592 914 594 924
rect 594 914 646 924
rect 592 872 646 914
rect 646 872 648 924
rect 672 924 728 926
rect 672 914 674 924
rect 674 914 726 924
rect 592 870 642 872
rect 642 870 648 872
rect 672 872 726 914
rect 726 872 728 924
rect 672 870 722 872
rect 722 870 728 872
rect 986 924 1042 926
rect 986 914 988 924
rect 988 914 1040 924
rect 986 872 1040 914
rect 1040 872 1042 924
rect 1066 924 1122 926
rect 1066 914 1068 924
rect 1068 914 1120 924
rect 986 870 1036 872
rect 1036 870 1042 872
rect 1066 872 1120 914
rect 1120 872 1122 924
rect 1066 870 1116 872
rect 1116 870 1122 872
rect 1380 924 1436 926
rect 1380 914 1382 924
rect 1382 914 1434 924
rect 1380 872 1434 914
rect 1434 872 1436 924
rect 1460 924 1516 926
rect 1460 914 1462 924
rect 1462 914 1514 924
rect 1380 870 1430 872
rect 1430 870 1436 872
rect 1460 872 1514 914
rect 1514 872 1516 924
rect 1460 870 1510 872
rect 1510 870 1516 872
rect 1774 924 1830 926
rect 1774 914 1776 924
rect 1776 914 1828 924
rect 1774 872 1828 914
rect 1828 872 1830 924
rect 1854 924 1910 926
rect 1854 914 1856 924
rect 1856 914 1908 924
rect 1774 870 1824 872
rect 1824 870 1830 872
rect 1854 872 1908 914
rect 1908 872 1910 924
rect 1854 870 1904 872
rect 1904 870 1910 872
rect 2152 914 2208 926
rect 2236 914 2292 926
rect 2152 870 2166 914
rect 2166 870 2208 914
rect 2236 870 2246 914
rect 2246 870 2292 914
rect 2316 870 2372 926
rect 2396 870 2452 926
rect 548 730 604 786
rect 628 730 684 786
rect 708 730 764 786
rect 548 650 604 706
rect 628 650 684 706
rect 708 650 764 706
rect 548 570 604 626
rect 628 570 684 626
rect 708 570 764 626
rect 942 730 998 786
rect 1022 730 1078 786
rect 1102 730 1158 786
rect 942 650 998 706
rect 1022 650 1078 706
rect 1102 650 1158 706
rect 942 570 998 626
rect 1022 570 1078 626
rect 1102 570 1158 626
rect 1336 730 1392 786
rect 1416 730 1472 786
rect 1496 730 1552 786
rect 1336 650 1392 706
rect 1416 650 1472 706
rect 1496 650 1552 706
rect 1336 570 1392 626
rect 1416 570 1472 626
rect 1496 570 1552 626
rect 1730 730 1786 786
rect 1810 730 1866 786
rect 1890 730 1946 786
rect 1730 650 1786 706
rect 1810 650 1866 706
rect 1890 650 1946 706
rect 1730 570 1786 626
rect 1810 570 1866 626
rect 1890 570 1946 626
rect 2124 730 2180 786
rect 2204 730 2260 786
rect 2284 730 2340 786
rect 2124 650 2180 706
rect 2204 650 2260 706
rect 2284 650 2340 706
rect 2124 570 2180 626
rect 2204 570 2260 626
rect 2284 570 2340 626
rect 548 418 604 474
rect 628 418 684 474
rect 708 418 764 474
rect 548 338 604 394
rect 628 338 684 394
rect 708 338 764 394
rect 548 258 604 314
rect 628 258 684 314
rect 708 258 764 314
rect 942 418 998 474
rect 1022 418 1078 474
rect 1102 418 1158 474
rect 942 338 998 394
rect 1022 338 1078 394
rect 1102 338 1158 394
rect 942 258 998 314
rect 1022 258 1078 314
rect 1102 258 1158 314
rect 592 174 648 176
rect 672 174 728 176
rect 592 122 646 174
rect 646 122 648 174
rect 672 122 726 174
rect 726 122 728 174
rect 592 120 648 122
rect 672 120 728 122
rect 986 174 1042 176
rect 1066 174 1122 176
rect 986 122 1040 174
rect 1040 122 1042 174
rect 1066 122 1120 174
rect 1120 122 1122 174
rect 986 120 1042 122
rect 1066 120 1122 122
rect 1730 418 1786 474
rect 1810 418 1866 474
rect 1890 418 1946 474
rect 1730 338 1786 394
rect 1810 338 1866 394
rect 1890 338 1946 394
rect 1730 258 1786 314
rect 1810 258 1866 314
rect 1890 258 1946 314
rect 2124 418 2180 474
rect 2204 418 2260 474
rect 2284 418 2340 474
rect 2124 338 2180 394
rect 2204 338 2260 394
rect 2284 338 2340 394
rect 2124 258 2180 314
rect 2204 258 2260 314
rect 2284 258 2340 314
rect 1774 174 1830 176
rect 1854 174 1910 176
rect 1774 122 1828 174
rect 1828 122 1830 174
rect 1854 122 1908 174
rect 1908 122 1910 174
rect 1774 120 1830 122
rect 1854 120 1910 122
rect 2152 122 2166 176
rect 2166 122 2208 176
rect 2236 122 2246 176
rect 2246 122 2292 176
rect 2152 120 2208 122
rect 2236 120 2292 122
rect 2316 120 2372 176
rect 2396 120 2452 176
rect 1336 -22 1392 34
rect 1416 -22 1472 34
rect 1496 -22 1552 34
rect 1336 -102 1392 -46
rect 1416 -102 1472 -46
rect 1496 -102 1552 -46
rect 1336 -182 1392 -126
rect 1416 -182 1472 -126
rect 1496 -182 1552 -126
rect 2400 -22 2456 34
rect 2400 -102 2456 -46
rect 2400 -182 2456 -126
rect 194 -350 196 -310
rect 196 -350 248 -310
rect 248 -350 250 -310
rect 274 -350 312 -310
rect 312 -350 324 -310
rect 324 -350 330 -310
rect 354 -350 376 -310
rect 376 -350 388 -310
rect 388 -350 410 -310
rect 434 -350 440 -310
rect 440 -350 452 -310
rect 452 -350 490 -310
rect 514 -350 516 -310
rect 516 -350 568 -310
rect 568 -350 570 -310
rect 194 -362 250 -350
rect 274 -362 330 -350
rect 354 -362 410 -350
rect 434 -362 490 -350
rect 514 -362 570 -350
rect 194 -366 196 -362
rect 196 -366 248 -362
rect 248 -366 250 -362
rect 274 -366 312 -362
rect 312 -366 324 -362
rect 324 -366 330 -362
rect 354 -366 376 -362
rect 376 -366 388 -362
rect 388 -366 410 -362
rect 434 -366 440 -362
rect 440 -366 452 -362
rect 452 -366 490 -362
rect 514 -366 516 -362
rect 516 -366 568 -362
rect 568 -366 570 -362
rect 194 -414 196 -390
rect 196 -414 248 -390
rect 248 -414 250 -390
rect 274 -414 312 -390
rect 312 -414 324 -390
rect 324 -414 330 -390
rect 354 -414 376 -390
rect 376 -414 388 -390
rect 388 -414 410 -390
rect 434 -414 440 -390
rect 440 -414 452 -390
rect 452 -414 490 -390
rect 514 -414 516 -390
rect 516 -414 568 -390
rect 568 -414 570 -390
rect 194 -426 250 -414
rect 274 -426 330 -414
rect 354 -426 410 -414
rect 434 -426 490 -414
rect 514 -426 570 -414
rect 194 -446 196 -426
rect 196 -446 248 -426
rect 248 -446 250 -426
rect 274 -446 312 -426
rect 312 -446 324 -426
rect 324 -446 330 -426
rect 354 -446 376 -426
rect 376 -446 388 -426
rect 388 -446 410 -426
rect 434 -446 440 -426
rect 440 -446 452 -426
rect 452 -446 490 -426
rect 514 -446 516 -426
rect 516 -446 568 -426
rect 568 -446 570 -426
rect 194 -478 196 -470
rect 196 -478 248 -470
rect 248 -478 250 -470
rect 274 -478 312 -470
rect 312 -478 324 -470
rect 324 -478 330 -470
rect 354 -478 376 -470
rect 376 -478 388 -470
rect 388 -478 410 -470
rect 434 -478 440 -470
rect 440 -478 452 -470
rect 452 -478 490 -470
rect 514 -478 516 -470
rect 516 -478 568 -470
rect 568 -478 570 -470
rect 194 -490 250 -478
rect 274 -490 330 -478
rect 354 -490 410 -478
rect 434 -490 490 -478
rect 514 -490 570 -478
rect 194 -526 196 -490
rect 196 -526 248 -490
rect 248 -526 250 -490
rect 274 -526 312 -490
rect 312 -526 324 -490
rect 324 -526 330 -490
rect 354 -526 376 -490
rect 376 -526 388 -490
rect 388 -526 410 -490
rect 434 -526 440 -490
rect 440 -526 452 -490
rect 452 -526 490 -490
rect 514 -526 516 -490
rect 516 -526 568 -490
rect 568 -526 570 -490
rect 194 -554 250 -550
rect 274 -554 330 -550
rect 354 -554 410 -550
rect 434 -554 490 -550
rect 514 -554 570 -550
rect 194 -606 196 -554
rect 196 -606 248 -554
rect 248 -606 250 -554
rect 274 -606 312 -554
rect 312 -606 324 -554
rect 324 -606 330 -554
rect 354 -606 376 -554
rect 376 -606 388 -554
rect 388 -606 410 -554
rect 434 -606 440 -554
rect 440 -606 452 -554
rect 452 -606 490 -554
rect 514 -606 516 -554
rect 516 -606 568 -554
rect 568 -606 570 -554
rect 194 -670 196 -630
rect 196 -670 248 -630
rect 248 -670 250 -630
rect 274 -670 312 -630
rect 312 -670 324 -630
rect 324 -670 330 -630
rect 354 -670 376 -630
rect 376 -670 388 -630
rect 388 -670 410 -630
rect 434 -670 440 -630
rect 440 -670 452 -630
rect 452 -670 490 -630
rect 514 -670 516 -630
rect 516 -670 568 -630
rect 568 -670 570 -630
rect 194 -682 250 -670
rect 274 -682 330 -670
rect 354 -682 410 -670
rect 434 -682 490 -670
rect 514 -682 570 -670
rect 194 -686 196 -682
rect 196 -686 248 -682
rect 248 -686 250 -682
rect 274 -686 312 -682
rect 312 -686 324 -682
rect 324 -686 330 -682
rect 354 -686 376 -682
rect 376 -686 388 -682
rect 388 -686 410 -682
rect 434 -686 440 -682
rect 440 -686 452 -682
rect 452 -686 490 -682
rect 514 -686 516 -682
rect 516 -686 568 -682
rect 568 -686 570 -682
rect 194 -734 196 -710
rect 196 -734 248 -710
rect 248 -734 250 -710
rect 274 -734 312 -710
rect 312 -734 324 -710
rect 324 -734 330 -710
rect 354 -734 376 -710
rect 376 -734 388 -710
rect 388 -734 410 -710
rect 434 -734 440 -710
rect 440 -734 452 -710
rect 452 -734 490 -710
rect 514 -734 516 -710
rect 516 -734 568 -710
rect 568 -734 570 -710
rect 194 -746 250 -734
rect 274 -746 330 -734
rect 354 -746 410 -734
rect 434 -746 490 -734
rect 514 -746 570 -734
rect 194 -766 196 -746
rect 196 -766 248 -746
rect 248 -766 250 -746
rect 274 -766 312 -746
rect 312 -766 324 -746
rect 324 -766 330 -746
rect 354 -766 376 -746
rect 376 -766 388 -746
rect 388 -766 410 -746
rect 434 -766 440 -746
rect 440 -766 452 -746
rect 452 -766 490 -746
rect 514 -766 516 -746
rect 516 -766 568 -746
rect 568 -766 570 -746
rect 194 -798 196 -790
rect 196 -798 248 -790
rect 248 -798 250 -790
rect 274 -798 312 -790
rect 312 -798 324 -790
rect 324 -798 330 -790
rect 354 -798 376 -790
rect 376 -798 388 -790
rect 388 -798 410 -790
rect 434 -798 440 -790
rect 440 -798 452 -790
rect 452 -798 490 -790
rect 514 -798 516 -790
rect 516 -798 568 -790
rect 568 -798 570 -790
rect 194 -810 250 -798
rect 274 -810 330 -798
rect 354 -810 410 -798
rect 434 -810 490 -798
rect 514 -810 570 -798
rect 194 -846 196 -810
rect 196 -846 248 -810
rect 248 -846 250 -810
rect 274 -846 312 -810
rect 312 -846 324 -810
rect 324 -846 330 -810
rect 354 -846 376 -810
rect 376 -846 388 -810
rect 388 -846 410 -810
rect 434 -846 440 -810
rect 440 -846 452 -810
rect 452 -846 490 -810
rect 514 -846 516 -810
rect 516 -846 568 -810
rect 568 -846 570 -810
rect 1326 -350 1328 -310
rect 1328 -350 1380 -310
rect 1380 -350 1382 -310
rect 1406 -350 1444 -310
rect 1444 -350 1456 -310
rect 1456 -350 1462 -310
rect 1486 -350 1508 -310
rect 1508 -350 1520 -310
rect 1520 -350 1542 -310
rect 1566 -350 1572 -310
rect 1572 -350 1584 -310
rect 1584 -350 1622 -310
rect 1646 -350 1648 -310
rect 1648 -350 1700 -310
rect 1700 -350 1702 -310
rect 1326 -362 1382 -350
rect 1406 -362 1462 -350
rect 1486 -362 1542 -350
rect 1566 -362 1622 -350
rect 1646 -362 1702 -350
rect 1326 -366 1328 -362
rect 1328 -366 1380 -362
rect 1380 -366 1382 -362
rect 1406 -366 1444 -362
rect 1444 -366 1456 -362
rect 1456 -366 1462 -362
rect 1486 -366 1508 -362
rect 1508 -366 1520 -362
rect 1520 -366 1542 -362
rect 1566 -366 1572 -362
rect 1572 -366 1584 -362
rect 1584 -366 1622 -362
rect 1646 -366 1648 -362
rect 1648 -366 1700 -362
rect 1700 -366 1702 -362
rect 1326 -414 1328 -390
rect 1328 -414 1380 -390
rect 1380 -414 1382 -390
rect 1406 -414 1444 -390
rect 1444 -414 1456 -390
rect 1456 -414 1462 -390
rect 1486 -414 1508 -390
rect 1508 -414 1520 -390
rect 1520 -414 1542 -390
rect 1566 -414 1572 -390
rect 1572 -414 1584 -390
rect 1584 -414 1622 -390
rect 1646 -414 1648 -390
rect 1648 -414 1700 -390
rect 1700 -414 1702 -390
rect 1326 -426 1382 -414
rect 1406 -426 1462 -414
rect 1486 -426 1542 -414
rect 1566 -426 1622 -414
rect 1646 -426 1702 -414
rect 1326 -446 1328 -426
rect 1328 -446 1380 -426
rect 1380 -446 1382 -426
rect 1406 -446 1444 -426
rect 1444 -446 1456 -426
rect 1456 -446 1462 -426
rect 1486 -446 1508 -426
rect 1508 -446 1520 -426
rect 1520 -446 1542 -426
rect 1566 -446 1572 -426
rect 1572 -446 1584 -426
rect 1584 -446 1622 -426
rect 1646 -446 1648 -426
rect 1648 -446 1700 -426
rect 1700 -446 1702 -426
rect 1326 -478 1328 -470
rect 1328 -478 1380 -470
rect 1380 -478 1382 -470
rect 1406 -478 1444 -470
rect 1444 -478 1456 -470
rect 1456 -478 1462 -470
rect 1486 -478 1508 -470
rect 1508 -478 1520 -470
rect 1520 -478 1542 -470
rect 1566 -478 1572 -470
rect 1572 -478 1584 -470
rect 1584 -478 1622 -470
rect 1646 -478 1648 -470
rect 1648 -478 1700 -470
rect 1700 -478 1702 -470
rect 1326 -490 1382 -478
rect 1406 -490 1462 -478
rect 1486 -490 1542 -478
rect 1566 -490 1622 -478
rect 1646 -490 1702 -478
rect 1326 -526 1328 -490
rect 1328 -526 1380 -490
rect 1380 -526 1382 -490
rect 1406 -526 1444 -490
rect 1444 -526 1456 -490
rect 1456 -526 1462 -490
rect 1486 -526 1508 -490
rect 1508 -526 1520 -490
rect 1520 -526 1542 -490
rect 1566 -526 1572 -490
rect 1572 -526 1584 -490
rect 1584 -526 1622 -490
rect 1646 -526 1648 -490
rect 1648 -526 1700 -490
rect 1700 -526 1702 -490
rect 1326 -554 1382 -550
rect 1406 -554 1462 -550
rect 1486 -554 1542 -550
rect 1566 -554 1622 -550
rect 1646 -554 1702 -550
rect 1326 -606 1328 -554
rect 1328 -606 1380 -554
rect 1380 -606 1382 -554
rect 1406 -606 1444 -554
rect 1444 -606 1456 -554
rect 1456 -606 1462 -554
rect 1486 -606 1508 -554
rect 1508 -606 1520 -554
rect 1520 -606 1542 -554
rect 1566 -606 1572 -554
rect 1572 -606 1584 -554
rect 1584 -606 1622 -554
rect 1646 -606 1648 -554
rect 1648 -606 1700 -554
rect 1700 -606 1702 -554
rect 1326 -670 1328 -630
rect 1328 -670 1380 -630
rect 1380 -670 1382 -630
rect 1406 -670 1444 -630
rect 1444 -670 1456 -630
rect 1456 -670 1462 -630
rect 1486 -670 1508 -630
rect 1508 -670 1520 -630
rect 1520 -670 1542 -630
rect 1566 -670 1572 -630
rect 1572 -670 1584 -630
rect 1584 -670 1622 -630
rect 1646 -670 1648 -630
rect 1648 -670 1700 -630
rect 1700 -670 1702 -630
rect 1326 -682 1382 -670
rect 1406 -682 1462 -670
rect 1486 -682 1542 -670
rect 1566 -682 1622 -670
rect 1646 -682 1702 -670
rect 1326 -686 1328 -682
rect 1328 -686 1380 -682
rect 1380 -686 1382 -682
rect 1406 -686 1444 -682
rect 1444 -686 1456 -682
rect 1456 -686 1462 -682
rect 1486 -686 1508 -682
rect 1508 -686 1520 -682
rect 1520 -686 1542 -682
rect 1566 -686 1572 -682
rect 1572 -686 1584 -682
rect 1584 -686 1622 -682
rect 1646 -686 1648 -682
rect 1648 -686 1700 -682
rect 1700 -686 1702 -682
rect 1326 -734 1328 -710
rect 1328 -734 1380 -710
rect 1380 -734 1382 -710
rect 1406 -734 1444 -710
rect 1444 -734 1456 -710
rect 1456 -734 1462 -710
rect 1486 -734 1508 -710
rect 1508 -734 1520 -710
rect 1520 -734 1542 -710
rect 1566 -734 1572 -710
rect 1572 -734 1584 -710
rect 1584 -734 1622 -710
rect 1646 -734 1648 -710
rect 1648 -734 1700 -710
rect 1700 -734 1702 -710
rect 1326 -746 1382 -734
rect 1406 -746 1462 -734
rect 1486 -746 1542 -734
rect 1566 -746 1622 -734
rect 1646 -746 1702 -734
rect 1326 -766 1328 -746
rect 1328 -766 1380 -746
rect 1380 -766 1382 -746
rect 1406 -766 1444 -746
rect 1444 -766 1456 -746
rect 1456 -766 1462 -746
rect 1486 -766 1508 -746
rect 1508 -766 1520 -746
rect 1520 -766 1542 -746
rect 1566 -766 1572 -746
rect 1572 -766 1584 -746
rect 1584 -766 1622 -746
rect 1646 -766 1648 -746
rect 1648 -766 1700 -746
rect 1700 -766 1702 -746
rect 1326 -798 1328 -790
rect 1328 -798 1380 -790
rect 1380 -798 1382 -790
rect 1406 -798 1444 -790
rect 1444 -798 1456 -790
rect 1456 -798 1462 -790
rect 1486 -798 1508 -790
rect 1508 -798 1520 -790
rect 1520 -798 1542 -790
rect 1566 -798 1572 -790
rect 1572 -798 1584 -790
rect 1584 -798 1622 -790
rect 1646 -798 1648 -790
rect 1648 -798 1700 -790
rect 1700 -798 1702 -790
rect 1326 -810 1382 -798
rect 1406 -810 1462 -798
rect 1486 -810 1542 -798
rect 1566 -810 1622 -798
rect 1646 -810 1702 -798
rect 1326 -846 1328 -810
rect 1328 -846 1380 -810
rect 1380 -846 1382 -810
rect 1406 -846 1444 -810
rect 1444 -846 1456 -810
rect 1456 -846 1462 -810
rect 1486 -846 1508 -810
rect 1508 -846 1520 -810
rect 1520 -846 1542 -810
rect 1566 -846 1572 -810
rect 1572 -846 1584 -810
rect 1584 -846 1622 -810
rect 1646 -846 1648 -810
rect 1648 -846 1700 -810
rect 1700 -846 1702 -810
<< metal3 >>
rect 172 2520 250 2550
rect 172 2456 178 2520
rect 244 2456 250 2520
rect 172 2440 250 2456
rect 172 2376 178 2440
rect 244 2376 250 2440
rect 172 2360 250 2376
rect 172 2296 178 2360
rect 244 2296 250 2360
rect 172 2280 250 2296
rect 172 2216 178 2280
rect 244 2216 250 2280
rect 172 2200 250 2216
rect 172 2136 178 2200
rect 244 2136 250 2200
rect 172 2120 250 2136
rect 172 2056 178 2120
rect 244 2056 250 2120
rect 172 2040 250 2056
rect 172 1976 178 2040
rect 244 1976 250 2040
rect 172 1950 250 1976
rect 1402 2520 1480 2550
rect 1402 2456 1408 2520
rect 1474 2456 1480 2520
rect 1402 2440 1480 2456
rect 1402 2376 1408 2440
rect 1474 2376 1480 2440
rect 1402 2360 1480 2376
rect 1402 2296 1408 2360
rect 1474 2296 1480 2360
rect 1402 2280 1480 2296
rect 1402 2216 1408 2280
rect 1474 2216 1480 2280
rect 1402 2200 1480 2216
rect 1402 2136 1408 2200
rect 1474 2136 1480 2200
rect 1402 2120 1480 2136
rect 1402 2056 1408 2120
rect 1474 2056 1480 2120
rect 1402 2040 1480 2056
rect 1402 1976 1408 2040
rect 1474 1976 1480 2040
rect 1402 1950 1480 1976
rect 2632 2520 2710 2550
rect 2632 2456 2638 2520
rect 2704 2456 2710 2520
rect 2632 2440 2710 2456
rect 2632 2376 2638 2440
rect 2704 2376 2710 2440
rect 2632 2360 2710 2376
rect 2632 2296 2638 2360
rect 2704 2296 2710 2360
rect 2632 2280 2710 2296
rect 2632 2216 2638 2280
rect 2704 2216 2710 2280
rect 2632 2200 2710 2216
rect 2632 2136 2638 2200
rect 2704 2136 2710 2200
rect 2632 2120 2710 2136
rect 2632 2056 2638 2120
rect 2704 2056 2710 2120
rect 2632 2040 2710 2056
rect 2632 1976 2638 2040
rect 2704 1976 2710 2040
rect 2632 1950 2710 1976
rect 558 1864 758 1870
rect 952 1864 1152 1870
rect 1740 1864 1940 1870
rect 2130 1864 2462 1870
rect 554 1862 2462 1864
rect 554 1806 592 1862
rect 648 1806 672 1862
rect 728 1806 986 1862
rect 1042 1806 1066 1862
rect 1122 1806 1774 1862
rect 1830 1806 1854 1862
rect 1910 1806 2152 1862
rect 2208 1806 2236 1862
rect 2292 1806 2316 1862
rect 2372 1806 2396 1862
rect 2452 1806 2462 1862
rect 554 1798 2462 1806
rect 148 1726 2346 1736
rect 148 1662 158 1726
rect 222 1662 238 1726
rect 302 1662 318 1726
rect 382 1722 2346 1726
rect 382 1666 548 1722
rect 604 1666 628 1722
rect 684 1666 708 1722
rect 764 1666 942 1722
rect 998 1666 1022 1722
rect 1078 1666 1102 1722
rect 1158 1666 1730 1722
rect 1786 1666 1810 1722
rect 1866 1666 1890 1722
rect 1946 1666 2124 1722
rect 2180 1666 2204 1722
rect 2260 1666 2284 1722
rect 2340 1666 2346 1722
rect 382 1662 2346 1666
rect 148 1646 2346 1662
rect 148 1582 158 1646
rect 222 1582 238 1646
rect 302 1582 318 1646
rect 382 1642 2346 1646
rect 382 1586 548 1642
rect 604 1586 628 1642
rect 684 1586 708 1642
rect 764 1586 942 1642
rect 998 1586 1022 1642
rect 1078 1586 1102 1642
rect 1158 1586 1730 1642
rect 1786 1586 1810 1642
rect 1866 1586 1890 1642
rect 1946 1586 2124 1642
rect 2180 1586 2204 1642
rect 2260 1586 2284 1642
rect 2340 1586 2346 1642
rect 382 1582 2346 1586
rect 148 1566 2346 1582
rect 148 1502 158 1566
rect 222 1502 238 1566
rect 302 1502 318 1566
rect 382 1562 2346 1566
rect 382 1506 548 1562
rect 604 1506 628 1562
rect 684 1506 708 1562
rect 764 1506 942 1562
rect 998 1506 1022 1562
rect 1078 1506 1102 1562
rect 1158 1506 1730 1562
rect 1786 1506 1810 1562
rect 1866 1506 1890 1562
rect 1946 1506 2124 1562
rect 2180 1506 2204 1562
rect 2260 1506 2284 1562
rect 2340 1506 2346 1562
rect 382 1502 2346 1506
rect 148 1492 2346 1502
rect 542 1420 2740 1430
rect 542 1416 2506 1420
rect 542 1360 548 1416
rect 604 1360 628 1416
rect 684 1360 708 1416
rect 764 1360 942 1416
rect 998 1360 1022 1416
rect 1078 1360 1102 1416
rect 1158 1360 1730 1416
rect 1786 1360 1810 1416
rect 1866 1360 1890 1416
rect 1946 1360 2124 1416
rect 2180 1360 2204 1416
rect 2260 1360 2284 1416
rect 2340 1360 2506 1416
rect 542 1356 2506 1360
rect 2570 1356 2586 1420
rect 2650 1356 2666 1420
rect 2730 1356 2740 1420
rect 542 1340 2740 1356
rect 542 1336 2506 1340
rect 542 1280 548 1336
rect 604 1280 628 1336
rect 684 1280 708 1336
rect 764 1280 942 1336
rect 998 1280 1022 1336
rect 1078 1280 1102 1336
rect 1158 1280 1730 1336
rect 1786 1280 1810 1336
rect 1866 1280 1890 1336
rect 1946 1280 2124 1336
rect 2180 1280 2204 1336
rect 2260 1280 2284 1336
rect 2340 1280 2506 1336
rect 542 1276 2506 1280
rect 2570 1276 2586 1340
rect 2650 1276 2666 1340
rect 2730 1276 2740 1340
rect 542 1260 2740 1276
rect 542 1256 2506 1260
rect 542 1200 548 1256
rect 604 1200 628 1256
rect 684 1200 708 1256
rect 764 1200 942 1256
rect 998 1200 1022 1256
rect 1078 1200 1102 1256
rect 1158 1200 1730 1256
rect 1786 1200 1810 1256
rect 1866 1200 1890 1256
rect 1946 1200 2124 1256
rect 2180 1200 2204 1256
rect 2260 1200 2284 1256
rect 2340 1200 2506 1256
rect 542 1196 2506 1200
rect 2570 1196 2586 1260
rect 2650 1196 2666 1260
rect 2730 1196 2740 1260
rect 542 1186 2740 1196
rect 554 1116 2462 1124
rect 554 1060 592 1116
rect 648 1060 672 1116
rect 728 1060 986 1116
rect 1042 1060 1066 1116
rect 1122 1060 1774 1116
rect 1830 1060 1854 1116
rect 1910 1060 2152 1116
rect 2208 1060 2236 1116
rect 2292 1060 2316 1116
rect 2372 1060 2396 1116
rect 2452 1060 2462 1116
rect 554 1058 2462 1060
rect 558 1052 758 1058
rect 952 1052 1152 1058
rect 1740 1052 1940 1058
rect 2130 1052 2462 1058
rect 558 928 758 934
rect 952 928 1152 934
rect 1346 928 1546 934
rect 1740 928 1940 934
rect 2130 928 2462 934
rect 554 926 2462 928
rect 554 870 592 926
rect 648 870 672 926
rect 728 870 986 926
rect 1042 870 1066 926
rect 1122 870 1380 926
rect 1436 870 1460 926
rect 1516 870 1774 926
rect 1830 870 1854 926
rect 1910 870 2152 926
rect 2208 870 2236 926
rect 2292 870 2316 926
rect 2372 870 2396 926
rect 2452 870 2462 926
rect 554 862 2462 870
rect 148 790 2346 800
rect 148 726 158 790
rect 222 726 238 790
rect 302 726 318 790
rect 382 786 2346 790
rect 382 730 548 786
rect 604 730 628 786
rect 684 730 708 786
rect 764 730 942 786
rect 998 730 1022 786
rect 1078 730 1102 786
rect 1158 730 1336 786
rect 1392 730 1416 786
rect 1472 730 1496 786
rect 1552 730 1730 786
rect 1786 730 1810 786
rect 1866 730 1890 786
rect 1946 730 2124 786
rect 2180 730 2204 786
rect 2260 730 2284 786
rect 2340 730 2346 786
rect 382 726 2346 730
rect 148 710 2346 726
rect 148 646 158 710
rect 222 646 238 710
rect 302 646 318 710
rect 382 706 2346 710
rect 382 650 548 706
rect 604 650 628 706
rect 684 650 708 706
rect 764 650 942 706
rect 998 650 1022 706
rect 1078 650 1102 706
rect 1158 650 1336 706
rect 1392 650 1416 706
rect 1472 650 1496 706
rect 1552 650 1730 706
rect 1786 650 1810 706
rect 1866 650 1890 706
rect 1946 650 2124 706
rect 2180 650 2204 706
rect 2260 650 2284 706
rect 2340 650 2346 706
rect 382 646 2346 650
rect 148 630 2346 646
rect 148 566 158 630
rect 222 566 238 630
rect 302 566 318 630
rect 382 626 2346 630
rect 382 570 548 626
rect 604 570 628 626
rect 684 570 708 626
rect 764 570 942 626
rect 998 570 1022 626
rect 1078 570 1102 626
rect 1158 570 1336 626
rect 1392 570 1416 626
rect 1472 570 1496 626
rect 1552 570 1730 626
rect 1786 570 1810 626
rect 1866 570 1890 626
rect 1946 570 2124 626
rect 2180 570 2204 626
rect 2260 570 2284 626
rect 2340 570 2346 626
rect 382 566 2346 570
rect 148 556 2346 566
rect 542 478 2740 488
rect 542 474 2506 478
rect 542 418 548 474
rect 604 418 628 474
rect 684 418 708 474
rect 764 418 942 474
rect 998 418 1022 474
rect 1078 418 1102 474
rect 1158 418 1730 474
rect 1786 418 1810 474
rect 1866 418 1890 474
rect 1946 418 2124 474
rect 2180 418 2204 474
rect 2260 418 2284 474
rect 2340 418 2506 474
rect 542 414 2506 418
rect 2570 414 2586 478
rect 2650 414 2666 478
rect 2730 414 2740 478
rect 542 398 2740 414
rect 542 394 2506 398
rect 542 338 548 394
rect 604 338 628 394
rect 684 338 708 394
rect 764 338 942 394
rect 998 338 1022 394
rect 1078 338 1102 394
rect 1158 338 1730 394
rect 1786 338 1810 394
rect 1866 338 1890 394
rect 1946 338 2124 394
rect 2180 338 2204 394
rect 2260 338 2284 394
rect 2340 338 2506 394
rect 542 334 2506 338
rect 2570 334 2586 398
rect 2650 334 2666 398
rect 2730 334 2740 398
rect 542 318 2740 334
rect 542 314 2506 318
rect 542 258 548 314
rect 604 258 628 314
rect 684 258 708 314
rect 764 258 942 314
rect 998 258 1022 314
rect 1078 258 1102 314
rect 1158 258 1730 314
rect 1786 258 1810 314
rect 1866 258 1890 314
rect 1946 258 2124 314
rect 2180 258 2204 314
rect 2260 258 2284 314
rect 2340 258 2506 314
rect 542 254 2506 258
rect 2570 254 2586 318
rect 2650 254 2666 318
rect 2730 254 2740 318
rect 542 244 2740 254
rect 554 176 2462 184
rect 554 120 592 176
rect 648 120 672 176
rect 728 120 986 176
rect 1042 120 1066 176
rect 1122 120 1774 176
rect 1830 120 1854 176
rect 1910 120 2152 176
rect 2208 120 2236 176
rect 2292 120 2316 176
rect 2372 120 2396 176
rect 2452 120 2462 176
rect 554 118 2462 120
rect 558 112 758 118
rect 952 112 1152 118
rect 1740 112 1940 118
rect 2130 112 2462 118
rect 1298 36 1730 48
rect 2388 36 2468 42
rect 1298 34 2468 36
rect 1298 -22 1336 34
rect 1392 -22 1416 34
rect 1472 -22 1496 34
rect 1552 -22 2400 34
rect 2456 -22 2468 34
rect 1298 -46 2468 -22
rect 1298 -102 1336 -46
rect 1392 -102 1416 -46
rect 1472 -102 1496 -46
rect 1552 -102 2400 -46
rect 2456 -102 2468 -46
rect 1298 -126 2468 -102
rect 1298 -182 1336 -126
rect 1392 -182 1416 -126
rect 1472 -182 1496 -126
rect 1552 -182 2400 -126
rect 2456 -182 2468 -126
rect 1298 -192 2468 -182
rect 0 -310 598 -294
rect 0 -366 194 -310
rect 250 -366 274 -310
rect 330 -366 354 -310
rect 410 -366 434 -310
rect 490 -366 514 -310
rect 570 -366 598 -310
rect 0 -390 598 -366
rect 0 -446 194 -390
rect 250 -446 274 -390
rect 330 -446 354 -390
rect 410 -446 434 -390
rect 490 -446 514 -390
rect 570 -446 598 -390
rect 0 -470 598 -446
rect 0 -526 194 -470
rect 250 -526 274 -470
rect 330 -526 354 -470
rect 410 -526 434 -470
rect 490 -526 514 -470
rect 570 -526 598 -470
rect 0 -550 598 -526
rect 0 -606 194 -550
rect 250 -606 274 -550
rect 330 -606 354 -550
rect 410 -606 434 -550
rect 490 -606 514 -550
rect 570 -606 598 -550
rect 0 -630 598 -606
rect 0 -686 194 -630
rect 250 -686 274 -630
rect 330 -686 354 -630
rect 410 -686 434 -630
rect 490 -686 514 -630
rect 570 -686 598 -630
rect 0 -710 598 -686
rect 0 -766 194 -710
rect 250 -766 274 -710
rect 330 -766 354 -710
rect 410 -766 434 -710
rect 490 -766 514 -710
rect 570 -766 598 -710
rect 0 -790 598 -766
rect 0 -846 194 -790
rect 250 -846 274 -790
rect 330 -846 354 -790
rect 410 -846 434 -790
rect 490 -846 514 -790
rect 570 -846 598 -790
rect 0 -864 598 -846
rect 1298 -310 1730 -192
rect 1298 -366 1326 -310
rect 1382 -366 1406 -310
rect 1462 -366 1486 -310
rect 1542 -366 1566 -310
rect 1622 -366 1646 -310
rect 1702 -366 1730 -310
rect 1298 -390 1730 -366
rect 1298 -446 1326 -390
rect 1382 -446 1406 -390
rect 1462 -446 1486 -390
rect 1542 -446 1566 -390
rect 1622 -446 1646 -390
rect 1702 -446 1730 -390
rect 1298 -470 1730 -446
rect 1298 -526 1326 -470
rect 1382 -526 1406 -470
rect 1462 -526 1486 -470
rect 1542 -526 1566 -470
rect 1622 -526 1646 -470
rect 1702 -526 1730 -470
rect 1298 -550 1730 -526
rect 1298 -606 1326 -550
rect 1382 -606 1406 -550
rect 1462 -606 1486 -550
rect 1542 -606 1566 -550
rect 1622 -606 1646 -550
rect 1702 -606 1730 -550
rect 1298 -630 1730 -606
rect 1298 -686 1326 -630
rect 1382 -686 1406 -630
rect 1462 -686 1486 -630
rect 1542 -686 1566 -630
rect 1622 -686 1646 -630
rect 1702 -686 1730 -630
rect 1298 -710 1730 -686
rect 1298 -766 1326 -710
rect 1382 -766 1406 -710
rect 1462 -766 1486 -710
rect 1542 -766 1566 -710
rect 1622 -766 1646 -710
rect 1702 -766 1730 -710
rect 1298 -790 1730 -766
rect 1298 -846 1326 -790
rect 1382 -846 1406 -790
rect 1462 -846 1486 -790
rect 1542 -846 1566 -790
rect 1622 -846 1646 -790
rect 1702 -846 1730 -790
rect 1298 -864 1730 -846
<< via3 >>
rect 178 2516 244 2520
rect 178 2460 182 2516
rect 182 2460 240 2516
rect 240 2460 244 2516
rect 178 2456 244 2460
rect 178 2436 244 2440
rect 178 2380 182 2436
rect 182 2380 240 2436
rect 240 2380 244 2436
rect 178 2376 244 2380
rect 178 2356 244 2360
rect 178 2300 182 2356
rect 182 2300 240 2356
rect 240 2300 244 2356
rect 178 2296 244 2300
rect 178 2276 244 2280
rect 178 2220 182 2276
rect 182 2220 240 2276
rect 240 2220 244 2276
rect 178 2216 244 2220
rect 178 2196 244 2200
rect 178 2140 182 2196
rect 182 2140 240 2196
rect 240 2140 244 2196
rect 178 2136 244 2140
rect 178 2116 244 2120
rect 178 2060 182 2116
rect 182 2060 240 2116
rect 240 2060 244 2116
rect 178 2056 244 2060
rect 178 2036 244 2040
rect 178 1980 182 2036
rect 182 1980 240 2036
rect 240 1980 244 2036
rect 178 1976 244 1980
rect 1408 2516 1474 2520
rect 1408 2460 1412 2516
rect 1412 2460 1470 2516
rect 1470 2460 1474 2516
rect 1408 2456 1474 2460
rect 1408 2436 1474 2440
rect 1408 2380 1412 2436
rect 1412 2380 1470 2436
rect 1470 2380 1474 2436
rect 1408 2376 1474 2380
rect 1408 2356 1474 2360
rect 1408 2300 1412 2356
rect 1412 2300 1470 2356
rect 1470 2300 1474 2356
rect 1408 2296 1474 2300
rect 1408 2276 1474 2280
rect 1408 2220 1412 2276
rect 1412 2220 1470 2276
rect 1470 2220 1474 2276
rect 1408 2216 1474 2220
rect 1408 2196 1474 2200
rect 1408 2140 1412 2196
rect 1412 2140 1470 2196
rect 1470 2140 1474 2196
rect 1408 2136 1474 2140
rect 1408 2116 1474 2120
rect 1408 2060 1412 2116
rect 1412 2060 1470 2116
rect 1470 2060 1474 2116
rect 1408 2056 1474 2060
rect 1408 2036 1474 2040
rect 1408 1980 1412 2036
rect 1412 1980 1470 2036
rect 1470 1980 1474 2036
rect 1408 1976 1474 1980
rect 2638 2516 2704 2520
rect 2638 2460 2642 2516
rect 2642 2460 2700 2516
rect 2700 2460 2704 2516
rect 2638 2456 2704 2460
rect 2638 2436 2704 2440
rect 2638 2380 2642 2436
rect 2642 2380 2700 2436
rect 2700 2380 2704 2436
rect 2638 2376 2704 2380
rect 2638 2356 2704 2360
rect 2638 2300 2642 2356
rect 2642 2300 2700 2356
rect 2700 2300 2704 2356
rect 2638 2296 2704 2300
rect 2638 2276 2704 2280
rect 2638 2220 2642 2276
rect 2642 2220 2700 2276
rect 2700 2220 2704 2276
rect 2638 2216 2704 2220
rect 2638 2196 2704 2200
rect 2638 2140 2642 2196
rect 2642 2140 2700 2196
rect 2700 2140 2704 2196
rect 2638 2136 2704 2140
rect 2638 2116 2704 2120
rect 2638 2060 2642 2116
rect 2642 2060 2700 2116
rect 2700 2060 2704 2116
rect 2638 2056 2704 2060
rect 2638 2036 2704 2040
rect 2638 1980 2642 2036
rect 2642 1980 2700 2036
rect 2700 1980 2704 2036
rect 2638 1976 2704 1980
rect 158 1662 222 1726
rect 238 1662 302 1726
rect 318 1662 382 1726
rect 158 1582 222 1646
rect 238 1582 302 1646
rect 318 1582 382 1646
rect 158 1502 222 1566
rect 238 1502 302 1566
rect 318 1502 382 1566
rect 2506 1356 2570 1420
rect 2586 1356 2650 1420
rect 2666 1356 2730 1420
rect 2506 1276 2570 1340
rect 2586 1276 2650 1340
rect 2666 1276 2730 1340
rect 2506 1196 2570 1260
rect 2586 1196 2650 1260
rect 2666 1196 2730 1260
rect 158 726 222 790
rect 238 726 302 790
rect 318 726 382 790
rect 158 646 222 710
rect 238 646 302 710
rect 318 646 382 710
rect 158 566 222 630
rect 238 566 302 630
rect 318 566 382 630
rect 2506 414 2570 478
rect 2586 414 2650 478
rect 2666 414 2730 478
rect 2506 334 2570 398
rect 2586 334 2650 398
rect 2666 334 2730 398
rect 2506 254 2570 318
rect 2586 254 2650 318
rect 2666 254 2730 318
<< metal4 >>
rect 36 2526 392 2550
rect 36 2290 94 2526
rect 330 2290 392 2526
rect 36 2280 392 2290
rect 36 2216 178 2280
rect 244 2216 392 2280
rect 36 2206 392 2216
rect 36 1970 94 2206
rect 330 1970 392 2206
rect 36 1946 392 1970
rect 1266 2526 1622 2550
rect 1266 2290 1324 2526
rect 1560 2290 1622 2526
rect 1266 2280 1622 2290
rect 1266 2216 1408 2280
rect 1474 2216 1622 2280
rect 1266 2206 1622 2216
rect 1266 1970 1324 2206
rect 1560 1970 1622 2206
rect 1266 1946 1622 1970
rect 2496 2526 2852 2550
rect 2496 2290 2554 2526
rect 2790 2290 2852 2526
rect 2496 2280 2852 2290
rect 2496 2216 2638 2280
rect 2704 2216 2852 2280
rect 2496 2206 2852 2216
rect 2496 1970 2554 2206
rect 2790 1970 2852 2206
rect 2496 1946 2852 1970
rect 148 1726 392 1946
rect 148 1662 158 1726
rect 222 1662 238 1726
rect 302 1662 318 1726
rect 382 1662 392 1726
rect 148 1646 392 1662
rect 148 1582 158 1646
rect 222 1582 238 1646
rect 302 1582 318 1646
rect 382 1582 392 1646
rect 148 1566 392 1582
rect 148 1502 158 1566
rect 222 1502 238 1566
rect 302 1502 318 1566
rect 382 1502 392 1566
rect 148 790 392 1502
rect 148 726 158 790
rect 222 726 238 790
rect 302 726 318 790
rect 382 726 392 790
rect 148 710 392 726
rect 148 646 158 710
rect 222 646 238 710
rect 302 646 318 710
rect 382 646 392 710
rect 148 630 392 646
rect 148 566 158 630
rect 222 566 238 630
rect 302 566 318 630
rect 382 566 392 630
rect 148 556 392 566
rect 2496 1420 2740 1430
rect 2496 1356 2506 1420
rect 2570 1356 2586 1420
rect 2650 1356 2666 1420
rect 2730 1356 2740 1420
rect 2496 1340 2740 1356
rect 2496 1276 2506 1340
rect 2570 1276 2586 1340
rect 2650 1276 2666 1340
rect 2730 1276 2740 1340
rect 2496 1260 2740 1276
rect 2496 1196 2506 1260
rect 2570 1196 2586 1260
rect 2650 1196 2666 1260
rect 2730 1196 2740 1260
rect 2496 478 2740 1196
rect 2496 414 2506 478
rect 2570 414 2586 478
rect 2650 414 2666 478
rect 2730 414 2740 478
rect 2496 398 2740 414
rect 2496 334 2506 398
rect 2570 334 2586 398
rect 2650 334 2666 398
rect 2730 334 2740 398
rect 2496 318 2740 334
rect 2496 254 2506 318
rect 2570 254 2586 318
rect 2650 254 2666 318
rect 2730 254 2740 318
rect 2496 -192 2740 254
<< via4 >>
rect 94 2520 330 2526
rect 94 2456 178 2520
rect 178 2456 244 2520
rect 244 2456 330 2520
rect 94 2440 330 2456
rect 94 2376 178 2440
rect 178 2376 244 2440
rect 244 2376 330 2440
rect 94 2360 330 2376
rect 94 2296 178 2360
rect 178 2296 244 2360
rect 244 2296 330 2360
rect 94 2290 330 2296
rect 94 2200 330 2206
rect 94 2136 178 2200
rect 178 2136 244 2200
rect 244 2136 330 2200
rect 94 2120 330 2136
rect 94 2056 178 2120
rect 178 2056 244 2120
rect 244 2056 330 2120
rect 94 2040 330 2056
rect 94 1976 178 2040
rect 178 1976 244 2040
rect 244 1976 330 2040
rect 94 1970 330 1976
rect 1324 2520 1560 2526
rect 1324 2456 1408 2520
rect 1408 2456 1474 2520
rect 1474 2456 1560 2520
rect 1324 2440 1560 2456
rect 1324 2376 1408 2440
rect 1408 2376 1474 2440
rect 1474 2376 1560 2440
rect 1324 2360 1560 2376
rect 1324 2296 1408 2360
rect 1408 2296 1474 2360
rect 1474 2296 1560 2360
rect 1324 2290 1560 2296
rect 1324 2200 1560 2206
rect 1324 2136 1408 2200
rect 1408 2136 1474 2200
rect 1474 2136 1560 2200
rect 1324 2120 1560 2136
rect 1324 2056 1408 2120
rect 1408 2056 1474 2120
rect 1474 2056 1560 2120
rect 1324 2040 1560 2056
rect 1324 1976 1408 2040
rect 1408 1976 1474 2040
rect 1474 1976 1560 2040
rect 1324 1970 1560 1976
rect 2554 2520 2790 2526
rect 2554 2456 2638 2520
rect 2638 2456 2704 2520
rect 2704 2456 2790 2520
rect 2554 2440 2790 2456
rect 2554 2376 2638 2440
rect 2638 2376 2704 2440
rect 2704 2376 2790 2440
rect 2554 2360 2790 2376
rect 2554 2296 2638 2360
rect 2638 2296 2704 2360
rect 2704 2296 2790 2360
rect 2554 2290 2790 2296
rect 2554 2200 2790 2206
rect 2554 2136 2638 2200
rect 2638 2136 2704 2200
rect 2704 2136 2790 2200
rect 2554 2120 2790 2136
rect 2554 2056 2638 2120
rect 2638 2056 2704 2120
rect 2704 2056 2790 2120
rect 2554 2040 2790 2056
rect 2554 1976 2638 2040
rect 2638 1976 2704 2040
rect 2704 1976 2790 2040
rect 2554 1970 2790 1976
<< metal5 >>
rect 36 2526 2852 2550
rect 36 2290 94 2526
rect 330 2290 1324 2526
rect 1560 2290 2554 2526
rect 2790 2290 2852 2526
rect 36 2206 2852 2290
rect 36 1970 94 2206
rect 330 1970 1324 2206
rect 1560 1970 2554 2206
rect 2790 1970 2852 2206
rect 36 1950 2852 1970
rect 36 1946 392 1950
rect 1266 1946 1622 1950
rect 2496 1946 2852 1950
use sky130_fd_pr__res_high_po_2p85_5ZUK6C  sky130_fd_pr__res_high_po_2p85_5ZUK6C_0
timestamp 1654612214
transform 0 1 948 -1 0 -579
box -451 -948 451 948
use vco_pmirr_base  vco_pmirr_base_0
timestamp 1654600796
transform -1 0 3018 0 1 1058
box 130 -1058 3018 928
<< labels >>
flabel metal4 s 2574 -176 2628 -156 0 FreeSans 800 0 0 0 IND_CT
port 0 nsew
flabel metal5 s 60 2228 74 2266 0 FreeSans 800 0 0 0 VDD
port 2 nsew
flabel metal3 s 12 -594 26 -556 0 FreeSans 800 0 0 0 VBIAS
port 1 nsew
flabel metal1 s 1838 -1014 1884 -992 0 FreeSans 800 0 0 0 GND
port 3 nsew
<< end >>
