** sch_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/capbank.sch
.subckt capbank VDD GND bit0 bit1 bit2 bit3 bit4 bit5 OUT_P OUT_N
*.iopin VDD
*.iopin GND
*.ipin bit0
*.ipin bit1
*.ipin bit2
*.ipin bit3
*.ipin bit4
*.ipin bit5
*.iopin OUT_P
*.iopin OUT_N
X1 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X2 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X3 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X4 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X5 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X6 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X7 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X8 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X9 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X10 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X11 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X12 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X13 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X14 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X15 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X16 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X17 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X18 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X19 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X20 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X21 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X22 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X23 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X24 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X25 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X26 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X27 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X28 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X29 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X30 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X31 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X32 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X33 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X34 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X35 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X36 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X37 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X38 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X39 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X40 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X41 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X42 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X43 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X44 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X45 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X46 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X47 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X48 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X49 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X50 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X51 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X52 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X53 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X54 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X55 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X56 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X57 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X58 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X59 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X60 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X61 w_inv1 bit1 OUT_P GND OUT_N cell_unit
X62 w_inv1 bit1 OUT_P GND OUT_N cell_unit
X63 w_inv0 bit0 OUT_P GND OUT_N cell_unit
X64 bit0 w_inv0 VDD GND inv
X65 bit1 w_inv1 VDD GND inv
X66 bit2 w_inv2 VDD GND inv
X67 bit3 w_inv3 VDD GND inv
X68 bit4 w_inv4 VDD GND inv
X69 bit5 w_inv5 VDD GND inv
.ends

* expanding   symbol:  cell_unit.sym # of pins=5
** sym_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/cell_unit.sym
** sch_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/cell_unit.sch
.subckt cell_unit  V_bias ON OUT_N GND OUT_P
*.iopin OUT_N
*.iopin OUT_P
*.iopin GND
*.ipin ON
*.ipin V_bias
XC1 OUT_N net1 sky130_fd_pr__cap_mim_m3_1 W=3.3 L=3.3 MF=1 m=1
XC2 OUT_P net2 sky130_fd_pr__cap_mim_m3_1 W=3.3 L=3.3 MF=1 m=1
XR1 net1 V_bias GND sky130_fd_pr__res_xhigh_po_0p35 L=1.5 mult=1 m=1
XR2 net2 V_bias GND sky130_fd_pr__res_xhigh_po_0p35 L=1.5 mult=1 m=1
X1 net2 ON net1 GND sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15
.ends


* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/inv.sym
** sch_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/inv.sch
.subckt inv  IN OUT VDD GND
*.ipin IN
*.opin OUT
*.iopin VDD
*.iopin GND
XM1 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15.sym # of pins=4
** sym_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15.sym
** sch_path: /home/asic/Desktop/ASIC_ONE/magic_workdir/VCO_xshem/sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15.sch
.subckt sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15  DRAIN GATE SOURCE SUBSTRATE
*.iopin SOURCE
*.iopin DRAIN
*.ipin GATE
*.ipin SUBSTRATE
**** begin user architecture code


X0 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 w=1.65e+06u l=150000u
X1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 w=1.65e+06u l=150000u


**** end user architecture code
.ends

.end
