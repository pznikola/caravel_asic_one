magic
tech sky130B
timestamp 1654600796
<< nwell >>
rect 65 23 1509 464
rect 65 6 89 23
rect 106 6 286 23
rect 303 6 483 23
rect 500 6 680 23
rect 697 6 877 23
rect 894 6 1074 23
rect 1091 6 1271 23
rect 1288 6 1468 23
rect 1485 6 1509 23
rect 65 -529 1509 6
<< nsubdiff >>
rect 83 440 1491 446
rect 83 423 106 440
rect 123 423 146 440
rect 163 423 186 440
rect 203 423 226 440
rect 243 423 266 440
rect 283 423 306 440
rect 323 423 346 440
rect 363 423 386 440
rect 403 423 426 440
rect 443 423 466 440
rect 483 423 506 440
rect 523 423 546 440
rect 563 423 586 440
rect 603 423 626 440
rect 643 423 666 440
rect 683 423 706 440
rect 723 423 746 440
rect 763 423 786 440
rect 803 423 826 440
rect 843 423 866 440
rect 883 423 906 440
rect 923 423 946 440
rect 963 423 986 440
rect 1003 423 1026 440
rect 1043 423 1066 440
rect 1083 423 1106 440
rect 1123 423 1146 440
rect 1163 423 1186 440
rect 1203 423 1226 440
rect 1243 423 1266 440
rect 1283 423 1306 440
rect 1323 423 1346 440
rect 1363 423 1386 440
rect 1403 423 1426 440
rect 1443 423 1491 440
rect 83 417 1491 423
rect 83 376 112 417
rect 83 359 89 376
rect 106 359 112 376
rect 83 352 112 359
rect 280 376 309 417
rect 280 359 286 376
rect 303 359 309 376
rect 280 352 309 359
rect 477 376 506 417
rect 477 359 483 376
rect 500 359 506 376
rect 477 352 506 359
rect 674 376 703 417
rect 674 359 680 376
rect 697 359 703 376
rect 674 352 703 359
rect 871 376 900 417
rect 871 359 877 376
rect 894 359 900 376
rect 871 352 900 359
rect 1068 376 1097 417
rect 1068 359 1074 376
rect 1091 359 1097 376
rect 1068 352 1097 359
rect 1265 376 1294 417
rect 1265 359 1271 376
rect 1288 359 1294 376
rect 1265 352 1294 359
rect 1462 376 1491 417
rect 1462 359 1468 376
rect 1485 359 1491 376
rect 1462 352 1491 359
rect 83 28 112 51
rect 83 11 89 28
rect 106 11 112 28
rect 83 -12 112 11
rect 83 -29 89 -12
rect 106 -29 112 -12
rect 83 -52 112 -29
rect 83 -69 89 -52
rect 106 -69 112 -52
rect 83 -92 112 -69
rect 83 -109 89 -92
rect 106 -109 112 -92
rect 83 -116 112 -109
rect 280 28 309 51
rect 280 11 286 28
rect 303 11 309 28
rect 280 -12 309 11
rect 280 -29 286 -12
rect 303 -29 309 -12
rect 280 -52 309 -29
rect 280 -69 286 -52
rect 303 -69 309 -52
rect 280 -92 309 -69
rect 280 -109 286 -92
rect 303 -109 309 -92
rect 280 -116 309 -109
rect 477 28 506 51
rect 477 11 483 28
rect 500 11 506 28
rect 477 -12 506 11
rect 477 -29 483 -12
rect 500 -29 506 -12
rect 477 -52 506 -29
rect 477 -69 483 -52
rect 500 -69 506 -52
rect 477 -92 506 -69
rect 477 -109 483 -92
rect 500 -109 506 -92
rect 477 -116 506 -109
rect 674 28 703 51
rect 674 11 680 28
rect 697 11 703 28
rect 674 -12 703 11
rect 674 -29 680 -12
rect 697 -29 703 -12
rect 674 -52 703 -29
rect 674 -69 680 -52
rect 697 -69 703 -52
rect 674 -92 703 -69
rect 674 -109 680 -92
rect 697 -109 703 -92
rect 674 -116 703 -109
rect 871 28 900 51
rect 871 11 877 28
rect 894 11 900 28
rect 871 -12 900 11
rect 871 -29 877 -12
rect 894 -29 900 -12
rect 871 -52 900 -29
rect 871 -69 877 -52
rect 894 -69 900 -52
rect 871 -92 900 -69
rect 871 -109 877 -92
rect 894 -109 900 -92
rect 871 -116 900 -109
rect 1068 28 1097 51
rect 1068 11 1074 28
rect 1091 11 1097 28
rect 1068 -12 1097 11
rect 1068 -29 1074 -12
rect 1091 -29 1097 -12
rect 1068 -52 1097 -29
rect 1068 -69 1074 -52
rect 1091 -69 1097 -52
rect 1068 -92 1097 -69
rect 1068 -109 1074 -92
rect 1091 -109 1097 -92
rect 1068 -116 1097 -109
rect 1265 28 1294 51
rect 1265 11 1271 28
rect 1288 11 1294 28
rect 1265 -12 1294 11
rect 1265 -29 1271 -12
rect 1288 -29 1294 -12
rect 1265 -52 1294 -29
rect 1265 -69 1271 -52
rect 1288 -69 1294 -52
rect 1265 -92 1294 -69
rect 1265 -109 1271 -92
rect 1288 -109 1294 -92
rect 1265 -116 1294 -109
rect 1462 28 1491 51
rect 1462 11 1468 28
rect 1485 11 1491 28
rect 1462 -12 1491 11
rect 1462 -29 1468 -12
rect 1485 -29 1491 -12
rect 1462 -52 1491 -29
rect 1462 -69 1468 -52
rect 1485 -69 1491 -52
rect 1462 -92 1491 -69
rect 1462 -109 1468 -92
rect 1485 -109 1491 -92
rect 1462 -116 1491 -109
rect 83 -424 112 -417
rect 83 -441 89 -424
rect 106 -441 112 -424
rect 83 -482 112 -441
rect 280 -424 309 -417
rect 280 -441 286 -424
rect 303 -441 309 -424
rect 280 -482 309 -441
rect 477 -424 506 -417
rect 477 -441 483 -424
rect 500 -441 506 -424
rect 477 -482 506 -441
rect 674 -424 703 -417
rect 674 -441 680 -424
rect 697 -441 703 -424
rect 674 -482 703 -441
rect 871 -424 900 -417
rect 871 -441 877 -424
rect 894 -441 900 -424
rect 871 -482 900 -441
rect 1068 -424 1097 -417
rect 1068 -441 1074 -424
rect 1091 -441 1097 -424
rect 1068 -482 1097 -441
rect 1265 -424 1294 -417
rect 1265 -441 1271 -424
rect 1288 -441 1294 -424
rect 1265 -482 1294 -441
rect 1462 -424 1491 -417
rect 1462 -441 1468 -424
rect 1485 -441 1491 -424
rect 1462 -482 1491 -441
rect 83 -488 1491 -482
rect 83 -505 106 -488
rect 123 -505 146 -488
rect 163 -505 186 -488
rect 203 -505 226 -488
rect 243 -505 266 -488
rect 283 -505 306 -488
rect 323 -505 346 -488
rect 363 -505 386 -488
rect 403 -505 426 -488
rect 443 -505 466 -488
rect 483 -505 506 -488
rect 523 -505 546 -488
rect 563 -505 586 -488
rect 603 -505 626 -488
rect 643 -505 666 -488
rect 683 -505 706 -488
rect 723 -505 746 -488
rect 763 -505 786 -488
rect 803 -505 826 -488
rect 843 -505 866 -488
rect 883 -505 906 -488
rect 923 -505 946 -488
rect 963 -505 986 -488
rect 1003 -505 1026 -488
rect 1043 -505 1066 -488
rect 1083 -505 1106 -488
rect 1123 -505 1146 -488
rect 1163 -505 1186 -488
rect 1203 -505 1226 -488
rect 1243 -505 1266 -488
rect 1283 -505 1306 -488
rect 1323 -505 1346 -488
rect 1363 -505 1386 -488
rect 1403 -505 1426 -488
rect 1443 -505 1491 -488
rect 83 -511 1491 -505
<< nsubdiffcont >>
rect 106 423 123 440
rect 146 423 163 440
rect 186 423 203 440
rect 226 423 243 440
rect 266 423 283 440
rect 306 423 323 440
rect 346 423 363 440
rect 386 423 403 440
rect 426 423 443 440
rect 466 423 483 440
rect 506 423 523 440
rect 546 423 563 440
rect 586 423 603 440
rect 626 423 643 440
rect 666 423 683 440
rect 706 423 723 440
rect 746 423 763 440
rect 786 423 803 440
rect 826 423 843 440
rect 866 423 883 440
rect 906 423 923 440
rect 946 423 963 440
rect 986 423 1003 440
rect 1026 423 1043 440
rect 1066 423 1083 440
rect 1106 423 1123 440
rect 1146 423 1163 440
rect 1186 423 1203 440
rect 1226 423 1243 440
rect 1266 423 1283 440
rect 1306 423 1323 440
rect 1346 423 1363 440
rect 1386 423 1403 440
rect 1426 423 1443 440
rect 89 359 106 376
rect 286 359 303 376
rect 483 359 500 376
rect 680 359 697 376
rect 877 359 894 376
rect 1074 359 1091 376
rect 1271 359 1288 376
rect 1468 359 1485 376
rect 89 11 106 28
rect 89 -29 106 -12
rect 89 -69 106 -52
rect 89 -109 106 -92
rect 286 11 303 28
rect 286 -29 303 -12
rect 286 -69 303 -52
rect 286 -109 303 -92
rect 483 11 500 28
rect 483 -29 500 -12
rect 483 -69 500 -52
rect 483 -109 500 -92
rect 680 11 697 28
rect 680 -29 697 -12
rect 680 -69 697 -52
rect 680 -109 697 -92
rect 877 11 894 28
rect 877 -29 894 -12
rect 877 -69 894 -52
rect 877 -109 894 -92
rect 1074 11 1091 28
rect 1074 -29 1091 -12
rect 1074 -69 1091 -52
rect 1074 -109 1091 -92
rect 1271 11 1288 28
rect 1271 -29 1288 -12
rect 1271 -69 1288 -52
rect 1271 -109 1288 -92
rect 1468 11 1485 28
rect 1468 -29 1485 -12
rect 1468 -69 1485 -52
rect 1468 -109 1485 -92
rect 89 -441 106 -424
rect 286 -441 303 -424
rect 483 -441 500 -424
rect 680 -441 697 -424
rect 877 -441 894 -424
rect 1074 -441 1091 -424
rect 1271 -441 1288 -424
rect 1468 -441 1485 -424
rect 106 -505 123 -488
rect 146 -505 163 -488
rect 186 -505 203 -488
rect 226 -505 243 -488
rect 266 -505 283 -488
rect 306 -505 323 -488
rect 346 -505 363 -488
rect 386 -505 403 -488
rect 426 -505 443 -488
rect 466 -505 483 -488
rect 506 -505 523 -488
rect 546 -505 563 -488
rect 586 -505 603 -488
rect 626 -505 643 -488
rect 666 -505 683 -488
rect 706 -505 723 -488
rect 746 -505 763 -488
rect 786 -505 803 -488
rect 826 -505 843 -488
rect 866 -505 883 -488
rect 906 -505 923 -488
rect 946 -505 963 -488
rect 986 -505 1003 -488
rect 1026 -505 1043 -488
rect 1066 -505 1083 -488
rect 1106 -505 1123 -488
rect 1146 -505 1163 -488
rect 1186 -505 1203 -488
rect 1226 -505 1243 -488
rect 1266 -505 1283 -488
rect 1306 -505 1323 -488
rect 1346 -505 1363 -488
rect 1386 -505 1403 -488
rect 1426 -505 1443 -488
<< locali >>
rect 89 376 106 440
rect 123 423 146 440
rect 163 423 186 440
rect 203 423 226 440
rect 243 423 266 440
rect 283 423 306 440
rect 323 423 346 440
rect 363 423 386 440
rect 403 423 426 440
rect 443 423 466 440
rect 483 423 506 440
rect 523 423 546 440
rect 563 423 586 440
rect 603 423 626 440
rect 643 423 666 440
rect 683 423 706 440
rect 723 423 746 440
rect 763 423 786 440
rect 803 423 826 440
rect 843 423 866 440
rect 883 423 906 440
rect 923 423 946 440
rect 963 423 986 440
rect 1003 423 1026 440
rect 1043 423 1066 440
rect 1083 423 1106 440
rect 1123 423 1146 440
rect 1163 423 1186 440
rect 1203 423 1226 440
rect 1243 423 1266 440
rect 1283 423 1306 440
rect 1323 423 1346 440
rect 1363 423 1386 440
rect 1403 423 1426 440
rect 1443 423 1485 440
rect 89 337 106 359
rect 286 376 303 423
rect 286 337 303 359
rect 483 376 500 423
rect 483 337 500 359
rect 680 376 697 423
rect 680 337 697 359
rect 877 376 894 423
rect 877 337 894 359
rect 1074 376 1091 423
rect 1074 337 1091 359
rect 1271 376 1288 423
rect 1271 337 1288 359
rect 1468 376 1485 423
rect 1468 337 1485 359
rect 89 28 106 66
rect 89 -12 106 11
rect 89 -52 106 -29
rect 89 -92 106 -69
rect 89 -131 106 -109
rect 286 28 303 66
rect 286 -12 303 11
rect 286 -52 303 -29
rect 286 -92 303 -69
rect 286 -131 303 -109
rect 483 28 500 66
rect 483 -12 500 11
rect 483 -52 500 -29
rect 483 -92 500 -69
rect 483 -131 500 -109
rect 680 28 697 66
rect 680 -12 697 11
rect 680 -52 697 -29
rect 680 -92 697 -69
rect 680 -131 697 -109
rect 877 28 894 66
rect 877 -12 894 11
rect 877 -52 894 -29
rect 877 -92 894 -69
rect 877 -131 894 -109
rect 1074 28 1091 66
rect 1074 -12 1091 11
rect 1074 -52 1091 -29
rect 1074 -92 1091 -69
rect 1074 -131 1091 -109
rect 1271 28 1288 66
rect 1271 -12 1288 11
rect 1271 -52 1288 -29
rect 1271 -92 1288 -69
rect 1271 -131 1288 -109
rect 1468 28 1485 66
rect 1468 -12 1485 11
rect 1468 -52 1485 -29
rect 1468 -92 1485 -69
rect 1468 -131 1485 -109
rect 89 -424 106 -402
rect 89 -505 106 -441
rect 286 -424 303 -402
rect 286 -488 303 -441
rect 483 -424 500 -402
rect 483 -488 500 -441
rect 680 -424 697 -402
rect 680 -488 697 -441
rect 877 -424 894 -402
rect 877 -488 894 -441
rect 1074 -424 1091 -402
rect 1074 -488 1091 -441
rect 1271 -424 1288 -402
rect 1271 -488 1288 -441
rect 1468 -424 1485 -402
rect 1468 -488 1485 -441
rect 123 -505 146 -488
rect 163 -505 186 -488
rect 203 -505 226 -488
rect 243 -505 266 -488
rect 283 -505 306 -488
rect 323 -505 346 -488
rect 363 -505 386 -488
rect 403 -505 426 -488
rect 443 -505 466 -488
rect 483 -505 506 -488
rect 523 -505 546 -488
rect 563 -505 586 -488
rect 603 -505 626 -488
rect 643 -505 666 -488
rect 683 -505 706 -488
rect 723 -505 746 -488
rect 763 -505 786 -488
rect 803 -505 826 -488
rect 843 -505 866 -488
rect 883 -505 906 -488
rect 923 -505 946 -488
rect 963 -505 986 -488
rect 1003 -505 1026 -488
rect 1043 -505 1066 -488
rect 1083 -505 1106 -488
rect 1123 -505 1146 -488
rect 1163 -505 1186 -488
rect 1203 -505 1226 -488
rect 1243 -505 1266 -488
rect 1283 -505 1306 -488
rect 1323 -505 1346 -488
rect 1363 -505 1386 -488
rect 1403 -505 1426 -488
rect 1443 -505 1485 -488
<< viali >>
rect 106 423 123 440
rect 146 423 163 440
rect 186 423 203 440
rect 226 423 243 440
rect 266 423 283 440
rect 306 423 323 440
rect 346 423 363 440
rect 386 423 403 440
rect 426 423 443 440
rect 466 423 483 440
rect 506 423 523 440
rect 546 423 563 440
rect 586 423 603 440
rect 626 423 643 440
rect 666 423 683 440
rect 706 423 723 440
rect 746 423 763 440
rect 786 423 803 440
rect 826 423 843 440
rect 866 423 883 440
rect 906 423 923 440
rect 946 423 963 440
rect 986 423 1003 440
rect 1026 423 1043 440
rect 1066 423 1083 440
rect 1106 423 1123 440
rect 1146 423 1163 440
rect 1186 423 1203 440
rect 1226 423 1243 440
rect 1266 423 1283 440
rect 1306 423 1323 440
rect 1346 423 1363 440
rect 1386 423 1403 440
rect 1426 423 1443 440
rect 89 359 106 376
rect 286 359 303 376
rect 483 359 500 376
rect 680 359 697 376
rect 877 359 894 376
rect 1074 359 1091 376
rect 1271 359 1288 376
rect 1468 359 1485 376
rect 89 11 106 28
rect 89 -29 106 -12
rect 89 -69 106 -52
rect 89 -109 106 -92
rect 286 11 303 28
rect 286 -29 303 -12
rect 286 -69 303 -52
rect 286 -109 303 -92
rect 483 11 500 28
rect 483 -29 500 -12
rect 483 -69 500 -52
rect 483 -109 500 -92
rect 680 11 697 28
rect 680 -29 697 -12
rect 680 -69 697 -52
rect 680 -109 697 -92
rect 877 11 894 28
rect 877 -29 894 -12
rect 877 -69 894 -52
rect 877 -109 894 -92
rect 1074 11 1091 28
rect 1074 -29 1091 -12
rect 1074 -69 1091 -52
rect 1074 -109 1091 -92
rect 1271 11 1288 28
rect 1271 -29 1288 -12
rect 1271 -69 1288 -52
rect 1271 -109 1288 -92
rect 1468 11 1485 28
rect 1468 -29 1485 -12
rect 1468 -69 1485 -52
rect 1468 -109 1485 -92
rect 89 -441 106 -424
rect 286 -441 303 -424
rect 483 -441 500 -424
rect 680 -441 697 -424
rect 877 -441 894 -424
rect 1074 -441 1091 -424
rect 1271 -441 1288 -424
rect 1468 -441 1485 -424
rect 106 -505 123 -488
rect 146 -505 163 -488
rect 186 -505 203 -488
rect 226 -505 243 -488
rect 266 -505 283 -488
rect 306 -505 323 -488
rect 346 -505 363 -488
rect 386 -505 403 -488
rect 426 -505 443 -488
rect 466 -505 483 -488
rect 506 -505 523 -488
rect 546 -505 563 -488
rect 586 -505 603 -488
rect 626 -505 643 -488
rect 666 -505 683 -488
rect 706 -505 723 -488
rect 746 -505 763 -488
rect 786 -505 803 -488
rect 826 -505 843 -488
rect 866 -505 883 -488
rect 906 -505 923 -488
rect 946 -505 963 -488
rect 986 -505 1003 -488
rect 1026 -505 1043 -488
rect 1066 -505 1083 -488
rect 1106 -505 1123 -488
rect 1146 -505 1163 -488
rect 1186 -505 1203 -488
rect 1226 -505 1243 -488
rect 1266 -505 1283 -488
rect 1306 -505 1323 -488
rect 1346 -505 1363 -488
rect 1386 -505 1403 -488
rect 1426 -505 1443 -488
<< metal1 >>
rect 83 440 1491 446
rect 83 423 106 440
rect 123 423 146 440
rect 163 423 186 440
rect 203 423 226 440
rect 243 423 266 440
rect 283 423 306 440
rect 323 423 346 440
rect 363 423 386 440
rect 403 423 426 440
rect 443 423 466 440
rect 483 423 506 440
rect 523 423 546 440
rect 563 423 586 440
rect 603 423 626 440
rect 643 423 666 440
rect 683 423 706 440
rect 723 423 746 440
rect 763 423 786 440
rect 803 423 826 440
rect 843 423 866 440
rect 883 423 906 440
rect 923 423 946 440
rect 963 423 986 440
rect 1003 423 1026 440
rect 1043 423 1066 440
rect 1083 423 1106 440
rect 1123 423 1146 440
rect 1163 423 1186 440
rect 1203 423 1226 440
rect 1243 423 1266 440
rect 1283 423 1306 440
rect 1323 423 1346 440
rect 1363 423 1386 440
rect 1403 423 1426 440
rect 1443 423 1491 440
rect 83 417 1491 423
rect 83 376 309 417
rect 83 359 89 376
rect 106 370 286 376
rect 106 359 112 370
rect 83 342 112 359
rect 140 342 166 370
rect 183 342 209 370
rect 226 342 252 370
rect 280 359 286 370
rect 303 359 309 376
rect 280 342 309 359
rect 477 376 506 417
rect 477 359 483 376
rect 500 359 506 376
rect 477 342 506 359
rect 674 376 900 417
rect 674 359 680 376
rect 697 370 877 376
rect 697 359 703 370
rect 674 342 703 359
rect 731 342 757 370
rect 774 342 800 370
rect 817 342 843 370
rect 871 359 877 370
rect 894 359 900 376
rect 871 342 900 359
rect 1068 376 1097 417
rect 1068 359 1074 376
rect 1091 359 1097 376
rect 1068 342 1097 359
rect 1265 376 1491 417
rect 1265 359 1271 376
rect 1288 370 1468 376
rect 1288 359 1294 370
rect 1265 342 1294 359
rect 1322 342 1348 370
rect 1365 342 1391 370
rect 1408 342 1434 370
rect 1462 359 1468 370
rect 1485 359 1491 376
rect 1462 342 1491 359
rect 83 33 112 61
rect 140 33 166 61
rect 183 33 209 61
rect 226 33 252 61
rect 280 33 309 61
rect 83 28 309 33
rect 83 11 89 28
rect 106 11 286 28
rect 303 11 309 28
rect 83 0 309 11
rect 83 -12 112 0
rect 83 -29 89 -12
rect 106 -29 112 -12
rect 83 -52 112 -29
rect 83 -69 89 -52
rect 106 -65 112 -52
rect 280 -12 309 0
rect 280 -29 286 -12
rect 303 -29 309 -12
rect 280 -52 309 -29
rect 280 -65 286 -52
rect 106 -69 286 -65
rect 303 -69 309 -52
rect 83 -92 309 -69
rect 83 -109 89 -92
rect 106 -98 286 -92
rect 106 -109 112 -98
rect 83 -126 112 -109
rect 140 -126 166 -98
rect 183 -126 209 -98
rect 226 -126 252 -98
rect 280 -109 286 -98
rect 303 -109 309 -92
rect 280 -126 309 -109
rect 477 28 506 61
rect 477 11 483 28
rect 500 11 506 28
rect 477 -12 506 11
rect 477 -29 483 -12
rect 500 -29 506 -12
rect 477 -52 506 -29
rect 477 -69 483 -52
rect 500 -69 506 -52
rect 477 -92 506 -69
rect 477 -109 483 -92
rect 500 -109 506 -92
rect 477 -126 506 -109
rect 674 33 703 61
rect 731 33 757 61
rect 774 33 800 61
rect 817 33 843 61
rect 871 33 900 61
rect 674 28 900 33
rect 674 11 680 28
rect 697 11 877 28
rect 894 11 900 28
rect 674 0 900 11
rect 674 -12 703 0
rect 674 -29 680 -12
rect 697 -29 703 -12
rect 674 -52 703 -29
rect 674 -69 680 -52
rect 697 -69 703 -52
rect 674 -92 703 -69
rect 674 -109 680 -92
rect 697 -109 703 -92
rect 674 -126 703 -109
rect 871 -12 900 0
rect 871 -29 877 -12
rect 894 -29 900 -12
rect 871 -52 900 -29
rect 871 -69 877 -52
rect 894 -69 900 -52
rect 871 -92 900 -69
rect 871 -109 877 -92
rect 894 -109 900 -92
rect 871 -126 900 -109
rect 1068 28 1097 61
rect 1068 11 1074 28
rect 1091 11 1097 28
rect 1068 -12 1097 11
rect 1068 -29 1074 -12
rect 1091 -29 1097 -12
rect 1068 -52 1097 -29
rect 1068 -69 1074 -52
rect 1091 -69 1097 -52
rect 1068 -92 1097 -69
rect 1068 -109 1074 -92
rect 1091 -109 1097 -92
rect 1068 -126 1097 -109
rect 1265 33 1294 61
rect 1322 33 1348 61
rect 1365 33 1391 61
rect 1408 33 1434 61
rect 1462 33 1491 61
rect 1265 28 1364 33
rect 1265 11 1271 28
rect 1288 11 1364 28
rect 1265 0 1364 11
rect 1365 0 1407 33
rect 1408 28 1491 33
rect 1408 11 1468 28
rect 1485 11 1491 28
rect 1408 0 1491 11
rect 1265 -12 1294 0
rect 1265 -29 1271 -12
rect 1288 -29 1294 -12
rect 1265 -52 1294 -29
rect 1265 -69 1271 -52
rect 1288 -65 1294 -52
rect 1462 -12 1491 0
rect 1462 -29 1468 -12
rect 1485 -29 1491 -12
rect 1462 -52 1491 -29
rect 1462 -65 1468 -52
rect 1288 -69 1468 -65
rect 1485 -69 1491 -52
rect 1265 -92 1491 -69
rect 1265 -109 1271 -92
rect 1288 -98 1468 -92
rect 1288 -109 1294 -98
rect 1265 -126 1294 -109
rect 1322 -126 1348 -98
rect 1365 -126 1391 -98
rect 1408 -126 1434 -98
rect 1462 -109 1468 -98
rect 1485 -109 1491 -92
rect 1462 -126 1491 -109
rect 83 -424 112 -407
rect 83 -441 89 -424
rect 106 -435 112 -424
rect 140 -435 166 -407
rect 183 -435 209 -407
rect 226 -435 252 -407
rect 280 -424 309 -407
rect 280 -435 286 -424
rect 106 -441 286 -435
rect 303 -441 309 -424
rect 83 -482 309 -441
rect 477 -424 506 -407
rect 477 -441 483 -424
rect 500 -441 506 -424
rect 477 -482 506 -441
rect 674 -424 703 -407
rect 674 -441 680 -424
rect 697 -441 703 -424
rect 674 -482 703 -441
rect 871 -424 900 -407
rect 871 -441 877 -424
rect 894 -441 900 -424
rect 871 -482 900 -441
rect 1068 -424 1097 -407
rect 1068 -441 1074 -424
rect 1091 -441 1097 -424
rect 1068 -482 1097 -441
rect 1265 -424 1294 -407
rect 1265 -441 1271 -424
rect 1288 -435 1294 -424
rect 1322 -435 1348 -407
rect 1365 -435 1391 -407
rect 1408 -435 1434 -407
rect 1462 -424 1491 -407
rect 1462 -435 1468 -424
rect 1288 -441 1468 -435
rect 1485 -441 1491 -424
rect 1265 -482 1491 -441
rect 83 -488 1491 -482
rect 83 -505 106 -488
rect 123 -505 146 -488
rect 163 -505 186 -488
rect 203 -505 226 -488
rect 243 -505 266 -488
rect 283 -505 306 -488
rect 323 -505 346 -488
rect 363 -505 386 -488
rect 403 -505 426 -488
rect 443 -505 466 -488
rect 483 -505 506 -488
rect 523 -505 546 -488
rect 563 -505 586 -488
rect 603 -505 626 -488
rect 643 -505 666 -488
rect 683 -505 706 -488
rect 723 -505 746 -488
rect 763 -505 786 -488
rect 803 -505 826 -488
rect 843 -505 866 -488
rect 883 -505 906 -488
rect 923 -505 946 -488
rect 963 -505 986 -488
rect 1003 -505 1026 -488
rect 1043 -505 1066 -488
rect 1083 -505 1106 -488
rect 1123 -505 1146 -488
rect 1163 -505 1186 -488
rect 1203 -505 1226 -488
rect 1243 -505 1266 -488
rect 1283 -505 1306 -488
rect 1323 -505 1346 -488
rect 1363 -505 1386 -488
rect 1403 -505 1426 -488
rect 1443 -505 1491 -488
rect 83 -511 1491 -505
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_0
timestamp 1654596980
transform 1 0 65 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_1
timestamp 1654596980
transform 1 0 262 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_2
timestamp 1654596980
transform 1 0 459 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_3
timestamp 1654596980
transform 1 0 656 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_4
timestamp 1654596980
transform 1 0 853 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_5
timestamp 1654596980
transform 1 0 1050 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_6
timestamp 1654596980
transform 1 0 1247 0 1 0
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_7
timestamp 1654596980
transform 1 0 65 0 1 -468
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_8
timestamp 1654596980
transform 1 0 262 0 1 -468
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_9
timestamp 1654596980
transform 1 0 459 0 1 -468
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_10
timestamp 1654596980
transform 1 0 656 0 1 -468
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_11
timestamp 1654596980
transform 1 0 853 0 1 -468
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_12
timestamp 1654596980
transform 1 0 1050 0 1 -468
box 0 0 262 403
use rf_pfet_01v8_aM02W3p00L0p15  rf_pfet_01v8_aM02W3p00L0p15_13
timestamp 1654596980
transform 1 0 1247 0 1 -468
box 0 0 262 403
<< end >>
