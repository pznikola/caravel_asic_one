magic
tech sky130B
magscale 1 2
timestamp 1654523624
<< psubdiff >>
rect 3858 2454 4882 2520
rect 3858 360 3924 2454
rect 4816 360 4882 2454
rect 3858 294 4882 360
rect 3858 226 3924 294
rect 3858 192 3874 226
rect 3908 192 3924 226
rect 3858 146 3924 192
rect 3858 112 3874 146
rect 3908 112 3924 146
rect 32 42 92 72
rect 32 8 46 42
rect 80 8 92 42
rect 32 -38 92 8
rect 32 -72 46 -38
rect 80 -72 92 -38
rect 32 -118 92 -72
rect 32 -152 46 -118
rect 80 -152 92 -118
rect 32 -198 92 -152
rect 32 -232 46 -198
rect 80 -232 92 -198
rect 32 -278 92 -232
rect 32 -312 46 -278
rect 80 -312 92 -278
rect 32 -358 92 -312
rect 32 -392 46 -358
rect 80 -392 92 -358
rect 32 -482 92 -392
rect 2710 36 2770 72
rect 2710 2 2722 36
rect 2756 2 2770 36
rect 2710 -44 2770 2
rect 2710 -78 2722 -44
rect 2756 -78 2770 -44
rect 2710 -124 2770 -78
rect 2710 -158 2722 -124
rect 2756 -158 2770 -124
rect 2710 -204 2770 -158
rect 2710 -238 2722 -204
rect 2756 -238 2770 -204
rect 2710 -284 2770 -238
rect 2710 -318 2722 -284
rect 2756 -318 2770 -284
rect 2710 -364 2770 -318
rect 2710 -398 2722 -364
rect 2756 -398 2770 -364
rect 2710 -482 2770 -398
rect 3858 66 3924 112
rect 3858 32 3874 66
rect 3908 32 3924 66
rect 3858 -14 3924 32
rect 3858 -48 3874 -14
rect 3908 -48 3924 -14
rect 3858 -94 3924 -48
rect 3858 -128 3874 -94
rect 3908 -128 3924 -94
rect 3858 -174 3924 -128
rect 3858 -208 3874 -174
rect 3908 -208 3924 -174
rect 3858 -254 3924 -208
rect 3858 -288 3874 -254
rect 3908 -288 3924 -254
rect 3858 -334 3924 -288
rect 3858 -368 3874 -334
rect 3908 -368 3924 -334
rect 3858 -414 3924 -368
rect 3858 -448 3874 -414
rect 3908 -448 3924 -414
rect 3858 -494 3924 -448
rect 4816 226 4882 294
rect 4816 192 4832 226
rect 4866 192 4882 226
rect 4816 146 4882 192
rect 4816 112 4832 146
rect 4866 112 4882 146
rect 4816 66 4882 112
rect 4816 32 4832 66
rect 4866 32 4882 66
rect 4816 -14 4882 32
rect 4816 -48 4832 -14
rect 4866 -48 4882 -14
rect 4816 -94 4882 -48
rect 4816 -128 4832 -94
rect 4866 -128 4882 -94
rect 4816 -174 4882 -128
rect 4816 -208 4832 -174
rect 4866 -208 4882 -174
rect 4816 -254 4882 -208
rect 4816 -288 4832 -254
rect 4866 -288 4882 -254
rect 4816 -334 4882 -288
rect 4816 -368 4832 -334
rect 4866 -368 4882 -334
rect 4816 -414 4882 -368
rect 4816 -448 4832 -414
rect 4866 -448 4882 -414
rect 4816 -494 4882 -448
<< psubdiffcont >>
rect 3874 192 3908 226
rect 3874 112 3908 146
rect 46 8 80 42
rect 46 -72 80 -38
rect 46 -152 80 -118
rect 46 -232 80 -198
rect 46 -312 80 -278
rect 46 -392 80 -358
rect 2722 2 2756 36
rect 2722 -78 2756 -44
rect 2722 -158 2756 -124
rect 2722 -238 2756 -204
rect 2722 -318 2756 -284
rect 2722 -398 2756 -364
rect 3874 32 3908 66
rect 3874 -48 3908 -14
rect 3874 -128 3908 -94
rect 3874 -208 3908 -174
rect 3874 -288 3908 -254
rect 3874 -368 3908 -334
rect 3874 -448 3908 -414
rect 4832 192 4866 226
rect 4832 112 4866 146
rect 4832 32 4866 66
rect 4832 -48 4866 -14
rect 4832 -128 4866 -94
rect 4832 -208 4866 -174
rect 4832 -288 4866 -254
rect 4832 -368 4866 -334
rect 4832 -448 4866 -414
<< locali >>
rect 3874 2466 3890 2488
rect 4754 2454 4788 2488
rect 4850 2466 4866 2488
rect 3874 2386 3890 2432
rect 4850 2386 4866 2432
rect 3874 2306 3890 2352
rect 4850 2306 4866 2352
rect 3874 2226 3890 2272
rect 4850 2226 4866 2272
rect 3874 2146 3890 2192
rect 4850 2146 4866 2192
rect 3874 2066 3890 2112
rect 4850 2066 4866 2112
rect 3874 1986 3890 2032
rect 4850 1986 4866 2032
rect 3874 1906 3890 1952
rect 4850 1906 4866 1952
rect 3874 1826 3890 1872
rect 4850 1826 4866 1872
rect 3874 1746 3890 1792
rect 4850 1746 4866 1792
rect 3874 1666 3890 1712
rect 4850 1666 4866 1712
rect 3874 1586 3890 1632
rect 4850 1586 4866 1632
rect 3874 1506 3890 1552
rect 4850 1506 4866 1552
rect 3874 1426 3890 1472
rect 4850 1426 4866 1472
rect 3874 1346 3890 1392
rect 4850 1346 4866 1392
rect 3874 1266 3890 1312
rect 4850 1266 4866 1312
rect 3874 1186 3890 1232
rect 4850 1186 4866 1232
rect 3874 1106 3890 1152
rect 4850 1106 4866 1152
rect 3874 1026 3890 1072
rect 4850 1026 4866 1072
rect 3874 946 3890 992
rect 4850 946 4866 992
rect 3874 866 3890 912
rect 4850 866 4866 912
rect 3874 786 3890 832
rect 4850 786 4866 832
rect 3874 706 3890 752
rect 4850 706 4866 752
rect 3874 626 3890 672
rect 4850 626 4866 672
rect 3874 546 3890 592
rect 4850 546 4866 592
rect 3874 466 3890 512
rect 4850 466 4866 512
rect 3874 386 3890 432
rect 4850 386 4866 432
rect 3874 310 3890 352
rect 4850 310 4866 352
rect 3874 306 3924 310
rect 3908 272 3924 306
rect 3874 266 3924 272
rect 4816 306 4866 310
rect 4816 272 4832 306
rect 4816 266 4866 272
rect 3874 226 3908 266
rect 3874 146 3908 192
rect 46 42 80 84
rect 46 -38 80 8
rect 46 -118 80 -72
rect 46 -198 80 -152
rect 46 -278 80 -232
rect 46 -358 80 -312
rect 46 -494 80 -392
rect 2722 36 2756 84
rect 2722 -44 2756 2
rect 2722 -124 2756 -78
rect 2722 -204 2756 -158
rect 2722 -284 2756 -238
rect 2722 -364 2756 -318
rect 2722 -494 2756 -398
rect 3874 66 3908 112
rect 3874 -14 3908 32
rect 3874 -94 3908 -48
rect 3874 -174 3908 -128
rect 3874 -254 3908 -208
rect 3874 -334 3908 -288
rect 3874 -414 3908 -368
rect 3874 -494 3908 -448
rect 4832 226 4866 266
rect 4832 146 4866 192
rect 4832 66 4866 112
rect 4832 -14 4866 32
rect 4832 -94 4866 -48
rect 4832 -174 4866 -128
rect 4832 -254 4866 -208
rect 4832 -334 4866 -288
rect 4832 -414 4866 -368
rect 4832 -494 4866 -448
<< viali >>
rect 3874 2432 3908 2466
rect 4832 2432 4866 2466
rect 3874 2352 3908 2386
rect 4832 2352 4866 2386
rect 3874 2272 3908 2306
rect 4832 2272 4866 2306
rect 3874 2192 3908 2226
rect 4832 2192 4866 2226
rect 3874 2112 3908 2146
rect 4832 2112 4866 2146
rect 3874 2032 3908 2066
rect 4832 2032 4866 2066
rect 3874 1952 3908 1986
rect 4832 1952 4866 1986
rect 3874 1872 3908 1906
rect 4832 1872 4866 1906
rect 3874 1792 3908 1826
rect 4832 1792 4866 1826
rect 3874 1712 3908 1746
rect 4832 1712 4866 1746
rect 3874 1632 3908 1666
rect 4832 1632 4866 1666
rect 3874 1552 3908 1586
rect 4832 1552 4866 1586
rect 3874 1472 3908 1506
rect 4832 1472 4866 1506
rect 3874 1392 3908 1426
rect 4832 1392 4866 1426
rect 3874 1312 3908 1346
rect 4832 1312 4866 1346
rect 3874 1232 3908 1266
rect 4832 1232 4866 1266
rect 3874 1152 3908 1186
rect 4832 1152 4866 1186
rect 3874 1072 3908 1106
rect 4832 1072 4866 1106
rect 3874 992 3908 1026
rect 4832 992 4866 1026
rect 3874 912 3908 946
rect 4832 912 4866 946
rect 3874 832 3908 866
rect 4832 832 4866 866
rect 3874 752 3908 786
rect 4832 752 4866 786
rect 3874 672 3908 706
rect 4832 672 4866 706
rect 3874 592 3908 626
rect 4832 592 4866 626
rect 3874 512 3908 546
rect 4832 512 4866 546
rect 3874 432 3908 466
rect 4832 432 4866 466
rect 3874 352 3908 386
rect 4832 352 4866 386
rect 3874 272 3908 306
rect 4832 272 4866 306
rect 3874 192 3908 226
rect 3874 112 3908 146
rect 46 8 80 42
rect 46 -72 80 -38
rect 46 -152 80 -118
rect 46 -232 80 -198
rect 46 -312 80 -278
rect 46 -392 80 -358
rect 2722 2 2756 36
rect 2722 -78 2756 -44
rect 2722 -158 2756 -124
rect 2722 -238 2756 -204
rect 2722 -318 2756 -284
rect 2722 -398 2756 -364
rect 3874 32 3908 66
rect 3874 -48 3908 -14
rect 3874 -128 3908 -94
rect 3874 -208 3908 -174
rect 3874 -288 3908 -254
rect 3874 -368 3908 -334
rect 3874 -448 3908 -414
rect 4832 192 4866 226
rect 4832 112 4866 146
rect 4832 32 4866 66
rect 4832 -48 4866 -14
rect 4832 -128 4866 -94
rect 4832 -208 4866 -174
rect 4832 -288 4866 -254
rect 4832 -368 4866 -334
rect 4832 -448 4866 -414
<< metal1 >>
rect 3858 2466 3924 2520
rect 3858 2432 3874 2466
rect 3908 2432 3924 2466
rect 3858 2386 3924 2432
rect 3858 2352 3874 2386
rect 3908 2352 3924 2386
rect 3858 2306 3924 2352
rect 3858 2272 3874 2306
rect 3908 2272 3924 2306
rect 4020 2510 4720 2534
rect 4020 2458 4044 2510
rect 4096 2458 4144 2510
rect 4196 2458 4244 2510
rect 4296 2458 4344 2510
rect 4396 2458 4444 2510
rect 4496 2458 4544 2510
rect 4596 2458 4644 2510
rect 4696 2458 4720 2510
rect 4020 2410 4720 2458
rect 4020 2358 4044 2410
rect 4096 2358 4144 2410
rect 4196 2358 4244 2410
rect 4296 2358 4344 2410
rect 4396 2358 4444 2410
rect 4496 2358 4544 2410
rect 4596 2358 4644 2410
rect 4696 2358 4720 2410
rect 4020 2286 4720 2358
rect 4816 2466 4882 2520
rect 4816 2432 4832 2466
rect 4866 2432 4882 2466
rect 4816 2386 4882 2432
rect 4816 2352 4832 2386
rect 4866 2352 4882 2386
rect 4816 2306 4882 2352
rect 3858 2226 3924 2272
rect 3858 2192 3874 2226
rect 3908 2192 3924 2226
rect 3858 2146 3924 2192
rect 3858 2112 3874 2146
rect 3908 2112 3924 2146
rect 3858 2066 3924 2112
rect 3858 2032 3874 2066
rect 3908 2032 3924 2066
rect 3858 1986 3924 2032
rect 3858 1952 3874 1986
rect 3908 1952 3924 1986
rect 3858 1906 3924 1952
rect 3858 1872 3874 1906
rect 3908 1872 3924 1906
rect 3858 1826 3924 1872
rect 3858 1792 3874 1826
rect 3908 1792 3924 1826
rect 3858 1746 3924 1792
rect 3858 1712 3874 1746
rect 3908 1712 3924 1746
rect 3858 1666 3924 1712
rect 3858 1632 3874 1666
rect 3908 1632 3924 1666
rect 3858 1586 3924 1632
rect 3858 1552 3874 1586
rect 3908 1552 3924 1586
rect 4816 2272 4832 2306
rect 4866 2272 4882 2306
rect 4816 2226 4882 2272
rect 4816 2192 4832 2226
rect 4866 2192 4882 2226
rect 4816 2146 4882 2192
rect 4816 2112 4832 2146
rect 4866 2112 4882 2146
rect 4816 2066 4882 2112
rect 4816 2032 4832 2066
rect 4866 2032 4882 2066
rect 4816 1986 4882 2032
rect 4816 1952 4832 1986
rect 4866 1952 4882 1986
rect 4816 1906 4882 1952
rect 4816 1872 4832 1906
rect 4866 1872 4882 1906
rect 4816 1826 4882 1872
rect 4816 1792 4832 1826
rect 4866 1792 4882 1826
rect 4816 1746 4882 1792
rect 4816 1712 4832 1746
rect 4866 1712 4882 1746
rect 4816 1666 4882 1712
rect 4816 1632 4832 1666
rect 4866 1632 4882 1666
rect 4816 1586 4882 1632
rect 3858 1506 3924 1552
rect 3858 1472 3874 1506
rect 3908 1472 3924 1506
rect 3858 1426 3924 1472
rect 3858 1392 3874 1426
rect 3908 1392 3924 1426
rect 3858 1346 3924 1392
rect 3858 1312 3874 1346
rect 3908 1312 3924 1346
rect 3858 1266 3924 1312
rect 3858 1232 3874 1266
rect 3908 1232 3924 1266
rect 3858 1186 3924 1232
rect 4020 1514 4720 1584
rect 4020 1462 4040 1514
rect 4092 1462 4140 1514
rect 4192 1462 4240 1514
rect 4292 1462 4340 1514
rect 4392 1462 4440 1514
rect 4492 1462 4540 1514
rect 4592 1462 4640 1514
rect 4692 1462 4720 1514
rect 4020 1414 4720 1462
rect 4020 1362 4040 1414
rect 4092 1362 4140 1414
rect 4192 1362 4240 1414
rect 4292 1362 4340 1414
rect 4392 1362 4440 1414
rect 4492 1362 4540 1414
rect 4592 1362 4640 1414
rect 4692 1362 4720 1414
rect 4020 1314 4720 1362
rect 4020 1262 4040 1314
rect 4092 1262 4140 1314
rect 4192 1262 4240 1314
rect 4292 1262 4340 1314
rect 4392 1262 4440 1314
rect 4492 1262 4540 1314
rect 4592 1262 4640 1314
rect 4692 1262 4720 1314
rect 4020 1214 4720 1262
rect 4816 1552 4832 1586
rect 4866 1552 4882 1586
rect 4816 1506 4882 1552
rect 4816 1472 4832 1506
rect 4866 1472 4882 1506
rect 4816 1426 4882 1472
rect 4816 1392 4832 1426
rect 4866 1392 4882 1426
rect 4816 1346 4882 1392
rect 4816 1312 4832 1346
rect 4866 1312 4882 1346
rect 4816 1266 4882 1312
rect 4816 1232 4832 1266
rect 4866 1232 4882 1266
rect 3858 1152 3874 1186
rect 3908 1152 3924 1186
rect 3858 1106 3924 1152
rect 3858 1072 3874 1106
rect 3908 1072 3924 1106
rect 3858 1026 3924 1072
rect 3858 992 3874 1026
rect 3908 992 3924 1026
rect 3858 946 3924 992
rect 3858 912 3874 946
rect 3908 912 3924 946
rect 3858 866 3924 912
rect 3858 832 3874 866
rect 3908 832 3924 866
rect 3858 786 3924 832
rect 3858 752 3874 786
rect 3908 752 3924 786
rect 3858 706 3924 752
rect 3858 672 3874 706
rect 3908 672 3924 706
rect 3858 626 3924 672
rect 3858 592 3874 626
rect 3908 592 3924 626
rect 3858 546 3924 592
rect 3858 512 3874 546
rect 3908 512 3924 546
rect 4816 1186 4882 1232
rect 4816 1152 4832 1186
rect 4866 1152 4882 1186
rect 4816 1106 4882 1152
rect 4816 1072 4832 1106
rect 4866 1072 4882 1106
rect 4816 1026 4882 1072
rect 4816 992 4832 1026
rect 4866 992 4882 1026
rect 4816 946 4882 992
rect 4816 912 4832 946
rect 4866 912 4882 946
rect 4816 866 4882 912
rect 4816 832 4832 866
rect 4866 832 4882 866
rect 4816 786 4882 832
rect 4816 752 4832 786
rect 4866 752 4882 786
rect 4816 706 4882 752
rect 4816 672 4832 706
rect 4866 672 4882 706
rect 4816 626 4882 672
rect 4816 592 4832 626
rect 4866 592 4882 626
rect 4816 546 4882 592
rect 4816 512 4832 546
rect 4866 512 4882 546
rect 3858 466 3924 512
rect 3858 432 3874 466
rect 3908 432 3924 466
rect 3858 386 3924 432
rect 3858 352 3874 386
rect 3908 352 3924 386
rect 3858 306 3924 352
rect 3858 272 3874 306
rect 3908 272 3924 306
rect 3858 226 3924 272
rect 4020 442 4720 512
rect 4020 390 4044 442
rect 4096 390 4144 442
rect 4196 390 4244 442
rect 4296 390 4344 442
rect 4396 390 4444 442
rect 4496 390 4544 442
rect 4596 390 4644 442
rect 4696 390 4720 442
rect 4020 342 4720 390
rect 4020 290 4044 342
rect 4096 290 4144 342
rect 4196 290 4244 342
rect 4296 290 4344 342
rect 4396 290 4444 342
rect 4496 290 4544 342
rect 4596 290 4644 342
rect 4696 290 4720 342
rect 4020 266 4720 290
rect 4816 466 4882 512
rect 4816 432 4832 466
rect 4866 432 4882 466
rect 4816 386 4882 432
rect 4816 352 4832 386
rect 4866 352 4882 386
rect 4816 306 4882 352
rect 4816 272 4832 306
rect 4866 272 4882 306
rect 3858 192 3874 226
rect 3908 192 3924 226
rect 3858 146 3924 192
rect 3858 112 3874 146
rect 3908 112 3924 146
rect 32 42 92 72
rect 32 8 46 42
rect 80 8 92 42
rect 32 -38 92 8
rect 32 -72 46 -38
rect 80 -72 92 -38
rect 32 -118 92 -72
rect 32 -152 46 -118
rect 80 -152 92 -118
rect 32 -198 92 -152
rect 32 -232 46 -198
rect 80 -232 92 -198
rect 32 -278 92 -232
rect 32 -312 46 -278
rect 80 -312 92 -278
rect 32 -358 92 -312
rect 32 -392 46 -358
rect 80 -392 92 -358
rect 32 -482 92 -392
rect 2710 36 2770 72
rect 2710 2 2722 36
rect 2756 2 2770 36
rect 2710 -44 2770 2
rect 2710 -78 2722 -44
rect 2756 -78 2770 -44
rect 2710 -124 2770 -78
rect 2710 -158 2722 -124
rect 2756 -158 2770 -124
rect 2710 -204 2770 -158
rect 2710 -238 2722 -204
rect 2756 -238 2770 -204
rect 2710 -284 2770 -238
rect 2710 -318 2722 -284
rect 2756 -318 2770 -284
rect 2710 -364 2770 -318
rect 2710 -398 2722 -364
rect 2756 -398 2770 -364
rect 2710 -482 2770 -398
rect 3858 66 3924 112
rect 3858 32 3874 66
rect 3908 32 3924 66
rect 3858 -14 3924 32
rect 3858 -48 3874 -14
rect 3908 -48 3924 -14
rect 3858 -94 3924 -48
rect 3858 -128 3874 -94
rect 3908 -128 3924 -94
rect 3858 -174 3924 -128
rect 3858 -208 3874 -174
rect 3908 -208 3924 -174
rect 3858 -254 3924 -208
rect 3858 -288 3874 -254
rect 3908 -288 3924 -254
rect 3858 -334 3924 -288
rect 3858 -368 3874 -334
rect 3908 -368 3924 -334
rect 3858 -414 3924 -368
rect 3858 -448 3874 -414
rect 3908 -448 3924 -414
rect 3858 -482 3924 -448
rect 4816 226 4882 272
rect 4816 192 4832 226
rect 4866 192 4882 226
rect 4816 146 4882 192
rect 4816 112 4832 146
rect 4866 112 4882 146
rect 4816 66 4882 112
rect 4816 32 4832 66
rect 4866 32 4882 66
rect 4816 -14 4882 32
rect 4816 -48 4832 -14
rect 4866 -48 4882 -14
rect 4816 -94 4882 -48
rect 4816 -128 4832 -94
rect 4866 -128 4882 -94
rect 4816 -174 4882 -128
rect 4816 -208 4832 -174
rect 4866 -208 4882 -174
rect 4816 -254 4882 -208
rect 4816 -288 4832 -254
rect 4866 -288 4882 -254
rect 4816 -334 4882 -288
rect 4816 -368 4832 -334
rect 4866 -368 4882 -334
rect 4816 -414 4882 -368
rect 4816 -448 4832 -414
rect 4866 -448 4882 -414
rect 4816 -482 4882 -448
<< via1 >>
rect 4044 2458 4096 2510
rect 4144 2458 4196 2510
rect 4244 2458 4296 2510
rect 4344 2458 4396 2510
rect 4444 2458 4496 2510
rect 4544 2458 4596 2510
rect 4644 2458 4696 2510
rect 4044 2358 4096 2410
rect 4144 2358 4196 2410
rect 4244 2358 4296 2410
rect 4344 2358 4396 2410
rect 4444 2358 4496 2410
rect 4544 2358 4596 2410
rect 4644 2358 4696 2410
rect 4040 1462 4092 1514
rect 4140 1462 4192 1514
rect 4240 1462 4292 1514
rect 4340 1462 4392 1514
rect 4440 1462 4492 1514
rect 4540 1462 4592 1514
rect 4640 1462 4692 1514
rect 4040 1362 4092 1414
rect 4140 1362 4192 1414
rect 4240 1362 4292 1414
rect 4340 1362 4392 1414
rect 4440 1362 4492 1414
rect 4540 1362 4592 1414
rect 4640 1362 4692 1414
rect 4040 1262 4092 1314
rect 4140 1262 4192 1314
rect 4240 1262 4292 1314
rect 4340 1262 4392 1314
rect 4440 1262 4492 1314
rect 4540 1262 4592 1314
rect 4640 1262 4692 1314
rect 4044 390 4096 442
rect 4144 390 4196 442
rect 4244 390 4296 442
rect 4344 390 4396 442
rect 4444 390 4496 442
rect 4544 390 4596 442
rect 4644 390 4696 442
rect 4044 290 4096 342
rect 4144 290 4196 342
rect 4244 290 4296 342
rect 4344 290 4396 342
rect 4444 290 4496 342
rect 4544 290 4596 342
rect 4644 290 4696 342
<< metal2 >>
rect 4020 2514 4720 2534
rect 4020 2454 4040 2514
rect 4100 2454 4140 2514
rect 4200 2454 4240 2514
rect 4300 2454 4340 2514
rect 4400 2454 4440 2514
rect 4500 2454 4540 2514
rect 4600 2454 4640 2514
rect 4700 2454 4720 2514
rect 4020 2414 4720 2454
rect 4020 2354 4040 2414
rect 4100 2354 4140 2414
rect 4200 2354 4240 2414
rect 4300 2354 4340 2414
rect 4400 2354 4440 2414
rect 4500 2354 4540 2414
rect 4600 2354 4640 2414
rect 4700 2354 4720 2414
rect 4020 2334 4720 2354
rect 4020 1518 4720 1584
rect 4020 1458 4036 1518
rect 4096 1458 4136 1518
rect 4196 1458 4236 1518
rect 4296 1458 4336 1518
rect 4396 1458 4436 1518
rect 4496 1458 4536 1518
rect 4596 1458 4636 1518
rect 4696 1458 4720 1518
rect 4020 1418 4720 1458
rect 4020 1358 4036 1418
rect 4096 1358 4136 1418
rect 4196 1358 4236 1418
rect 4296 1358 4336 1418
rect 4396 1358 4436 1418
rect 4496 1358 4536 1418
rect 4596 1358 4636 1418
rect 4696 1358 4720 1418
rect 4020 1318 4720 1358
rect 4020 1258 4036 1318
rect 4096 1258 4136 1318
rect 4196 1258 4236 1318
rect 4296 1258 4336 1318
rect 4396 1258 4436 1318
rect 4496 1258 4536 1318
rect 4596 1258 4636 1318
rect 4696 1258 4720 1318
rect 4020 1214 4720 1258
rect 4020 446 4720 466
rect 4020 386 4040 446
rect 4100 386 4140 446
rect 4200 386 4240 446
rect 4300 386 4340 446
rect 4400 386 4440 446
rect 4500 386 4540 446
rect 4600 386 4640 446
rect 4700 386 4720 446
rect 4020 346 4720 386
rect 4020 286 4040 346
rect 4100 286 4140 346
rect 4200 286 4240 346
rect 4300 286 4340 346
rect 4400 286 4440 346
rect 4500 286 4540 346
rect 4600 286 4640 346
rect 4700 286 4720 346
rect 4020 266 4720 286
<< via2 >>
rect 4040 2510 4100 2514
rect 4040 2458 4044 2510
rect 4044 2458 4096 2510
rect 4096 2458 4100 2510
rect 4040 2454 4100 2458
rect 4140 2510 4200 2514
rect 4140 2458 4144 2510
rect 4144 2458 4196 2510
rect 4196 2458 4200 2510
rect 4140 2454 4200 2458
rect 4240 2510 4300 2514
rect 4240 2458 4244 2510
rect 4244 2458 4296 2510
rect 4296 2458 4300 2510
rect 4240 2454 4300 2458
rect 4340 2510 4400 2514
rect 4340 2458 4344 2510
rect 4344 2458 4396 2510
rect 4396 2458 4400 2510
rect 4340 2454 4400 2458
rect 4440 2510 4500 2514
rect 4440 2458 4444 2510
rect 4444 2458 4496 2510
rect 4496 2458 4500 2510
rect 4440 2454 4500 2458
rect 4540 2510 4600 2514
rect 4540 2458 4544 2510
rect 4544 2458 4596 2510
rect 4596 2458 4600 2510
rect 4540 2454 4600 2458
rect 4640 2510 4700 2514
rect 4640 2458 4644 2510
rect 4644 2458 4696 2510
rect 4696 2458 4700 2510
rect 4640 2454 4700 2458
rect 4040 2410 4100 2414
rect 4040 2358 4044 2410
rect 4044 2358 4096 2410
rect 4096 2358 4100 2410
rect 4040 2354 4100 2358
rect 4140 2410 4200 2414
rect 4140 2358 4144 2410
rect 4144 2358 4196 2410
rect 4196 2358 4200 2410
rect 4140 2354 4200 2358
rect 4240 2410 4300 2414
rect 4240 2358 4244 2410
rect 4244 2358 4296 2410
rect 4296 2358 4300 2410
rect 4240 2354 4300 2358
rect 4340 2410 4400 2414
rect 4340 2358 4344 2410
rect 4344 2358 4396 2410
rect 4396 2358 4400 2410
rect 4340 2354 4400 2358
rect 4440 2410 4500 2414
rect 4440 2358 4444 2410
rect 4444 2358 4496 2410
rect 4496 2358 4500 2410
rect 4440 2354 4500 2358
rect 4540 2410 4600 2414
rect 4540 2358 4544 2410
rect 4544 2358 4596 2410
rect 4596 2358 4600 2410
rect 4540 2354 4600 2358
rect 4640 2410 4700 2414
rect 4640 2358 4644 2410
rect 4644 2358 4696 2410
rect 4696 2358 4700 2410
rect 4640 2354 4700 2358
rect 4036 1514 4096 1518
rect 4036 1462 4040 1514
rect 4040 1462 4092 1514
rect 4092 1462 4096 1514
rect 4036 1458 4096 1462
rect 4136 1514 4196 1518
rect 4136 1462 4140 1514
rect 4140 1462 4192 1514
rect 4192 1462 4196 1514
rect 4136 1458 4196 1462
rect 4236 1514 4296 1518
rect 4236 1462 4240 1514
rect 4240 1462 4292 1514
rect 4292 1462 4296 1514
rect 4236 1458 4296 1462
rect 4336 1514 4396 1518
rect 4336 1462 4340 1514
rect 4340 1462 4392 1514
rect 4392 1462 4396 1514
rect 4336 1458 4396 1462
rect 4436 1514 4496 1518
rect 4436 1462 4440 1514
rect 4440 1462 4492 1514
rect 4492 1462 4496 1514
rect 4436 1458 4496 1462
rect 4536 1514 4596 1518
rect 4536 1462 4540 1514
rect 4540 1462 4592 1514
rect 4592 1462 4596 1514
rect 4536 1458 4596 1462
rect 4636 1514 4696 1518
rect 4636 1462 4640 1514
rect 4640 1462 4692 1514
rect 4692 1462 4696 1514
rect 4636 1458 4696 1462
rect 4036 1414 4096 1418
rect 4036 1362 4040 1414
rect 4040 1362 4092 1414
rect 4092 1362 4096 1414
rect 4036 1358 4096 1362
rect 4136 1414 4196 1418
rect 4136 1362 4140 1414
rect 4140 1362 4192 1414
rect 4192 1362 4196 1414
rect 4136 1358 4196 1362
rect 4236 1414 4296 1418
rect 4236 1362 4240 1414
rect 4240 1362 4292 1414
rect 4292 1362 4296 1414
rect 4236 1358 4296 1362
rect 4336 1414 4396 1418
rect 4336 1362 4340 1414
rect 4340 1362 4392 1414
rect 4392 1362 4396 1414
rect 4336 1358 4396 1362
rect 4436 1414 4496 1418
rect 4436 1362 4440 1414
rect 4440 1362 4492 1414
rect 4492 1362 4496 1414
rect 4436 1358 4496 1362
rect 4536 1414 4596 1418
rect 4536 1362 4540 1414
rect 4540 1362 4592 1414
rect 4592 1362 4596 1414
rect 4536 1358 4596 1362
rect 4636 1414 4696 1418
rect 4636 1362 4640 1414
rect 4640 1362 4692 1414
rect 4692 1362 4696 1414
rect 4636 1358 4696 1362
rect 4036 1314 4096 1318
rect 4036 1262 4040 1314
rect 4040 1262 4092 1314
rect 4092 1262 4096 1314
rect 4036 1258 4096 1262
rect 4136 1314 4196 1318
rect 4136 1262 4140 1314
rect 4140 1262 4192 1314
rect 4192 1262 4196 1314
rect 4136 1258 4196 1262
rect 4236 1314 4296 1318
rect 4236 1262 4240 1314
rect 4240 1262 4292 1314
rect 4292 1262 4296 1314
rect 4236 1258 4296 1262
rect 4336 1314 4396 1318
rect 4336 1262 4340 1314
rect 4340 1262 4392 1314
rect 4392 1262 4396 1314
rect 4336 1258 4396 1262
rect 4436 1314 4496 1318
rect 4436 1262 4440 1314
rect 4440 1262 4492 1314
rect 4492 1262 4496 1314
rect 4436 1258 4496 1262
rect 4536 1314 4596 1318
rect 4536 1262 4540 1314
rect 4540 1262 4592 1314
rect 4592 1262 4596 1314
rect 4536 1258 4596 1262
rect 4636 1314 4696 1318
rect 4636 1262 4640 1314
rect 4640 1262 4692 1314
rect 4692 1262 4696 1314
rect 4636 1258 4696 1262
rect 4040 442 4100 446
rect 4040 390 4044 442
rect 4044 390 4096 442
rect 4096 390 4100 442
rect 4040 386 4100 390
rect 4140 442 4200 446
rect 4140 390 4144 442
rect 4144 390 4196 442
rect 4196 390 4200 442
rect 4140 386 4200 390
rect 4240 442 4300 446
rect 4240 390 4244 442
rect 4244 390 4296 442
rect 4296 390 4300 442
rect 4240 386 4300 390
rect 4340 442 4400 446
rect 4340 390 4344 442
rect 4344 390 4396 442
rect 4396 390 4400 442
rect 4340 386 4400 390
rect 4440 442 4500 446
rect 4440 390 4444 442
rect 4444 390 4496 442
rect 4496 390 4500 442
rect 4440 386 4500 390
rect 4540 442 4600 446
rect 4540 390 4544 442
rect 4544 390 4596 442
rect 4596 390 4600 442
rect 4540 386 4600 390
rect 4640 442 4700 446
rect 4640 390 4644 442
rect 4644 390 4696 442
rect 4696 390 4700 442
rect 4640 386 4700 390
rect 4040 342 4100 346
rect 4040 290 4044 342
rect 4044 290 4096 342
rect 4096 290 4100 342
rect 4040 286 4100 290
rect 4140 342 4200 346
rect 4140 290 4144 342
rect 4144 290 4196 342
rect 4196 290 4200 342
rect 4140 286 4200 290
rect 4240 342 4300 346
rect 4240 290 4244 342
rect 4244 290 4296 342
rect 4296 290 4300 342
rect 4240 286 4300 290
rect 4340 342 4400 346
rect 4340 290 4344 342
rect 4344 290 4396 342
rect 4396 290 4400 342
rect 4340 286 4400 290
rect 4440 342 4500 346
rect 4440 290 4444 342
rect 4444 290 4496 342
rect 4496 290 4500 342
rect 4440 286 4500 290
rect 4540 342 4600 346
rect 4540 290 4544 342
rect 4544 290 4596 342
rect 4596 290 4600 342
rect 4540 286 4600 290
rect 4640 342 4700 346
rect 4640 290 4644 342
rect 4644 290 4696 342
rect 4696 290 4700 342
rect 4640 286 4700 290
<< metal3 >>
rect 1357 2514 4908 2534
rect 1357 2454 4040 2514
rect 4100 2454 4140 2514
rect 4200 2454 4240 2514
rect 4300 2454 4340 2514
rect 4400 2454 4440 2514
rect 4500 2454 4540 2514
rect 4600 2454 4640 2514
rect 4700 2454 4908 2514
rect 1357 2414 4908 2454
rect 1357 2354 4040 2414
rect 4100 2354 4140 2414
rect 4200 2354 4240 2414
rect 4300 2354 4340 2414
rect 4400 2354 4440 2414
rect 4500 2354 4540 2414
rect 4600 2354 4640 2414
rect 4700 2354 4908 2414
rect 1357 2334 4908 2354
rect 3848 1550 4720 1584
rect 3848 1486 3876 1550
rect 3940 1486 3956 1550
rect 4020 1518 4720 1550
rect 4020 1486 4036 1518
rect 3848 1466 4036 1486
rect 3848 1402 3876 1466
rect 3940 1402 3956 1466
rect 4020 1458 4036 1466
rect 4096 1458 4136 1518
rect 4196 1458 4236 1518
rect 4296 1458 4336 1518
rect 4396 1458 4436 1518
rect 4496 1458 4536 1518
rect 4596 1458 4636 1518
rect 4696 1458 4720 1518
rect 4020 1418 4720 1458
rect 4020 1402 4036 1418
rect 3848 1382 4036 1402
rect 3848 1318 3876 1382
rect 3940 1318 3956 1382
rect 4020 1358 4036 1382
rect 4096 1358 4136 1418
rect 4196 1358 4236 1418
rect 4296 1358 4336 1418
rect 4396 1358 4436 1418
rect 4496 1358 4536 1418
rect 4596 1358 4636 1418
rect 4696 1358 4720 1418
rect 4020 1318 4720 1358
rect 3848 1302 4036 1318
rect 3848 1238 3876 1302
rect 3940 1238 3956 1302
rect 4020 1258 4036 1302
rect 4096 1258 4136 1318
rect 4196 1258 4236 1318
rect 4296 1258 4336 1318
rect 4396 1258 4436 1318
rect 4496 1258 4536 1318
rect 4596 1258 4636 1318
rect 4696 1258 4720 1318
rect 4020 1238 4720 1258
rect 3848 1214 4720 1238
rect 2994 538 3880 738
rect 3680 466 3880 538
rect 3680 446 4908 466
rect 3680 386 4040 446
rect 4100 386 4140 446
rect 4200 386 4240 446
rect 4300 386 4340 446
rect 4400 386 4440 446
rect 4500 386 4540 446
rect 4600 386 4640 446
rect 4700 386 4908 446
rect 3680 346 4908 386
rect 3680 286 4040 346
rect 4100 286 4140 346
rect 4200 286 4240 346
rect 4300 286 4340 346
rect 4400 286 4440 346
rect 4500 286 4540 346
rect 4600 286 4640 346
rect 4700 286 4908 346
rect 3680 266 4908 286
<< via3 >>
rect 3876 1486 3940 1550
rect 3956 1486 4020 1550
rect 3876 1402 3940 1466
rect 3956 1402 4020 1466
rect 3876 1318 3940 1382
rect 3956 1318 4020 1382
rect 3876 1238 3940 1302
rect 3956 1238 4020 1302
<< metal4 >>
rect 3770 3446 4130 3512
rect 3770 3210 3830 3446
rect 4066 3210 4130 3446
rect 3770 3126 4130 3210
rect 3770 2890 3828 3126
rect 4064 2890 4130 3126
rect 3770 2840 4130 2890
rect 3848 1550 4048 2840
rect 3848 1486 3876 1550
rect 3940 1486 3956 1550
rect 4020 1486 4048 1550
rect 3848 1466 4048 1486
rect 3848 1402 3876 1466
rect 3940 1402 3956 1466
rect 4020 1402 4048 1466
rect 3848 1382 4048 1402
rect 3848 1318 3876 1382
rect 3940 1318 3956 1382
rect 4020 1318 4048 1382
rect 3848 1302 4048 1318
rect 3848 1238 3876 1302
rect 3940 1238 3956 1302
rect 4020 1238 4048 1302
rect 3848 1214 4048 1238
rect 3316 -60 3650 904
rect 3316 -296 3368 -60
rect 3604 -296 3650 -60
rect 3316 -348 3650 -296
<< via4 >>
rect 3830 3210 4066 3446
rect 3828 2890 4064 3126
rect 3368 -296 3604 -60
<< metal5 >>
rect 32 3446 4908 3512
rect 32 3210 3830 3446
rect 4066 3210 4908 3446
rect 32 3126 4908 3210
rect 32 2890 3828 3126
rect 4064 2890 4908 3126
rect 32 2840 4908 2890
rect 3316 -60 4908 -14
rect 3316 -296 3368 -60
rect 3604 -296 4908 -60
rect 3316 -348 4908 -296
use buffer_input  buffer_input_0
timestamp 1654466164
transform 1 0 363 0 1 286
box -356 -286 3286 2508
use buffer_mirror  buffer_mirror_0
timestamp 1654467620
transform 1 0 7 0 1 -3214
box -7 -772 4900 3194
use sky130_fd_pr__res_generic_po_TC8HWG  sky130_fd_pr__res_generic_po_TC8HWG_0
timestamp 1654517990
transform 1 0 4370 0 1 1935
box -516 -589 516 589
use sky130_fd_pr__res_generic_po_TC8HWG  sky130_fd_pr__res_generic_po_TC8HWG_1
timestamp 1654517990
transform 1 0 4370 0 1 863
box -516 -589 516 589
<< labels >>
flabel metal5 s 134 -190 142 -162 0 FreeSans 800 0 0 0 VBIAS
port 0 nsew
flabel metal5 s 132 3160 140 3188 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal3 s 16 1460 24 1488 0 FreeSans 800 0 0 0 IN_P
port 5 nsew
flabel metal3 s 16 1312 24 1340 0 FreeSans 800 0 0 0 IN_N
port 6 nsew
flabel metal5 s 54 -3670 62 -3642 0 FreeSans 800 0 0 0 GND
port 2 nsew
flabel metal3 s 4886 344 4894 372 0 FreeSans 800 0 0 0 OUT_N
port 4 nsew
flabel metal3 s 4892 2414 4900 2442 0 FreeSans 800 0 0 0 OUT_P
port 3 nsew
<< end >>
