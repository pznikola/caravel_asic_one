* NGSPICE file created from vco_pair.ext - technology: sky130B

.subckt sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=1.414e+12p pd=1.066e+07u as=2.828e+12p ps=2.132e+07u w=5.05e+06u l=150000u
X1 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends

.subckt rf_nfet_01v8_aM02W5p00L0p15 DRAIN GATE SOURCE SUBSTRATE
X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 ad=1.414e+12p pd=1.066e+07u as=2.828e+12p ps=2.132e+07u w=5.05e+06u l=150000u
X1 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
.ends

.subckt vco_pair_base sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/DRAIN sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/DRAIN sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/SOURCE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/DRAIN sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/DRAIN sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/DRAIN sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/DRAIN sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/SOURCE
+ rf_nfet_01v8_aM02W5p00L0p15_0/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SOURCE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/SOURCE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/SOURCE
+ rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SOURCE SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/SOURCE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/DRAIN
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13 SUBSTRATE SUBSTRATE SUBSTRATE SUBSTRATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14 SUBSTRATE SUBSTRATE SUBSTRATE SUBSTRATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15 SUBSTRATE SUBSTRATE SUBSTRATE SUBSTRATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16 SUBSTRATE SUBSTRATE SUBSTRATE SUBSTRATE
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xrf_nfet_01v8_aM02W5p00L0p15_0 rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN rf_nfet_01v8_aM02W5p00L0p15_0/GATE
+ rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE SUBSTRATE rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
Xsky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8 sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/DRAIN
+ sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/GATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/SOURCE
+ SUBSTRATE sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15
.ends

.subckt vco_pair GND OUT_P OUT_N
Xvco_pair_base_0 GND OUT_P OUT_P OUT_N GND OUT_P OUT_N GND OUT_P OUT_N OUT_N OUT_N
+ OUT_P OUT_P OUT_N OUT_P GND OUT_N OUT_N GND OUT_P GND OUT_P OUT_P GND OUT_N OUT_P
+ GND GND OUT_N OUT_N GND OUT_N GND OUT_P GND GND OUT_N GND OUT_P GND OUT_P OUT_N
+ vco_pair_base
.ends

