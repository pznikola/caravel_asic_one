* NGSPICE file created from inv_1_pex.ext - technology: sky130B

.subckt inv_1_pex ON OUT VDD GND
X0 VDD.t1 ON.t0 OUT VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=150000u
X1 GND.t1 ON.t1 OUT GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=150000u
C0 VDD ON 0.12fF
C1 VDD OUT 1.48fF
C2 OUT ON 0.03fF
R0 ON.n1 ON.t0 552.693
R1 ON.n1 ON.t1 279.56
R2 ON.n2 ON.n1 119.785
R3 ON.n2 ON.n0 0.078
R4 ON ON.n2 0.002
R5 VDD.n5 VDD.t0 1362.76
R6 VDD.n2 VDD.t1 145.803
R7 VDD.n12 VDD.n11 35.555
R8 VDD.n15 VDD.n14 9.3
R9 VDD.n1 VDD.n0 9.3
R10 VDD VDD.n18 5.716
R11 VDD.n5 VDD.n4 4.68
R12 VDD.n13 VDD.n3 2.007
R13 VDD.n17 VDD.n1 1.65
R14 VDD.n15 VDD.n13 1.003
R15 VDD.n16 VDD.n15 0.535
R16 VDD.n8 VDD.n7 0.501
R17 VDD.n3 VDD.n2 0.125
R18 VDD.n18 VDD.n17 0.05
R19 VDD.n7 VDD.n6 0.032
R20 VDD.n6 VDD.n5 0.032
R21 VDD.n12 VDD.n10 0.008
R22 VDD.n10 VDD.n9 0.007
R23 VDD.n9 VDD.n8 0.007
R24 VDD.n13 VDD.n12 0.007
R25 VDD.n17 VDD.n16 0.003
R26 GND.n7 GND.t0 3941.67
R27 GND.n4 GND.t1 93.671
R28 GND.n5 GND.n1 73.875
R29 GND GND.n9 2.553
R30 GND.n4 GND.n3 2.461
R31 GND.n4 GND.n2 0.656
R32 GND.n5 GND.n4 0.152
R33 GND.n6 GND.n5 0.103
R34 GND.n7 GND.n6 0.049
R35 GND.n9 GND.n0 0.011
R36 GND.n9 GND.n8 0.011
R37 GND.n8 GND.n7 0.003
C3 OUT GND 6.12fF
C4 ON GND 1.34fF
C5 VDD GND 27.13fF
C6 VDD.n0 GND 0.00fF
C7 VDD.n1 GND 0.00fF
C8 VDD.t1 GND 0.05fF $ **FLOATING
C9 VDD.n2 GND 0.01fF
C10 VDD.n3 GND 0.00fF
C11 VDD.t0 GND 0.11fF $ **FLOATING
C12 VDD.n5 GND 0.04fF
C13 VDD.n6 GND 0.00fF
C14 VDD.n7 GND 0.00fF
C15 VDD.n8 GND 0.00fF
C16 VDD.n9 GND 0.00fF
C17 VDD.n10 GND 0.01fF
C18 VDD.n11 GND 0.00fF
C19 VDD.n12 GND 0.00fF
C20 VDD.n13 GND 0.00fF
C21 VDD.n14 GND 0.00fF
C22 VDD.n15 GND 0.00fF
C23 VDD.n16 GND 0.03fF
C24 VDD.n17 GND 0.00fF
C25 VDD.n18 GND 0.56fF
.ends
