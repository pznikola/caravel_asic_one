magic
tech sky130B
magscale 1 2
timestamp 1654466164
<< psubdiff >>
rect -330 2430 2406 2442
rect -330 2396 -284 2430
rect -250 2396 -210 2430
rect -176 2396 -136 2430
rect -102 2396 -62 2430
rect -28 2396 12 2430
rect 46 2396 86 2430
rect 120 2396 160 2430
rect 194 2396 234 2430
rect 268 2396 308 2430
rect 342 2396 382 2430
rect 416 2396 456 2430
rect 490 2396 530 2430
rect 564 2396 604 2430
rect 638 2396 678 2430
rect 712 2396 752 2430
rect 786 2396 826 2430
rect 860 2396 900 2430
rect 934 2396 974 2430
rect 1008 2396 1048 2430
rect 1082 2396 1122 2430
rect 1156 2396 1196 2430
rect 1230 2396 1270 2430
rect 1304 2396 1344 2430
rect 1378 2396 1418 2430
rect 1452 2396 1492 2430
rect 1526 2396 1566 2430
rect 1600 2396 1640 2430
rect 1674 2396 1714 2430
rect 1748 2396 1788 2430
rect 1822 2396 1862 2430
rect 1896 2396 1936 2430
rect 1970 2396 2010 2430
rect 2044 2396 2084 2430
rect 2118 2396 2158 2430
rect 2192 2396 2232 2430
rect 2266 2396 2306 2430
rect 2340 2396 2406 2430
rect -330 2384 2406 2396
rect -330 2256 -272 2384
rect 374 2256 432 2384
rect 940 2256 998 2384
rect 1078 2256 1136 2384
rect 1644 2256 1702 2384
rect 1782 2256 1840 2384
rect 2348 2210 2406 2384
rect -330 1184 -272 1246
rect -330 1150 -318 1184
rect -284 1150 -272 1184
rect -330 1110 -272 1150
rect -330 1076 -318 1110
rect -284 1076 -272 1110
rect -330 1036 -272 1076
rect -330 1002 -318 1036
rect -284 1002 -272 1036
rect -330 982 -272 1002
rect 236 1184 294 1246
rect 236 1150 248 1184
rect 282 1150 294 1184
rect 236 1110 294 1150
rect 236 1076 248 1110
rect 282 1076 294 1110
rect 236 1036 294 1076
rect 236 1002 248 1036
rect 282 1002 294 1036
rect 236 982 294 1002
rect 374 1184 432 1246
rect 374 1150 386 1184
rect 420 1150 432 1184
rect 374 1110 432 1150
rect 374 1076 386 1110
rect 420 1076 432 1110
rect 374 1036 432 1076
rect 374 1002 386 1036
rect 420 1002 432 1036
rect 374 982 432 1002
rect 940 1184 998 1246
rect 940 1150 952 1184
rect 986 1150 998 1184
rect 940 1110 998 1150
rect 940 1076 952 1110
rect 986 1076 998 1110
rect 940 1036 998 1076
rect 940 1002 952 1036
rect 986 1002 998 1036
rect 940 982 998 1002
rect 1078 1184 1136 1246
rect 1078 1150 1090 1184
rect 1124 1150 1136 1184
rect 1078 1110 1136 1150
rect 1078 1076 1090 1110
rect 1124 1076 1136 1110
rect 1078 1036 1136 1076
rect 1078 1002 1090 1036
rect 1124 1002 1136 1036
rect 1078 982 1136 1002
rect 1644 1184 1702 1246
rect 1644 1150 1656 1184
rect 1690 1150 1702 1184
rect 1644 1110 1702 1150
rect 1644 1076 1656 1110
rect 1690 1076 1702 1110
rect 1644 1036 1702 1076
rect 1644 1002 1656 1036
rect 1690 1002 1702 1036
rect 1644 982 1702 1002
rect 1782 1184 1840 1246
rect 1782 1150 1794 1184
rect 1828 1150 1840 1184
rect 1782 1110 1840 1150
rect 1782 1076 1794 1110
rect 1828 1076 1840 1110
rect 1782 1036 1840 1076
rect 1782 1002 1794 1036
rect 1828 1002 1840 1036
rect 1782 982 1840 1002
rect 2348 1184 2406 1246
rect 2348 1150 2360 1184
rect 2394 1150 2406 1184
rect 2348 1110 2406 1150
rect 2348 1076 2360 1110
rect 2394 1076 2406 1110
rect 2348 1036 2406 1076
rect 2348 1002 2360 1036
rect 2394 1002 2406 1036
rect 2348 982 2406 1002
rect -330 -148 -272 -28
rect 374 -148 432 -28
rect 940 -148 998 -28
rect 1078 -148 1136 -28
rect 1644 -148 1702 -28
rect 1782 -148 1840 -28
rect 2348 -148 2406 18
rect -330 -168 2406 -148
rect -330 -202 -284 -168
rect -250 -202 -210 -168
rect -176 -202 -136 -168
rect -102 -202 -62 -168
rect -28 -202 12 -168
rect 46 -202 86 -168
rect 120 -202 160 -168
rect 194 -202 234 -168
rect 268 -202 308 -168
rect 342 -202 382 -168
rect 416 -202 456 -168
rect 490 -202 530 -168
rect 564 -202 604 -168
rect 638 -202 678 -168
rect 712 -202 752 -168
rect 786 -202 826 -168
rect 860 -202 900 -168
rect 934 -202 974 -168
rect 1008 -202 1048 -168
rect 1082 -202 1122 -168
rect 1156 -202 1196 -168
rect 1230 -202 1270 -168
rect 1304 -202 1344 -168
rect 1378 -202 1418 -168
rect 1452 -202 1492 -168
rect 1526 -202 1566 -168
rect 1600 -202 1640 -168
rect 1674 -202 1714 -168
rect 1748 -202 1788 -168
rect 1822 -202 1862 -168
rect 1896 -202 1936 -168
rect 1970 -202 2010 -168
rect 2044 -202 2084 -168
rect 2118 -202 2158 -168
rect 2192 -202 2232 -168
rect 2266 -202 2306 -168
rect 2340 -202 2406 -168
rect -330 -214 2406 -202
<< psubdiffcont >>
rect -284 2396 -250 2430
rect -210 2396 -176 2430
rect -136 2396 -102 2430
rect -62 2396 -28 2430
rect 12 2396 46 2430
rect 86 2396 120 2430
rect 160 2396 194 2430
rect 234 2396 268 2430
rect 308 2396 342 2430
rect 382 2396 416 2430
rect 456 2396 490 2430
rect 530 2396 564 2430
rect 604 2396 638 2430
rect 678 2396 712 2430
rect 752 2396 786 2430
rect 826 2396 860 2430
rect 900 2396 934 2430
rect 974 2396 1008 2430
rect 1048 2396 1082 2430
rect 1122 2396 1156 2430
rect 1196 2396 1230 2430
rect 1270 2396 1304 2430
rect 1344 2396 1378 2430
rect 1418 2396 1452 2430
rect 1492 2396 1526 2430
rect 1566 2396 1600 2430
rect 1640 2396 1674 2430
rect 1714 2396 1748 2430
rect 1788 2396 1822 2430
rect 1862 2396 1896 2430
rect 1936 2396 1970 2430
rect 2010 2396 2044 2430
rect 2084 2396 2118 2430
rect 2158 2396 2192 2430
rect 2232 2396 2266 2430
rect 2306 2396 2340 2430
rect -318 1150 -284 1184
rect -318 1076 -284 1110
rect -318 1002 -284 1036
rect 248 1150 282 1184
rect 248 1076 282 1110
rect 248 1002 282 1036
rect 386 1150 420 1184
rect 386 1076 420 1110
rect 386 1002 420 1036
rect 952 1150 986 1184
rect 952 1076 986 1110
rect 952 1002 986 1036
rect 1090 1150 1124 1184
rect 1090 1076 1124 1110
rect 1090 1002 1124 1036
rect 1656 1150 1690 1184
rect 1656 1076 1690 1110
rect 1656 1002 1690 1036
rect 1794 1150 1828 1184
rect 1794 1076 1828 1110
rect 1794 1002 1828 1036
rect 2360 1150 2394 1184
rect 2360 1076 2394 1110
rect 2360 1002 2394 1036
rect -284 -202 -250 -168
rect -210 -202 -176 -168
rect -136 -202 -102 -168
rect -62 -202 -28 -168
rect 12 -202 46 -168
rect 86 -202 120 -168
rect 160 -202 194 -168
rect 234 -202 268 -168
rect 308 -202 342 -168
rect 382 -202 416 -168
rect 456 -202 490 -168
rect 530 -202 564 -168
rect 604 -202 638 -168
rect 678 -202 712 -168
rect 752 -202 786 -168
rect 826 -202 860 -168
rect 900 -202 934 -168
rect 974 -202 1008 -168
rect 1048 -202 1082 -168
rect 1122 -202 1156 -168
rect 1196 -202 1230 -168
rect 1270 -202 1304 -168
rect 1344 -202 1378 -168
rect 1418 -202 1452 -168
rect 1492 -202 1526 -168
rect 1566 -202 1600 -168
rect 1640 -202 1674 -168
rect 1714 -202 1748 -168
rect 1788 -202 1822 -168
rect 1862 -202 1896 -168
rect 1936 -202 1970 -168
rect 2010 -202 2044 -168
rect 2084 -202 2118 -168
rect 2158 -202 2192 -168
rect 2232 -202 2266 -168
rect 2306 -202 2340 -168
<< locali >>
rect -318 2236 -284 2430
rect -250 2396 -210 2430
rect -176 2396 -136 2430
rect -102 2396 -62 2430
rect -28 2396 12 2430
rect 46 2396 86 2430
rect 120 2396 160 2430
rect 194 2396 234 2430
rect 268 2396 308 2430
rect 342 2396 382 2430
rect 416 2396 456 2430
rect 490 2396 530 2430
rect 564 2396 604 2430
rect 638 2396 678 2430
rect 712 2396 752 2430
rect 786 2396 826 2430
rect 860 2396 900 2430
rect 934 2396 974 2430
rect 1008 2396 1048 2430
rect 1082 2396 1122 2430
rect 1156 2396 1196 2430
rect 1230 2396 1270 2430
rect 1304 2396 1344 2430
rect 1378 2396 1418 2430
rect 1452 2396 1492 2430
rect 1526 2396 1566 2430
rect 1600 2396 1640 2430
rect 1674 2396 1714 2430
rect 1748 2396 1788 2430
rect 1822 2396 1862 2430
rect 1896 2396 1936 2430
rect 1970 2396 2010 2430
rect 2044 2396 2084 2430
rect 2118 2396 2158 2430
rect 2192 2396 2232 2430
rect 2266 2396 2306 2430
rect 2340 2396 2394 2430
rect 386 2236 420 2396
rect 952 2236 986 2396
rect 1090 2236 1124 2396
rect 1656 2236 1690 2396
rect 1794 2236 1828 2396
rect 2360 2236 2394 2396
rect -318 1184 -284 1266
rect -318 1110 -284 1150
rect -318 1036 -284 1076
rect -318 962 -284 1002
rect 248 1184 282 1266
rect 248 1110 282 1150
rect 248 1036 282 1076
rect 248 962 282 1002
rect 386 1184 420 1266
rect 386 1110 420 1150
rect 386 1036 420 1076
rect 386 962 420 1002
rect 952 1184 986 1266
rect 952 1110 986 1150
rect 952 1036 986 1076
rect 952 962 986 1002
rect 1090 1184 1124 1266
rect 1090 1110 1124 1150
rect 1090 1036 1124 1076
rect 1090 962 1124 1002
rect 1656 1184 1690 1266
rect 1656 1110 1690 1150
rect 1656 1036 1690 1076
rect 1656 962 1690 1002
rect 1794 1184 1828 1266
rect 1794 1110 1828 1150
rect 1794 1036 1828 1076
rect 1794 962 1828 1002
rect 2360 1184 2394 1266
rect 2360 1110 2394 1150
rect 2360 1036 2394 1076
rect 2360 962 2394 1002
rect -318 -202 -284 0
rect 386 -168 420 -8
rect 952 -168 986 -8
rect 1090 -168 1124 -8
rect 1656 -168 1690 -8
rect 1794 -168 1828 -8
rect 2360 -168 2394 0
rect -250 -202 -210 -168
rect -176 -202 -136 -168
rect -102 -202 -62 -168
rect -28 -202 12 -168
rect 46 -202 86 -168
rect 120 -202 160 -168
rect 194 -202 234 -168
rect 268 -202 308 -168
rect 342 -202 382 -168
rect 416 -202 456 -168
rect 490 -202 530 -168
rect 564 -202 604 -168
rect 638 -202 678 -168
rect 712 -202 752 -168
rect 786 -202 826 -168
rect 860 -202 900 -168
rect 934 -202 974 -168
rect 1008 -202 1048 -168
rect 1082 -202 1122 -168
rect 1156 -202 1196 -168
rect 1230 -202 1270 -168
rect 1304 -202 1344 -168
rect 1378 -202 1418 -168
rect 1452 -202 1492 -168
rect 1526 -202 1566 -168
rect 1600 -202 1640 -168
rect 1674 -202 1714 -168
rect 1748 -202 1788 -168
rect 1822 -202 1862 -168
rect 1896 -202 1936 -168
rect 1970 -202 2010 -168
rect 2044 -202 2084 -168
rect 2118 -202 2158 -168
rect 2192 -202 2232 -168
rect 2266 -202 2306 -168
rect 2340 -202 2394 -168
<< viali >>
rect -284 2396 -250 2430
rect -210 2396 -176 2430
rect -136 2396 -102 2430
rect -62 2396 -28 2430
rect 12 2396 46 2430
rect 86 2396 120 2430
rect 160 2396 194 2430
rect 234 2396 268 2430
rect 308 2396 342 2430
rect 382 2396 416 2430
rect 456 2396 490 2430
rect 530 2396 564 2430
rect 604 2396 638 2430
rect 678 2396 712 2430
rect 752 2396 786 2430
rect 826 2396 860 2430
rect 900 2396 934 2430
rect 974 2396 1008 2430
rect 1048 2396 1082 2430
rect 1122 2396 1156 2430
rect 1196 2396 1230 2430
rect 1270 2396 1304 2430
rect 1344 2396 1378 2430
rect 1418 2396 1452 2430
rect 1492 2396 1526 2430
rect 1566 2396 1600 2430
rect 1640 2396 1674 2430
rect 1714 2396 1748 2430
rect 1788 2396 1822 2430
rect 1862 2396 1896 2430
rect 1936 2396 1970 2430
rect 2010 2396 2044 2430
rect 2084 2396 2118 2430
rect 2158 2396 2192 2430
rect 2232 2396 2266 2430
rect 2306 2396 2340 2430
rect -318 1150 -284 1184
rect -318 1076 -284 1110
rect -318 1002 -284 1036
rect 248 1150 282 1184
rect 248 1076 282 1110
rect 248 1002 282 1036
rect 386 1150 420 1184
rect 386 1076 420 1110
rect 386 1002 420 1036
rect 952 1150 986 1184
rect 952 1076 986 1110
rect 952 1002 986 1036
rect 1090 1150 1124 1184
rect 1090 1076 1124 1110
rect 1090 1002 1124 1036
rect 1656 1150 1690 1184
rect 1656 1076 1690 1110
rect 1656 1002 1690 1036
rect 1794 1150 1828 1184
rect 1794 1076 1828 1110
rect 1794 1002 1828 1036
rect 2360 1150 2394 1184
rect 2360 1076 2394 1110
rect 2360 1002 2394 1036
rect -284 -202 -250 -168
rect -210 -202 -176 -168
rect -136 -202 -102 -168
rect -62 -202 -28 -168
rect 12 -202 46 -168
rect 86 -202 120 -168
rect 160 -202 194 -168
rect 234 -202 268 -168
rect 308 -202 342 -168
rect 382 -202 416 -168
rect 456 -202 490 -168
rect 530 -202 564 -168
rect 604 -202 638 -168
rect 678 -202 712 -168
rect 752 -202 786 -168
rect 826 -202 860 -168
rect 900 -202 934 -168
rect 974 -202 1008 -168
rect 1048 -202 1082 -168
rect 1122 -202 1156 -168
rect 1196 -202 1230 -168
rect 1270 -202 1304 -168
rect 1344 -202 1378 -168
rect 1418 -202 1452 -168
rect 1492 -202 1526 -168
rect 1566 -202 1600 -168
rect 1640 -202 1674 -168
rect 1714 -202 1748 -168
rect 1788 -202 1822 -168
rect 1862 -202 1896 -168
rect 1936 -202 1970 -168
rect 2010 -202 2044 -168
rect 2084 -202 2118 -168
rect 2158 -202 2192 -168
rect 2232 -202 2266 -168
rect 2306 -202 2340 -168
<< metal1 >>
rect -330 2430 2406 2442
rect -330 2396 -284 2430
rect -250 2396 -210 2430
rect -176 2396 -136 2430
rect -102 2396 -62 2430
rect -28 2396 12 2430
rect 46 2396 86 2430
rect 120 2396 160 2430
rect 194 2396 234 2430
rect 268 2396 308 2430
rect 342 2396 382 2430
rect 416 2396 456 2430
rect 490 2396 530 2430
rect 564 2396 604 2430
rect 638 2396 678 2430
rect 712 2396 752 2430
rect 786 2396 826 2430
rect 860 2396 900 2430
rect 934 2396 974 2430
rect 1008 2396 1048 2430
rect 1082 2396 1122 2430
rect 1156 2396 1196 2430
rect 1230 2396 1270 2430
rect 1304 2396 1344 2430
rect 1378 2396 1418 2430
rect 1452 2396 1492 2430
rect 1526 2396 1566 2430
rect 1600 2396 1640 2430
rect 1674 2396 1714 2430
rect 1748 2396 1788 2430
rect 1822 2396 1862 2430
rect 1896 2396 1936 2430
rect 1970 2396 2010 2430
rect 2044 2396 2084 2430
rect 2118 2396 2158 2430
rect 2192 2396 2232 2430
rect 2266 2396 2306 2430
rect 2340 2396 2406 2430
rect -330 2376 2406 2396
rect -330 2282 294 2376
rect -330 2248 -272 2282
rect -216 2248 -164 2282
rect -130 2248 -78 2282
rect -44 2248 8 2282
rect 42 2248 94 2282
rect 128 2248 180 2282
rect 236 2248 294 2282
rect 374 2244 432 2376
rect 512 2340 860 2348
rect 512 2288 538 2340
rect 590 2288 602 2340
rect 654 2288 666 2340
rect 718 2288 730 2340
rect 782 2288 794 2340
rect 846 2288 860 2340
rect 512 2282 860 2288
rect 940 2244 998 2376
rect 1078 2244 1136 2376
rect 1216 2340 1564 2348
rect 1216 2288 1242 2340
rect 1294 2288 1306 2340
rect 1358 2288 1370 2340
rect 1422 2288 1434 2340
rect 1486 2288 1498 2340
rect 1550 2288 1564 2340
rect 1216 2282 1564 2288
rect 1644 2244 1702 2376
rect 1782 2282 2406 2376
rect 1782 2244 1840 2282
rect 1896 2248 1948 2282
rect 1982 2248 2034 2282
rect 2068 2248 2120 2282
rect 2154 2248 2206 2282
rect 2240 2248 2292 2282
rect 2348 2248 2406 2282
rect -330 1220 -272 1254
rect -216 1220 -164 1254
rect -130 1220 -78 1254
rect -44 1220 8 1254
rect 42 1220 94 1254
rect 128 1220 180 1254
rect 236 1220 294 1254
rect -330 1184 294 1220
rect -330 1150 -318 1184
rect -284 1154 248 1184
rect -284 1150 -272 1154
rect -330 1110 -272 1150
rect -330 1076 -318 1110
rect -284 1076 -272 1110
rect -330 1074 -272 1076
rect 236 1150 248 1154
rect 282 1150 294 1184
rect 236 1110 294 1150
rect 236 1076 248 1110
rect 282 1076 294 1110
rect 236 1074 294 1076
rect -330 1036 294 1074
rect -330 1002 -318 1036
rect -284 1008 248 1036
rect -284 1002 -272 1008
rect -330 974 -272 1002
rect -216 974 -164 1008
rect -130 974 -78 1008
rect -44 974 8 1008
rect 42 974 94 1008
rect 128 974 180 1008
rect 236 1002 248 1008
rect 282 1002 294 1036
rect 236 974 294 1002
rect 374 1184 432 1254
rect 374 1150 386 1184
rect 420 1150 432 1184
rect 512 1212 860 1220
rect 512 1160 518 1212
rect 570 1160 586 1212
rect 638 1160 658 1212
rect 710 1160 730 1212
rect 782 1160 802 1212
rect 854 1160 860 1212
rect 512 1154 860 1160
rect 940 1184 998 1254
rect 374 1110 432 1150
rect 374 1076 386 1110
rect 420 1076 432 1110
rect 374 1036 432 1076
rect 940 1150 952 1184
rect 986 1150 998 1184
rect 940 1110 998 1150
rect 940 1076 952 1110
rect 986 1076 998 1110
rect 374 1002 386 1036
rect 420 1002 432 1036
rect 512 1066 860 1074
rect 512 1014 518 1066
rect 570 1014 586 1066
rect 638 1014 658 1066
rect 710 1014 730 1066
rect 782 1014 802 1066
rect 854 1014 860 1066
rect 512 1008 860 1014
rect 940 1036 998 1076
rect 374 974 432 1002
rect 940 1002 952 1036
rect 986 1002 998 1036
rect 940 974 998 1002
rect 1078 1184 1136 1254
rect 1078 1150 1090 1184
rect 1124 1150 1136 1184
rect 1216 1212 1564 1220
rect 1216 1160 1222 1212
rect 1274 1160 1290 1212
rect 1342 1160 1362 1212
rect 1414 1160 1434 1212
rect 1486 1160 1506 1212
rect 1558 1160 1564 1212
rect 1216 1154 1564 1160
rect 1644 1184 1702 1254
rect 1078 1110 1136 1150
rect 1078 1076 1090 1110
rect 1124 1076 1136 1110
rect 1078 1036 1136 1076
rect 1644 1150 1656 1184
rect 1690 1150 1702 1184
rect 1644 1110 1702 1150
rect 1644 1076 1656 1110
rect 1690 1076 1702 1110
rect 1078 1002 1090 1036
rect 1124 1002 1136 1036
rect 1216 1066 1564 1074
rect 1216 1014 1224 1066
rect 1276 1014 1290 1066
rect 1342 1014 1362 1066
rect 1414 1014 1434 1066
rect 1486 1014 1506 1066
rect 1558 1014 1564 1066
rect 1216 1008 1564 1014
rect 1644 1036 1702 1076
rect 1078 974 1136 1002
rect 1644 1002 1656 1036
rect 1690 1002 1702 1036
rect 1644 974 1702 1002
rect 1782 1220 1840 1254
rect 1896 1220 1948 1254
rect 1982 1220 2034 1254
rect 2068 1220 2120 1254
rect 2154 1220 2206 1254
rect 2240 1220 2292 1254
rect 2348 1220 2406 1254
rect 1782 1184 2406 1220
rect 1782 1150 1794 1184
rect 1828 1154 2360 1184
rect 1828 1150 1840 1154
rect 1782 1110 1840 1150
rect 1782 1076 1794 1110
rect 1828 1076 1840 1110
rect 1782 1074 1840 1076
rect 2348 1150 2360 1154
rect 2394 1150 2406 1184
rect 2348 1110 2406 1150
rect 2348 1076 2360 1110
rect 2394 1076 2406 1110
rect 2348 1074 2406 1076
rect 1782 1036 2406 1074
rect 1782 1002 1794 1036
rect 1828 1008 2360 1036
rect 1828 1002 1840 1008
rect 1782 974 1840 1002
rect 1896 974 1948 1008
rect 1982 974 2034 1008
rect 2068 974 2120 1008
rect 2154 974 2206 1008
rect 2240 974 2292 1008
rect 2348 1002 2360 1008
rect 2394 1002 2406 1036
rect 2348 974 2406 1002
rect 236 -20 284 -6
rect -330 -54 -272 -20
rect -216 -54 -164 -20
rect -130 -54 -78 -20
rect -44 -54 8 -20
rect 42 -54 94 -20
rect 128 -54 180 -20
rect 236 -54 294 -20
rect -330 -148 294 -54
rect 374 -148 432 -20
rect 512 -60 860 -54
rect 512 -112 538 -60
rect 590 -112 602 -60
rect 654 -112 666 -60
rect 718 -112 730 -60
rect 782 -112 794 -60
rect 846 -112 860 -60
rect 512 -120 860 -112
rect 940 -148 998 -20
rect 1078 -148 1136 -20
rect 1216 -60 1564 -54
rect 1216 -112 1242 -60
rect 1294 -112 1306 -60
rect 1358 -112 1370 -60
rect 1422 -112 1434 -60
rect 1486 -112 1498 -60
rect 1550 -112 1564 -60
rect 1216 -120 1564 -112
rect 1644 -148 1702 -20
rect 1782 -54 1840 -20
rect 1896 -54 1948 -20
rect 1982 -54 2034 -20
rect 2068 -54 2120 -20
rect 2154 -54 2206 -20
rect 2240 -54 2292 -20
rect 2348 -54 2406 -20
rect 1782 -148 2406 -54
rect -330 -168 2406 -148
rect -330 -202 -284 -168
rect -250 -202 -210 -168
rect -176 -202 -136 -168
rect -102 -202 -62 -168
rect -28 -202 12 -168
rect 46 -202 86 -168
rect 120 -202 160 -168
rect 194 -202 234 -168
rect 268 -202 308 -168
rect 342 -202 382 -168
rect 416 -202 456 -168
rect 490 -202 530 -168
rect 564 -202 604 -168
rect 638 -202 678 -168
rect 712 -202 752 -168
rect 786 -202 826 -168
rect 860 -202 900 -168
rect 934 -202 974 -168
rect 1008 -202 1048 -168
rect 1082 -202 1122 -168
rect 1156 -202 1196 -168
rect 1230 -202 1270 -168
rect 1304 -202 1344 -168
rect 1378 -202 1418 -168
rect 1452 -202 1492 -168
rect 1526 -202 1566 -168
rect 1600 -202 1640 -168
rect 1674 -202 1714 -168
rect 1748 -202 1788 -168
rect 1822 -202 1862 -168
rect 1896 -202 1936 -168
rect 1970 -202 2010 -168
rect 2044 -202 2084 -168
rect 2118 -202 2158 -168
rect 2192 -202 2232 -168
rect 2266 -202 2306 -168
rect 2340 -202 2406 -168
rect -330 -214 2406 -202
<< via1 >>
rect 538 2288 590 2340
rect 602 2288 654 2340
rect 666 2288 718 2340
rect 730 2288 782 2340
rect 794 2288 846 2340
rect 1242 2288 1294 2340
rect 1306 2288 1358 2340
rect 1370 2288 1422 2340
rect 1434 2288 1486 2340
rect 1498 2288 1550 2340
rect 518 1160 570 1212
rect 586 1160 638 1212
rect 658 1160 710 1212
rect 730 1160 782 1212
rect 802 1160 854 1212
rect 518 1014 570 1066
rect 586 1014 638 1066
rect 658 1014 710 1066
rect 730 1014 782 1066
rect 802 1014 854 1066
rect 1222 1160 1274 1212
rect 1290 1160 1342 1212
rect 1362 1160 1414 1212
rect 1434 1160 1486 1212
rect 1506 1160 1558 1212
rect 1224 1014 1276 1066
rect 1290 1014 1342 1066
rect 1362 1014 1414 1066
rect 1434 1014 1486 1066
rect 1506 1014 1558 1066
rect 538 -112 590 -60
rect 602 -112 654 -60
rect 666 -112 718 -60
rect 730 -112 782 -60
rect 794 -112 846 -60
rect 1242 -112 1294 -60
rect 1306 -112 1358 -60
rect 1370 -112 1422 -60
rect 1434 -112 1486 -60
rect 1498 -112 1550 -60
<< metal2 >>
rect 512 2370 860 2378
rect 512 2340 544 2370
rect 600 2340 624 2370
rect 680 2340 704 2370
rect 760 2340 784 2370
rect 840 2340 860 2370
rect 512 2288 538 2340
rect 600 2314 602 2340
rect 782 2314 784 2340
rect 590 2288 602 2314
rect 654 2288 666 2314
rect 718 2288 730 2314
rect 782 2288 794 2314
rect 846 2288 860 2340
rect 512 2282 860 2288
rect 1216 2370 1564 2378
rect 1216 2340 1248 2370
rect 1304 2340 1328 2370
rect 1384 2340 1408 2370
rect 1464 2340 1488 2370
rect 1544 2340 1564 2370
rect 1216 2288 1242 2340
rect 1304 2314 1306 2340
rect 1486 2314 1488 2340
rect 1294 2288 1306 2314
rect 1358 2288 1370 2314
rect 1422 2288 1434 2314
rect 1486 2288 1498 2314
rect 1550 2288 1564 2340
rect 1216 2282 1564 2288
rect 348 2216 1024 2248
rect 348 2160 378 2216
rect 434 2160 458 2216
rect 514 2160 538 2216
rect 594 2160 618 2216
rect 674 2160 698 2216
rect 754 2160 778 2216
rect 834 2160 858 2216
rect 914 2160 938 2216
rect 994 2160 1024 2216
rect 348 2136 1024 2160
rect 348 2080 378 2136
rect 434 2080 458 2136
rect 514 2080 538 2136
rect 594 2080 618 2136
rect 674 2080 698 2136
rect 754 2080 778 2136
rect 834 2080 858 2136
rect 914 2080 938 2136
rect 994 2080 1024 2136
rect 348 2048 1024 2080
rect 1052 1944 1728 1976
rect 1052 1888 1082 1944
rect 1138 1888 1162 1944
rect 1218 1888 1242 1944
rect 1298 1888 1322 1944
rect 1378 1888 1402 1944
rect 1458 1888 1482 1944
rect 1538 1888 1562 1944
rect 1618 1888 1642 1944
rect 1698 1888 1728 1944
rect 1052 1864 1728 1888
rect 1052 1808 1082 1864
rect 1138 1808 1162 1864
rect 1218 1808 1242 1864
rect 1298 1808 1322 1864
rect 1378 1808 1402 1864
rect 1458 1808 1482 1864
rect 1538 1808 1562 1864
rect 1618 1808 1642 1864
rect 1698 1808 1728 1864
rect 1052 1776 1728 1808
rect 374 1588 998 1638
rect 374 1532 458 1588
rect 514 1532 538 1588
rect 594 1532 618 1588
rect 674 1532 698 1588
rect 754 1532 778 1588
rect 834 1532 858 1588
rect 914 1532 998 1588
rect 374 1508 998 1532
rect 374 1452 458 1508
rect 514 1452 538 1508
rect 594 1452 618 1508
rect 674 1452 698 1508
rect 754 1452 778 1508
rect 834 1452 858 1508
rect 914 1452 998 1508
rect 374 1424 998 1452
rect 374 1368 458 1424
rect 514 1368 538 1424
rect 594 1368 618 1424
rect 674 1368 698 1424
rect 754 1368 778 1424
rect 834 1368 858 1424
rect 914 1368 998 1424
rect 374 1318 998 1368
rect 1078 1588 1702 1638
rect 1078 1532 1162 1588
rect 1218 1532 1242 1588
rect 1298 1532 1322 1588
rect 1378 1532 1402 1588
rect 1458 1532 1482 1588
rect 1538 1532 1562 1588
rect 1618 1532 1702 1588
rect 1078 1508 1702 1532
rect 1078 1452 1162 1508
rect 1218 1452 1242 1508
rect 1298 1452 1322 1508
rect 1378 1452 1402 1508
rect 1458 1452 1482 1508
rect 1538 1452 1562 1508
rect 1618 1452 1702 1508
rect 1078 1424 1702 1452
rect 1078 1368 1162 1424
rect 1218 1368 1242 1424
rect 1298 1368 1322 1424
rect 1378 1368 1402 1424
rect 1458 1368 1482 1424
rect 1538 1368 1562 1424
rect 1618 1368 1702 1424
rect 1078 1318 1702 1368
rect 512 1220 860 1222
rect 512 1216 1070 1220
rect 512 1212 522 1216
rect 578 1212 612 1216
rect 668 1212 702 1216
rect 758 1212 794 1216
rect 850 1212 1070 1216
rect 512 1160 518 1212
rect 578 1160 586 1212
rect 782 1160 794 1212
rect 854 1160 1070 1212
rect 512 1154 1070 1160
rect 1216 1216 1564 1222
rect 1216 1212 1226 1216
rect 1282 1212 1316 1216
rect 1372 1212 1406 1216
rect 1462 1212 1498 1216
rect 1554 1212 1564 1216
rect 1216 1160 1222 1212
rect 1282 1160 1290 1212
rect 1486 1160 1498 1212
rect 1558 1160 1564 1212
rect 1216 1154 1564 1160
rect 1004 1074 1070 1154
rect 512 1068 860 1074
rect 512 1066 522 1068
rect 578 1066 612 1068
rect 668 1066 702 1068
rect 758 1066 794 1068
rect 850 1066 860 1068
rect 512 1014 518 1066
rect 578 1014 586 1066
rect 782 1014 794 1066
rect 854 1014 860 1066
rect 512 1012 522 1014
rect 578 1012 612 1014
rect 668 1012 702 1014
rect 758 1012 794 1014
rect 850 1012 860 1014
rect 512 1006 860 1012
rect 1004 1066 1564 1074
rect 1004 1014 1224 1066
rect 1276 1014 1290 1066
rect 1342 1014 1362 1066
rect 1414 1014 1434 1066
rect 1486 1014 1506 1066
rect 1558 1014 1564 1066
rect 1004 1008 1564 1014
rect 374 860 998 910
rect 374 804 458 860
rect 514 804 538 860
rect 594 804 618 860
rect 674 804 698 860
rect 754 804 778 860
rect 834 804 858 860
rect 914 804 998 860
rect 374 780 998 804
rect 374 724 458 780
rect 514 724 538 780
rect 594 724 618 780
rect 674 724 698 780
rect 754 724 778 780
rect 834 724 858 780
rect 914 724 998 780
rect 374 696 998 724
rect 374 640 458 696
rect 514 640 538 696
rect 594 640 618 696
rect 674 640 698 696
rect 754 640 778 696
rect 834 640 858 696
rect 914 640 998 696
rect 374 590 998 640
rect 1078 860 1702 910
rect 1078 804 1162 860
rect 1218 804 1242 860
rect 1298 804 1322 860
rect 1378 804 1402 860
rect 1458 804 1482 860
rect 1538 804 1562 860
rect 1618 804 1702 860
rect 1078 780 1702 804
rect 1078 724 1162 780
rect 1218 724 1242 780
rect 1298 724 1322 780
rect 1378 724 1402 780
rect 1458 724 1482 780
rect 1538 724 1562 780
rect 1618 724 1702 780
rect 1078 696 1702 724
rect 1078 640 1162 696
rect 1218 640 1242 696
rect 1298 640 1322 696
rect 1378 640 1402 696
rect 1458 640 1482 696
rect 1538 640 1562 696
rect 1618 640 1702 696
rect 1078 590 1702 640
rect 348 420 1024 452
rect 348 364 378 420
rect 434 364 458 420
rect 514 364 538 420
rect 594 364 618 420
rect 674 364 698 420
rect 754 364 778 420
rect 834 364 858 420
rect 914 364 938 420
rect 994 364 1024 420
rect 348 340 1024 364
rect 348 284 378 340
rect 434 284 458 340
rect 514 284 538 340
rect 594 284 618 340
rect 674 284 698 340
rect 754 284 778 340
rect 834 284 858 340
rect 914 284 938 340
rect 994 284 1024 340
rect 348 252 1024 284
rect 1052 148 1728 180
rect 1052 92 1082 148
rect 1138 92 1162 148
rect 1218 92 1242 148
rect 1298 92 1322 148
rect 1378 92 1402 148
rect 1458 92 1482 148
rect 1538 92 1562 148
rect 1618 92 1642 148
rect 1698 92 1728 148
rect 1052 68 1728 92
rect 1052 12 1082 68
rect 1138 12 1162 68
rect 1218 12 1242 68
rect 1298 12 1322 68
rect 1378 12 1402 68
rect 1458 12 1482 68
rect 1538 12 1562 68
rect 1618 12 1642 68
rect 1698 12 1728 68
rect 1052 -20 1728 12
rect 512 -60 860 -54
rect 512 -112 538 -60
rect 590 -86 602 -60
rect 654 -86 666 -60
rect 718 -86 730 -60
rect 782 -86 794 -60
rect 600 -112 602 -86
rect 782 -112 784 -86
rect 846 -112 860 -60
rect 512 -142 544 -112
rect 600 -142 624 -112
rect 680 -142 704 -112
rect 760 -142 784 -112
rect 840 -142 860 -112
rect 512 -150 860 -142
rect 1216 -60 1564 -54
rect 1216 -112 1242 -60
rect 1294 -86 1306 -60
rect 1358 -86 1370 -60
rect 1422 -86 1434 -60
rect 1486 -86 1498 -60
rect 1304 -112 1306 -86
rect 1486 -112 1488 -86
rect 1550 -112 1564 -60
rect 1216 -142 1248 -112
rect 1304 -142 1328 -112
rect 1384 -142 1408 -112
rect 1464 -142 1488 -112
rect 1544 -142 1564 -112
rect 1216 -150 1564 -142
<< via2 >>
rect 544 2340 600 2370
rect 624 2340 680 2370
rect 704 2340 760 2370
rect 784 2340 840 2370
rect 544 2314 590 2340
rect 590 2314 600 2340
rect 624 2314 654 2340
rect 654 2314 666 2340
rect 666 2314 680 2340
rect 704 2314 718 2340
rect 718 2314 730 2340
rect 730 2314 760 2340
rect 784 2314 794 2340
rect 794 2314 840 2340
rect 1248 2340 1304 2370
rect 1328 2340 1384 2370
rect 1408 2340 1464 2370
rect 1488 2340 1544 2370
rect 1248 2314 1294 2340
rect 1294 2314 1304 2340
rect 1328 2314 1358 2340
rect 1358 2314 1370 2340
rect 1370 2314 1384 2340
rect 1408 2314 1422 2340
rect 1422 2314 1434 2340
rect 1434 2314 1464 2340
rect 1488 2314 1498 2340
rect 1498 2314 1544 2340
rect 378 2160 434 2216
rect 458 2160 514 2216
rect 538 2160 594 2216
rect 618 2160 674 2216
rect 698 2160 754 2216
rect 778 2160 834 2216
rect 858 2160 914 2216
rect 938 2160 994 2216
rect 378 2080 434 2136
rect 458 2080 514 2136
rect 538 2080 594 2136
rect 618 2080 674 2136
rect 698 2080 754 2136
rect 778 2080 834 2136
rect 858 2080 914 2136
rect 938 2080 994 2136
rect 1082 1888 1138 1944
rect 1162 1888 1218 1944
rect 1242 1888 1298 1944
rect 1322 1888 1378 1944
rect 1402 1888 1458 1944
rect 1482 1888 1538 1944
rect 1562 1888 1618 1944
rect 1642 1888 1698 1944
rect 1082 1808 1138 1864
rect 1162 1808 1218 1864
rect 1242 1808 1298 1864
rect 1322 1808 1378 1864
rect 1402 1808 1458 1864
rect 1482 1808 1538 1864
rect 1562 1808 1618 1864
rect 1642 1808 1698 1864
rect 458 1532 514 1588
rect 538 1532 594 1588
rect 618 1532 674 1588
rect 698 1532 754 1588
rect 778 1532 834 1588
rect 858 1532 914 1588
rect 458 1452 514 1508
rect 538 1452 594 1508
rect 618 1452 674 1508
rect 698 1452 754 1508
rect 778 1452 834 1508
rect 858 1452 914 1508
rect 458 1368 514 1424
rect 538 1368 594 1424
rect 618 1368 674 1424
rect 698 1368 754 1424
rect 778 1368 834 1424
rect 858 1368 914 1424
rect 1162 1532 1218 1588
rect 1242 1532 1298 1588
rect 1322 1532 1378 1588
rect 1402 1532 1458 1588
rect 1482 1532 1538 1588
rect 1562 1532 1618 1588
rect 1162 1452 1218 1508
rect 1242 1452 1298 1508
rect 1322 1452 1378 1508
rect 1402 1452 1458 1508
rect 1482 1452 1538 1508
rect 1562 1452 1618 1508
rect 1162 1368 1218 1424
rect 1242 1368 1298 1424
rect 1322 1368 1378 1424
rect 1402 1368 1458 1424
rect 1482 1368 1538 1424
rect 1562 1368 1618 1424
rect 522 1212 578 1216
rect 612 1212 668 1216
rect 702 1212 758 1216
rect 794 1212 850 1216
rect 522 1160 570 1212
rect 570 1160 578 1212
rect 612 1160 638 1212
rect 638 1160 658 1212
rect 658 1160 668 1212
rect 702 1160 710 1212
rect 710 1160 730 1212
rect 730 1160 758 1212
rect 794 1160 802 1212
rect 802 1160 850 1212
rect 1226 1212 1282 1216
rect 1316 1212 1372 1216
rect 1406 1212 1462 1216
rect 1498 1212 1554 1216
rect 1226 1160 1274 1212
rect 1274 1160 1282 1212
rect 1316 1160 1342 1212
rect 1342 1160 1362 1212
rect 1362 1160 1372 1212
rect 1406 1160 1414 1212
rect 1414 1160 1434 1212
rect 1434 1160 1462 1212
rect 1498 1160 1506 1212
rect 1506 1160 1554 1212
rect 522 1066 578 1068
rect 612 1066 668 1068
rect 702 1066 758 1068
rect 794 1066 850 1068
rect 522 1014 570 1066
rect 570 1014 578 1066
rect 612 1014 638 1066
rect 638 1014 658 1066
rect 658 1014 668 1066
rect 702 1014 710 1066
rect 710 1014 730 1066
rect 730 1014 758 1066
rect 794 1014 802 1066
rect 802 1014 850 1066
rect 522 1012 578 1014
rect 612 1012 668 1014
rect 702 1012 758 1014
rect 794 1012 850 1014
rect 458 804 514 860
rect 538 804 594 860
rect 618 804 674 860
rect 698 804 754 860
rect 778 804 834 860
rect 858 804 914 860
rect 458 724 514 780
rect 538 724 594 780
rect 618 724 674 780
rect 698 724 754 780
rect 778 724 834 780
rect 858 724 914 780
rect 458 640 514 696
rect 538 640 594 696
rect 618 640 674 696
rect 698 640 754 696
rect 778 640 834 696
rect 858 640 914 696
rect 1162 804 1218 860
rect 1242 804 1298 860
rect 1322 804 1378 860
rect 1402 804 1458 860
rect 1482 804 1538 860
rect 1562 804 1618 860
rect 1162 724 1218 780
rect 1242 724 1298 780
rect 1322 724 1378 780
rect 1402 724 1458 780
rect 1482 724 1538 780
rect 1562 724 1618 780
rect 1162 640 1218 696
rect 1242 640 1298 696
rect 1322 640 1378 696
rect 1402 640 1458 696
rect 1482 640 1538 696
rect 1562 640 1618 696
rect 378 364 434 420
rect 458 364 514 420
rect 538 364 594 420
rect 618 364 674 420
rect 698 364 754 420
rect 778 364 834 420
rect 858 364 914 420
rect 938 364 994 420
rect 378 284 434 340
rect 458 284 514 340
rect 538 284 594 340
rect 618 284 674 340
rect 698 284 754 340
rect 778 284 834 340
rect 858 284 914 340
rect 938 284 994 340
rect 1082 92 1138 148
rect 1162 92 1218 148
rect 1242 92 1298 148
rect 1322 92 1378 148
rect 1402 92 1458 148
rect 1482 92 1538 148
rect 1562 92 1618 148
rect 1642 92 1698 148
rect 1082 12 1138 68
rect 1162 12 1218 68
rect 1242 12 1298 68
rect 1322 12 1378 68
rect 1402 12 1458 68
rect 1482 12 1538 68
rect 1562 12 1618 68
rect 1642 12 1698 68
rect 544 -112 590 -86
rect 590 -112 600 -86
rect 624 -112 654 -86
rect 654 -112 666 -86
rect 666 -112 680 -86
rect 704 -112 718 -86
rect 718 -112 730 -86
rect 730 -112 760 -86
rect 784 -112 794 -86
rect 794 -112 840 -86
rect 544 -142 600 -112
rect 624 -142 680 -112
rect 704 -142 760 -112
rect 784 -142 840 -112
rect 1248 -112 1294 -86
rect 1294 -112 1304 -86
rect 1328 -112 1358 -86
rect 1358 -112 1370 -86
rect 1370 -112 1384 -86
rect 1408 -112 1422 -86
rect 1422 -112 1434 -86
rect 1434 -112 1464 -86
rect 1488 -112 1498 -86
rect 1498 -112 1544 -86
rect 1248 -142 1304 -112
rect 1328 -142 1384 -112
rect 1408 -142 1464 -112
rect 1488 -142 1544 -112
<< metal3 >>
rect -228 2502 1564 2508
rect -228 2438 -222 2502
rect -158 2438 -142 2502
rect -78 2438 1564 2502
rect -228 2432 -72 2438
rect 32 2372 860 2378
rect 32 2308 38 2372
rect 102 2308 118 2372
rect 182 2370 860 2372
rect 182 2314 544 2370
rect 600 2314 624 2370
rect 680 2314 704 2370
rect 760 2314 784 2370
rect 840 2314 860 2370
rect 182 2308 860 2314
rect 1216 2370 1564 2438
rect 1216 2314 1248 2370
rect 1304 2314 1328 2370
rect 1384 2314 1408 2370
rect 1464 2314 1488 2370
rect 1544 2314 1564 2370
rect 1216 2308 1564 2314
rect 32 2302 188 2308
rect 348 2222 2892 2248
rect 348 2216 2720 2222
rect 348 2160 378 2216
rect 434 2160 458 2216
rect 514 2160 538 2216
rect 594 2160 618 2216
rect 674 2160 698 2216
rect 754 2160 778 2216
rect 834 2160 858 2216
rect 914 2160 938 2216
rect 994 2160 2720 2216
rect 348 2158 2720 2160
rect 2784 2158 2800 2222
rect 2864 2158 2892 2222
rect 348 2136 2892 2158
rect 348 2080 378 2136
rect 434 2080 458 2136
rect 514 2080 538 2136
rect 594 2080 618 2136
rect 674 2080 698 2136
rect 754 2080 778 2136
rect 834 2080 858 2136
rect 914 2080 938 2136
rect 994 2080 2720 2136
rect 348 2072 2720 2080
rect 2784 2072 2800 2136
rect 2864 2072 2892 2136
rect 348 2048 2892 2072
rect 348 1950 2632 1976
rect 348 1944 2460 1950
rect 348 1888 1082 1944
rect 1138 1888 1162 1944
rect 1218 1888 1242 1944
rect 1298 1888 1322 1944
rect 1378 1888 1402 1944
rect 1458 1888 1482 1944
rect 1538 1888 1562 1944
rect 1618 1888 1642 1944
rect 1698 1888 2460 1944
rect 348 1886 2460 1888
rect 2524 1886 2540 1950
rect 2604 1886 2632 1950
rect 348 1864 2632 1886
rect 348 1808 1082 1864
rect 1138 1808 1162 1864
rect 1218 1808 1242 1864
rect 1298 1808 1322 1864
rect 1378 1808 1402 1864
rect 1458 1808 1482 1864
rect 1538 1808 1562 1864
rect 1618 1808 1642 1864
rect 1698 1808 2460 1864
rect 348 1800 2460 1808
rect 2524 1800 2540 1864
rect 2604 1800 2632 1864
rect 348 1776 2632 1800
rect 374 1592 998 1638
rect 374 1528 454 1592
rect 518 1528 534 1592
rect 598 1528 614 1592
rect 678 1528 694 1592
rect 758 1528 774 1592
rect 838 1528 854 1592
rect 918 1528 998 1592
rect 374 1512 998 1528
rect 374 1448 454 1512
rect 518 1448 534 1512
rect 598 1448 614 1512
rect 678 1448 694 1512
rect 758 1448 774 1512
rect 838 1448 854 1512
rect 918 1448 998 1512
rect 374 1428 998 1448
rect 374 1364 454 1428
rect 518 1364 534 1428
rect 598 1364 614 1428
rect 678 1364 694 1428
rect 758 1364 774 1428
rect 838 1364 854 1428
rect 918 1364 998 1428
rect 374 1318 998 1364
rect 1078 1592 1702 1638
rect 1078 1528 1158 1592
rect 1222 1528 1238 1592
rect 1302 1528 1318 1592
rect 1382 1528 1398 1592
rect 1462 1528 1478 1592
rect 1542 1528 1558 1592
rect 1622 1528 1702 1592
rect 1078 1512 1702 1528
rect 1078 1448 1158 1512
rect 1222 1448 1238 1512
rect 1302 1448 1318 1512
rect 1382 1448 1398 1512
rect 1462 1448 1478 1512
rect 1542 1448 1558 1512
rect 1622 1448 1702 1512
rect 1078 1428 1702 1448
rect 1078 1364 1158 1428
rect 1222 1364 1238 1428
rect 1302 1364 1318 1428
rect 1382 1364 1398 1428
rect 1462 1364 1478 1428
rect 1542 1364 1558 1428
rect 1622 1364 1702 1428
rect 1078 1318 1702 1364
rect -98 1224 58 1230
rect -98 1220 -92 1224
rect -356 1160 -92 1220
rect -28 1160 -12 1224
rect 52 1220 58 1224
rect 512 1220 860 1222
rect 1216 1220 1564 1222
rect 52 1216 944 1220
rect 52 1160 522 1216
rect 578 1160 612 1216
rect 668 1160 702 1216
rect 758 1160 794 1216
rect 850 1160 944 1216
rect -356 1154 944 1160
rect 1004 1216 2432 1220
rect 1004 1160 1226 1216
rect 1282 1160 1316 1216
rect 1372 1160 1406 1216
rect 1462 1160 1498 1216
rect 1554 1160 2432 1216
rect 1004 1154 2432 1160
rect 1004 1074 1070 1154
rect -356 1068 2432 1074
rect -356 1008 -308 1068
rect -314 1004 -308 1008
rect -244 1004 -228 1068
rect -164 1008 38 1068
rect -164 1004 -158 1008
rect -314 998 -158 1004
rect 32 1004 38 1008
rect 102 1004 118 1068
rect 182 1012 522 1068
rect 578 1012 612 1068
rect 668 1012 702 1068
rect 758 1012 794 1068
rect 850 1012 2432 1068
rect 182 1008 2432 1012
rect 182 1004 188 1008
rect 512 1006 860 1008
rect 32 998 188 1004
rect 374 864 998 910
rect 374 800 454 864
rect 518 800 534 864
rect 598 800 614 864
rect 678 800 694 864
rect 758 800 774 864
rect 838 800 854 864
rect 918 800 998 864
rect 374 784 998 800
rect 374 720 454 784
rect 518 720 534 784
rect 598 720 614 784
rect 678 720 694 784
rect 758 720 774 784
rect 838 720 854 784
rect 918 720 998 784
rect 374 700 998 720
rect 374 636 454 700
rect 518 636 534 700
rect 598 636 614 700
rect 678 636 694 700
rect 758 636 774 700
rect 838 636 854 700
rect 918 636 998 700
rect 374 590 998 636
rect 1078 864 1702 910
rect 1078 800 1158 864
rect 1222 800 1238 864
rect 1302 800 1318 864
rect 1382 800 1398 864
rect 1462 800 1478 864
rect 1542 800 1558 864
rect 1622 800 1702 864
rect 1078 784 1702 800
rect 1078 720 1158 784
rect 1222 720 1238 784
rect 1302 720 1318 784
rect 1382 720 1398 784
rect 1462 720 1478 784
rect 1542 720 1558 784
rect 1622 720 1702 784
rect 1078 700 1702 720
rect 1078 636 1158 700
rect 1222 636 1238 700
rect 1302 636 1318 700
rect 1382 636 1398 700
rect 1462 636 1478 700
rect 1542 636 1558 700
rect 1622 636 1702 700
rect 1078 590 1702 636
rect 348 430 2632 452
rect 348 420 2458 430
rect 348 364 378 420
rect 434 364 458 420
rect 514 364 538 420
rect 594 364 618 420
rect 674 364 698 420
rect 754 364 778 420
rect 834 364 858 420
rect 914 364 938 420
rect 994 366 2458 420
rect 2522 366 2538 430
rect 2602 366 2632 430
rect 994 364 2632 366
rect 348 344 2632 364
rect 348 340 2458 344
rect 348 284 378 340
rect 434 284 458 340
rect 514 284 538 340
rect 594 284 618 340
rect 674 284 698 340
rect 754 284 778 340
rect 834 284 858 340
rect 914 284 938 340
rect 994 284 2458 340
rect 348 280 2458 284
rect 2522 280 2538 344
rect 2602 280 2632 344
rect 348 252 2632 280
rect 348 158 2892 180
rect 348 148 2718 158
rect 348 92 1082 148
rect 1138 92 1162 148
rect 1218 92 1242 148
rect 1298 92 1322 148
rect 1378 92 1402 148
rect 1458 92 1482 148
rect 1538 92 1562 148
rect 1618 92 1642 148
rect 1698 94 2718 148
rect 2782 94 2798 158
rect 2862 94 2892 158
rect 1698 92 2892 94
rect 348 72 2892 92
rect 348 68 2718 72
rect 348 12 1082 68
rect 1138 12 1162 68
rect 1218 12 1242 68
rect 1298 12 1322 68
rect 1378 12 1402 68
rect 1458 12 1482 68
rect 1538 12 1562 68
rect 1618 12 1642 68
rect 1698 12 2718 68
rect 348 8 2718 12
rect 2782 8 2798 72
rect 2862 8 2892 72
rect 348 -20 2892 8
rect 32 -80 188 -74
rect 32 -144 38 -80
rect 102 -144 118 -80
rect 182 -86 860 -80
rect 182 -142 544 -86
rect 600 -142 624 -86
rect 680 -142 704 -86
rect 760 -142 784 -86
rect 840 -142 860 -86
rect 182 -144 860 -142
rect 32 -150 860 -144
rect 1216 -86 1564 -80
rect 1216 -142 1248 -86
rect 1304 -142 1328 -86
rect 1384 -142 1408 -86
rect 1464 -142 1488 -86
rect 1544 -142 1564 -86
rect 1216 -210 1564 -142
rect -98 -216 1564 -210
rect -98 -280 -92 -216
rect -28 -280 -12 -216
rect 52 -280 1564 -216
rect -98 -286 58 -280
<< via3 >>
rect -222 2438 -158 2502
rect -142 2438 -78 2502
rect 38 2308 102 2372
rect 118 2308 182 2372
rect 2720 2158 2784 2222
rect 2800 2158 2864 2222
rect 2720 2072 2784 2136
rect 2800 2072 2864 2136
rect 2460 1886 2524 1950
rect 2540 1886 2604 1950
rect 2460 1800 2524 1864
rect 2540 1800 2604 1864
rect 454 1588 518 1592
rect 454 1532 458 1588
rect 458 1532 514 1588
rect 514 1532 518 1588
rect 454 1528 518 1532
rect 534 1588 598 1592
rect 534 1532 538 1588
rect 538 1532 594 1588
rect 594 1532 598 1588
rect 534 1528 598 1532
rect 614 1588 678 1592
rect 614 1532 618 1588
rect 618 1532 674 1588
rect 674 1532 678 1588
rect 614 1528 678 1532
rect 694 1588 758 1592
rect 694 1532 698 1588
rect 698 1532 754 1588
rect 754 1532 758 1588
rect 694 1528 758 1532
rect 774 1588 838 1592
rect 774 1532 778 1588
rect 778 1532 834 1588
rect 834 1532 838 1588
rect 774 1528 838 1532
rect 854 1588 918 1592
rect 854 1532 858 1588
rect 858 1532 914 1588
rect 914 1532 918 1588
rect 854 1528 918 1532
rect 454 1508 518 1512
rect 454 1452 458 1508
rect 458 1452 514 1508
rect 514 1452 518 1508
rect 454 1448 518 1452
rect 534 1508 598 1512
rect 534 1452 538 1508
rect 538 1452 594 1508
rect 594 1452 598 1508
rect 534 1448 598 1452
rect 614 1508 678 1512
rect 614 1452 618 1508
rect 618 1452 674 1508
rect 674 1452 678 1508
rect 614 1448 678 1452
rect 694 1508 758 1512
rect 694 1452 698 1508
rect 698 1452 754 1508
rect 754 1452 758 1508
rect 694 1448 758 1452
rect 774 1508 838 1512
rect 774 1452 778 1508
rect 778 1452 834 1508
rect 834 1452 838 1508
rect 774 1448 838 1452
rect 854 1508 918 1512
rect 854 1452 858 1508
rect 858 1452 914 1508
rect 914 1452 918 1508
rect 854 1448 918 1452
rect 454 1424 518 1428
rect 454 1368 458 1424
rect 458 1368 514 1424
rect 514 1368 518 1424
rect 454 1364 518 1368
rect 534 1424 598 1428
rect 534 1368 538 1424
rect 538 1368 594 1424
rect 594 1368 598 1424
rect 534 1364 598 1368
rect 614 1424 678 1428
rect 614 1368 618 1424
rect 618 1368 674 1424
rect 674 1368 678 1424
rect 614 1364 678 1368
rect 694 1424 758 1428
rect 694 1368 698 1424
rect 698 1368 754 1424
rect 754 1368 758 1424
rect 694 1364 758 1368
rect 774 1424 838 1428
rect 774 1368 778 1424
rect 778 1368 834 1424
rect 834 1368 838 1424
rect 774 1364 838 1368
rect 854 1424 918 1428
rect 854 1368 858 1424
rect 858 1368 914 1424
rect 914 1368 918 1424
rect 854 1364 918 1368
rect 1158 1588 1222 1592
rect 1158 1532 1162 1588
rect 1162 1532 1218 1588
rect 1218 1532 1222 1588
rect 1158 1528 1222 1532
rect 1238 1588 1302 1592
rect 1238 1532 1242 1588
rect 1242 1532 1298 1588
rect 1298 1532 1302 1588
rect 1238 1528 1302 1532
rect 1318 1588 1382 1592
rect 1318 1532 1322 1588
rect 1322 1532 1378 1588
rect 1378 1532 1382 1588
rect 1318 1528 1382 1532
rect 1398 1588 1462 1592
rect 1398 1532 1402 1588
rect 1402 1532 1458 1588
rect 1458 1532 1462 1588
rect 1398 1528 1462 1532
rect 1478 1588 1542 1592
rect 1478 1532 1482 1588
rect 1482 1532 1538 1588
rect 1538 1532 1542 1588
rect 1478 1528 1542 1532
rect 1558 1588 1622 1592
rect 1558 1532 1562 1588
rect 1562 1532 1618 1588
rect 1618 1532 1622 1588
rect 1558 1528 1622 1532
rect 1158 1508 1222 1512
rect 1158 1452 1162 1508
rect 1162 1452 1218 1508
rect 1218 1452 1222 1508
rect 1158 1448 1222 1452
rect 1238 1508 1302 1512
rect 1238 1452 1242 1508
rect 1242 1452 1298 1508
rect 1298 1452 1302 1508
rect 1238 1448 1302 1452
rect 1318 1508 1382 1512
rect 1318 1452 1322 1508
rect 1322 1452 1378 1508
rect 1378 1452 1382 1508
rect 1318 1448 1382 1452
rect 1398 1508 1462 1512
rect 1398 1452 1402 1508
rect 1402 1452 1458 1508
rect 1458 1452 1462 1508
rect 1398 1448 1462 1452
rect 1478 1508 1542 1512
rect 1478 1452 1482 1508
rect 1482 1452 1538 1508
rect 1538 1452 1542 1508
rect 1478 1448 1542 1452
rect 1558 1508 1622 1512
rect 1558 1452 1562 1508
rect 1562 1452 1618 1508
rect 1618 1452 1622 1508
rect 1558 1448 1622 1452
rect 1158 1424 1222 1428
rect 1158 1368 1162 1424
rect 1162 1368 1218 1424
rect 1218 1368 1222 1424
rect 1158 1364 1222 1368
rect 1238 1424 1302 1428
rect 1238 1368 1242 1424
rect 1242 1368 1298 1424
rect 1298 1368 1302 1424
rect 1238 1364 1302 1368
rect 1318 1424 1382 1428
rect 1318 1368 1322 1424
rect 1322 1368 1378 1424
rect 1378 1368 1382 1424
rect 1318 1364 1382 1368
rect 1398 1424 1462 1428
rect 1398 1368 1402 1424
rect 1402 1368 1458 1424
rect 1458 1368 1462 1424
rect 1398 1364 1462 1368
rect 1478 1424 1542 1428
rect 1478 1368 1482 1424
rect 1482 1368 1538 1424
rect 1538 1368 1542 1424
rect 1478 1364 1542 1368
rect 1558 1424 1622 1428
rect 1558 1368 1562 1424
rect 1562 1368 1618 1424
rect 1618 1368 1622 1424
rect 1558 1364 1622 1368
rect -92 1160 -28 1224
rect -12 1160 52 1224
rect -308 1004 -244 1068
rect -228 1004 -164 1068
rect 38 1004 102 1068
rect 118 1004 182 1068
rect 454 860 518 864
rect 454 804 458 860
rect 458 804 514 860
rect 514 804 518 860
rect 454 800 518 804
rect 534 860 598 864
rect 534 804 538 860
rect 538 804 594 860
rect 594 804 598 860
rect 534 800 598 804
rect 614 860 678 864
rect 614 804 618 860
rect 618 804 674 860
rect 674 804 678 860
rect 614 800 678 804
rect 694 860 758 864
rect 694 804 698 860
rect 698 804 754 860
rect 754 804 758 860
rect 694 800 758 804
rect 774 860 838 864
rect 774 804 778 860
rect 778 804 834 860
rect 834 804 838 860
rect 774 800 838 804
rect 854 860 918 864
rect 854 804 858 860
rect 858 804 914 860
rect 914 804 918 860
rect 854 800 918 804
rect 454 780 518 784
rect 454 724 458 780
rect 458 724 514 780
rect 514 724 518 780
rect 454 720 518 724
rect 534 780 598 784
rect 534 724 538 780
rect 538 724 594 780
rect 594 724 598 780
rect 534 720 598 724
rect 614 780 678 784
rect 614 724 618 780
rect 618 724 674 780
rect 674 724 678 780
rect 614 720 678 724
rect 694 780 758 784
rect 694 724 698 780
rect 698 724 754 780
rect 754 724 758 780
rect 694 720 758 724
rect 774 780 838 784
rect 774 724 778 780
rect 778 724 834 780
rect 834 724 838 780
rect 774 720 838 724
rect 854 780 918 784
rect 854 724 858 780
rect 858 724 914 780
rect 914 724 918 780
rect 854 720 918 724
rect 454 696 518 700
rect 454 640 458 696
rect 458 640 514 696
rect 514 640 518 696
rect 454 636 518 640
rect 534 696 598 700
rect 534 640 538 696
rect 538 640 594 696
rect 594 640 598 696
rect 534 636 598 640
rect 614 696 678 700
rect 614 640 618 696
rect 618 640 674 696
rect 674 640 678 696
rect 614 636 678 640
rect 694 696 758 700
rect 694 640 698 696
rect 698 640 754 696
rect 754 640 758 696
rect 694 636 758 640
rect 774 696 838 700
rect 774 640 778 696
rect 778 640 834 696
rect 834 640 838 696
rect 774 636 838 640
rect 854 696 918 700
rect 854 640 858 696
rect 858 640 914 696
rect 914 640 918 696
rect 854 636 918 640
rect 1158 860 1222 864
rect 1158 804 1162 860
rect 1162 804 1218 860
rect 1218 804 1222 860
rect 1158 800 1222 804
rect 1238 860 1302 864
rect 1238 804 1242 860
rect 1242 804 1298 860
rect 1298 804 1302 860
rect 1238 800 1302 804
rect 1318 860 1382 864
rect 1318 804 1322 860
rect 1322 804 1378 860
rect 1378 804 1382 860
rect 1318 800 1382 804
rect 1398 860 1462 864
rect 1398 804 1402 860
rect 1402 804 1458 860
rect 1458 804 1462 860
rect 1398 800 1462 804
rect 1478 860 1542 864
rect 1478 804 1482 860
rect 1482 804 1538 860
rect 1538 804 1542 860
rect 1478 800 1542 804
rect 1558 860 1622 864
rect 1558 804 1562 860
rect 1562 804 1618 860
rect 1618 804 1622 860
rect 1558 800 1622 804
rect 1158 780 1222 784
rect 1158 724 1162 780
rect 1162 724 1218 780
rect 1218 724 1222 780
rect 1158 720 1222 724
rect 1238 780 1302 784
rect 1238 724 1242 780
rect 1242 724 1298 780
rect 1298 724 1302 780
rect 1238 720 1302 724
rect 1318 780 1382 784
rect 1318 724 1322 780
rect 1322 724 1378 780
rect 1378 724 1382 780
rect 1318 720 1382 724
rect 1398 780 1462 784
rect 1398 724 1402 780
rect 1402 724 1458 780
rect 1458 724 1462 780
rect 1398 720 1462 724
rect 1478 780 1542 784
rect 1478 724 1482 780
rect 1482 724 1538 780
rect 1538 724 1542 780
rect 1478 720 1542 724
rect 1558 780 1622 784
rect 1558 724 1562 780
rect 1562 724 1618 780
rect 1618 724 1622 780
rect 1558 720 1622 724
rect 1158 696 1222 700
rect 1158 640 1162 696
rect 1162 640 1218 696
rect 1218 640 1222 696
rect 1158 636 1222 640
rect 1238 696 1302 700
rect 1238 640 1242 696
rect 1242 640 1298 696
rect 1298 640 1302 696
rect 1238 636 1302 640
rect 1318 696 1382 700
rect 1318 640 1322 696
rect 1322 640 1378 696
rect 1378 640 1382 696
rect 1318 636 1382 640
rect 1398 696 1462 700
rect 1398 640 1402 696
rect 1402 640 1458 696
rect 1458 640 1462 696
rect 1398 636 1462 640
rect 1478 696 1542 700
rect 1478 640 1482 696
rect 1482 640 1538 696
rect 1538 640 1542 696
rect 1478 636 1542 640
rect 1558 696 1622 700
rect 1558 640 1562 696
rect 1562 640 1618 696
rect 1618 640 1622 696
rect 1558 636 1622 640
rect 2458 366 2522 430
rect 2538 366 2602 430
rect 2458 280 2522 344
rect 2538 280 2602 344
rect 2718 94 2782 158
rect 2798 94 2862 158
rect 2718 8 2782 72
rect 2798 8 2862 72
rect 38 -144 102 -80
rect 118 -144 182 -80
rect -92 -280 -28 -216
rect -12 -280 52 -216
<< metal4 >>
rect -228 2502 -72 2508
rect -228 2438 -222 2502
rect -158 2438 -142 2502
rect -78 2438 -72 2502
rect -228 2432 -72 2438
rect -228 1074 -158 2432
rect 32 2372 188 2378
rect 32 2308 38 2372
rect 102 2308 118 2372
rect 182 2308 188 2372
rect 32 2302 188 2308
rect 32 1230 102 2302
rect 2692 2222 2892 2248
rect 2692 2158 2720 2222
rect 2784 2158 2800 2222
rect 2864 2158 2892 2222
rect 2692 2136 2892 2158
rect 2692 2072 2720 2136
rect 2784 2072 2800 2136
rect 2864 2072 2892 2136
rect 2432 1950 2632 1976
rect 2432 1886 2460 1950
rect 2524 1886 2540 1950
rect 2604 1886 2632 1950
rect 2432 1864 2632 1886
rect 2432 1800 2460 1864
rect 2524 1800 2540 1864
rect 2604 1800 2632 1864
rect 374 1596 998 1638
rect 374 1360 408 1596
rect 644 1592 728 1596
rect 678 1528 694 1592
rect 644 1512 728 1528
rect 678 1448 694 1512
rect 644 1428 728 1448
rect 678 1364 694 1428
rect 644 1360 728 1364
rect 964 1360 998 1596
rect 374 1318 998 1360
rect 1078 1596 1702 1638
rect 1078 1360 1112 1596
rect 1348 1592 1432 1596
rect 1382 1528 1398 1592
rect 1348 1512 1432 1528
rect 1382 1448 1398 1512
rect 1348 1428 1432 1448
rect 1382 1364 1398 1428
rect 1348 1360 1432 1364
rect 1668 1360 1702 1596
rect 1078 1318 1702 1360
rect -314 1068 -158 1074
rect -314 1004 -308 1068
rect -244 1004 -228 1068
rect -164 1004 -158 1068
rect -314 998 -158 1004
rect -98 1224 102 1230
rect -98 1160 -92 1224
rect -28 1160 -12 1224
rect 52 1160 102 1224
rect -98 1154 102 1160
rect -98 -210 -28 1154
rect 32 1068 188 1074
rect 32 1004 38 1068
rect 102 1004 118 1068
rect 182 1004 188 1068
rect 32 998 188 1004
rect 32 -74 102 998
rect 374 868 998 910
rect 374 632 408 868
rect 644 864 728 868
rect 678 800 694 864
rect 644 784 728 800
rect 678 720 694 784
rect 644 700 728 720
rect 678 636 694 700
rect 644 632 728 636
rect 964 632 998 868
rect 374 590 998 632
rect 1078 868 1702 910
rect 1078 632 1112 868
rect 1348 864 1432 868
rect 1382 800 1398 864
rect 1348 784 1432 800
rect 1382 720 1398 784
rect 1348 700 1432 720
rect 1382 636 1398 700
rect 1348 632 1432 636
rect 1668 632 1702 868
rect 1078 590 1702 632
rect 1894 590 2294 910
rect 2432 430 2632 1800
rect 2432 366 2458 430
rect 2522 366 2538 430
rect 2602 366 2632 430
rect 2432 344 2632 366
rect 2432 280 2458 344
rect 2522 280 2538 344
rect 2602 280 2632 344
rect 2432 252 2632 280
rect 2692 158 2892 2072
rect 2952 1596 3286 1638
rect 2952 1360 3000 1596
rect 3236 1360 3286 1596
rect 2952 868 3286 1360
rect 2952 632 3000 868
rect 3236 632 3286 868
rect 2952 590 3286 632
rect 2692 94 2718 158
rect 2782 94 2798 158
rect 2862 94 2892 158
rect 2692 72 2892 94
rect 2692 8 2718 72
rect 2782 8 2798 72
rect 2862 8 2892 72
rect 2692 -20 2892 8
rect 32 -80 188 -74
rect 32 -144 38 -80
rect 102 -144 118 -80
rect 182 -144 188 -80
rect 32 -150 188 -144
rect -98 -216 58 -210
rect -98 -280 -92 -216
rect -28 -280 -12 -216
rect 52 -280 58 -216
rect -98 -286 58 -280
<< via4 >>
rect 408 1592 644 1596
rect 728 1592 964 1596
rect 408 1528 454 1592
rect 454 1528 518 1592
rect 518 1528 534 1592
rect 534 1528 598 1592
rect 598 1528 614 1592
rect 614 1528 644 1592
rect 728 1528 758 1592
rect 758 1528 774 1592
rect 774 1528 838 1592
rect 838 1528 854 1592
rect 854 1528 918 1592
rect 918 1528 964 1592
rect 408 1512 644 1528
rect 728 1512 964 1528
rect 408 1448 454 1512
rect 454 1448 518 1512
rect 518 1448 534 1512
rect 534 1448 598 1512
rect 598 1448 614 1512
rect 614 1448 644 1512
rect 728 1448 758 1512
rect 758 1448 774 1512
rect 774 1448 838 1512
rect 838 1448 854 1512
rect 854 1448 918 1512
rect 918 1448 964 1512
rect 408 1428 644 1448
rect 728 1428 964 1448
rect 408 1364 454 1428
rect 454 1364 518 1428
rect 518 1364 534 1428
rect 534 1364 598 1428
rect 598 1364 614 1428
rect 614 1364 644 1428
rect 728 1364 758 1428
rect 758 1364 774 1428
rect 774 1364 838 1428
rect 838 1364 854 1428
rect 854 1364 918 1428
rect 918 1364 964 1428
rect 408 1360 644 1364
rect 728 1360 964 1364
rect 1112 1592 1348 1596
rect 1432 1592 1668 1596
rect 1112 1528 1158 1592
rect 1158 1528 1222 1592
rect 1222 1528 1238 1592
rect 1238 1528 1302 1592
rect 1302 1528 1318 1592
rect 1318 1528 1348 1592
rect 1432 1528 1462 1592
rect 1462 1528 1478 1592
rect 1478 1528 1542 1592
rect 1542 1528 1558 1592
rect 1558 1528 1622 1592
rect 1622 1528 1668 1592
rect 1112 1512 1348 1528
rect 1432 1512 1668 1528
rect 1112 1448 1158 1512
rect 1158 1448 1222 1512
rect 1222 1448 1238 1512
rect 1238 1448 1302 1512
rect 1302 1448 1318 1512
rect 1318 1448 1348 1512
rect 1432 1448 1462 1512
rect 1462 1448 1478 1512
rect 1478 1448 1542 1512
rect 1542 1448 1558 1512
rect 1558 1448 1622 1512
rect 1622 1448 1668 1512
rect 1112 1428 1348 1448
rect 1432 1428 1668 1448
rect 1112 1364 1158 1428
rect 1158 1364 1222 1428
rect 1222 1364 1238 1428
rect 1238 1364 1302 1428
rect 1302 1364 1318 1428
rect 1318 1364 1348 1428
rect 1432 1364 1462 1428
rect 1462 1364 1478 1428
rect 1478 1364 1542 1428
rect 1542 1364 1558 1428
rect 1558 1364 1622 1428
rect 1622 1364 1668 1428
rect 1112 1360 1348 1364
rect 1432 1360 1668 1364
rect 408 864 644 868
rect 728 864 964 868
rect 408 800 454 864
rect 454 800 518 864
rect 518 800 534 864
rect 534 800 598 864
rect 598 800 614 864
rect 614 800 644 864
rect 728 800 758 864
rect 758 800 774 864
rect 774 800 838 864
rect 838 800 854 864
rect 854 800 918 864
rect 918 800 964 864
rect 408 784 644 800
rect 728 784 964 800
rect 408 720 454 784
rect 454 720 518 784
rect 518 720 534 784
rect 534 720 598 784
rect 598 720 614 784
rect 614 720 644 784
rect 728 720 758 784
rect 758 720 774 784
rect 774 720 838 784
rect 838 720 854 784
rect 854 720 918 784
rect 918 720 964 784
rect 408 700 644 720
rect 728 700 964 720
rect 408 636 454 700
rect 454 636 518 700
rect 518 636 534 700
rect 534 636 598 700
rect 598 636 614 700
rect 614 636 644 700
rect 728 636 758 700
rect 758 636 774 700
rect 774 636 838 700
rect 838 636 854 700
rect 854 636 918 700
rect 918 636 964 700
rect 408 632 644 636
rect 728 632 964 636
rect 1112 864 1348 868
rect 1432 864 1668 868
rect 1112 800 1158 864
rect 1158 800 1222 864
rect 1222 800 1238 864
rect 1238 800 1302 864
rect 1302 800 1318 864
rect 1318 800 1348 864
rect 1432 800 1462 864
rect 1462 800 1478 864
rect 1478 800 1542 864
rect 1542 800 1558 864
rect 1558 800 1622 864
rect 1622 800 1668 864
rect 1112 784 1348 800
rect 1432 784 1668 800
rect 1112 720 1158 784
rect 1158 720 1222 784
rect 1222 720 1238 784
rect 1238 720 1302 784
rect 1302 720 1318 784
rect 1318 720 1348 784
rect 1432 720 1462 784
rect 1462 720 1478 784
rect 1478 720 1542 784
rect 1542 720 1558 784
rect 1558 720 1622 784
rect 1622 720 1668 784
rect 1112 700 1348 720
rect 1432 700 1668 720
rect 1112 636 1158 700
rect 1158 636 1222 700
rect 1222 636 1238 700
rect 1238 636 1302 700
rect 1302 636 1318 700
rect 1318 636 1348 700
rect 1432 636 1462 700
rect 1462 636 1478 700
rect 1478 636 1542 700
rect 1542 636 1558 700
rect 1558 636 1622 700
rect 1622 636 1668 700
rect 1112 632 1348 636
rect 1432 632 1668 636
rect 3000 1360 3236 1596
rect 3000 632 3236 868
<< metal5 >>
rect 374 1596 3286 1638
rect 374 1360 408 1596
rect 644 1360 728 1596
rect 964 1360 1112 1596
rect 1348 1360 1432 1596
rect 1668 1360 3000 1596
rect 3236 1360 3286 1596
rect 374 1318 3286 1360
rect 348 868 3286 910
rect 348 632 408 868
rect 644 632 728 868
rect 964 632 1112 868
rect 1348 632 1432 868
rect 1668 632 3000 868
rect 3236 632 3286 868
rect 348 590 3286 632
use buffer_input_base  buffer_input_base_0
timestamp 1654464469
transform 1 0 -218 0 1 -100
box -138 -20 2650 2448
<< labels >>
flabel metal1 s -57 2299 25 2324 0 FreeSans 300 0 0 0 GATE
port 2 nsew
<< end >>
