magic
tech sky130B
timestamp 1654424727
<< metal1 >>
rect -1940 49375 -940 55395
rect -1940 26195 -935 29655
rect 36780 28135 38800 29135
rect -1940 25195 20 26195
rect -1940 24675 -935 25195
rect 37800 24195 38800 28135
rect 36780 23195 38800 24195
rect -1940 16315 -935 19775
rect 36780 18255 38800 19255
rect -1940 15315 20 16315
rect -1940 11375 -935 15315
rect 37800 14315 38800 18255
rect 36780 13315 38800 14315
rect -1940 10375 20 11375
rect -1940 6435 -935 10375
rect 37800 9375 38800 13315
rect 36780 8375 38800 9375
rect -1940 5435 20 6435
rect -1940 4915 -935 5435
rect 37800 4435 38800 8375
rect 36780 3435 38800 4435
<< metal2 >>
rect -3440 49375 -2440 55395
rect 4580 46205 41300 47205
rect 9180 41265 41300 42265
rect 18380 36325 41300 37325
rect 36780 31385 41300 32385
rect -3440 24675 -2435 29655
rect 36780 26445 40800 27445
rect 39800 22505 40800 26445
rect 36780 21505 41300 22505
rect -3440 4915 -2435 19775
rect 36780 16565 40800 17565
rect 39800 12625 40800 16565
rect 36780 11625 40800 12625
rect 39800 7685 40800 11625
rect 36780 6685 40800 7685
rect 39800 2745 40800 6685
rect 36780 1745 41300 2745
<< metal3 >>
rect -3437 54895 35363 54898
rect -4880 53905 3110 54895
rect 4100 53905 7710 54895
rect 8700 53905 12310 54895
rect 13300 53905 16910 54895
rect 17900 53905 21510 54895
rect 22500 53905 26110 54895
rect 27100 54890 35363 54895
rect 36305 54890 41300 54900
rect 27100 53905 30710 54890
rect -4880 53900 30710 53905
rect 31700 53900 35310 54890
rect 36300 53900 41300 54890
rect -4880 53895 36305 53900
rect -4880 51890 35360 51895
rect 36305 51890 41300 51895
rect -4880 50900 505 51890
rect 1495 50900 5105 51890
rect 6095 50900 9705 51890
rect 10695 50900 14305 51890
rect 15295 50900 18905 51890
rect 19895 50900 23505 51890
rect 24495 50900 28105 51890
rect 29095 50900 32705 51890
rect 33695 50900 41300 51890
rect -4880 50895 41300 50900
<< via3 >>
rect 3110 53905 4100 54895
rect 7710 53905 8700 54895
rect 12310 53905 13300 54895
rect 16910 53905 17900 54895
rect 21510 53905 22500 54895
rect 26110 53905 27100 54895
rect 30710 53900 31700 54890
rect 35310 53900 36300 54890
rect 505 50900 1495 51890
rect 5105 50900 6095 51890
rect 9705 50900 10695 51890
rect 14305 50900 15295 51890
rect 18905 50900 19895 51890
rect 23505 50900 24495 51890
rect 28105 50900 29095 51890
rect 32705 50900 33695 51890
<< metal4 >>
rect 500 51890 1500 55395
rect 500 50900 505 51890
rect 1495 50900 1500 51890
rect 500 49375 1500 50900
rect 3105 54895 4105 55395
rect 3105 53905 3110 54895
rect 4100 53905 4105 54895
rect 3105 49375 4105 53905
rect 5100 51890 6100 55395
rect 5100 50900 5105 51890
rect 6095 50900 6100 51890
rect 5100 44435 6100 50900
rect 7705 54895 8705 55395
rect 7705 53905 7710 54895
rect 8700 53905 8705 54895
rect 7705 44435 8705 53905
rect 9700 51890 10700 55395
rect 9700 50900 9705 51890
rect 10695 50900 10700 51890
rect 9700 39495 10700 50900
rect 12305 54895 13305 55395
rect 12305 53905 12310 54895
rect 13300 53905 13305 54895
rect 12305 39495 13305 53905
rect 14300 51890 15300 55395
rect 14300 50900 14305 51890
rect 15295 50900 15300 51890
rect 14300 39495 15300 50900
rect 16905 54895 17905 55395
rect 16905 53905 16910 54895
rect 17900 53905 17905 54895
rect 16905 39495 17905 53905
rect 18900 51890 19900 55395
rect 18900 50900 18905 51890
rect 19895 50900 19900 51890
rect 18900 34555 19900 50900
rect 21505 54895 22505 55395
rect 21505 53905 21510 54895
rect 22500 53905 22505 54895
rect 21505 34555 22505 53905
rect 23500 51890 24500 55395
rect 23500 50900 23505 51890
rect 24495 50900 24500 51890
rect 23500 34555 24500 50900
rect 26105 54895 27105 55395
rect 26105 53905 26110 54895
rect 27100 53905 27105 54895
rect 26105 34555 27105 53905
rect 28100 51890 29100 55395
rect 28100 50900 28105 51890
rect 29095 50900 29100 51890
rect 28100 34555 29100 50900
rect 30705 54890 31705 55395
rect 30705 53900 30710 54890
rect 31700 53900 31705 54890
rect 30705 34555 31705 53900
rect 32700 51890 33700 55395
rect 32700 50900 32705 51890
rect 33695 50900 33700 51890
rect 32700 34555 33700 50900
rect 35305 54890 36305 55395
rect 35305 53900 35310 54890
rect 36300 53900 36305 54890
rect 35305 34555 36305 53900
use cell_unit  cell_unit_0
timestamp 1654419664
transform 1 0 2110 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_1
timestamp 1654419664
transform 1 0 6710 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_2
timestamp 1654419664
transform 1 0 11310 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_3
timestamp 1654419664
transform 1 0 15910 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_4
timestamp 1654419664
transform 1 0 20510 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_5
timestamp 1654419664
transform 1 0 25110 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_6
timestamp 1654419664
transform 1 0 29710 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_7
timestamp 1654419664
transform 1 0 34310 0 1 2975
box -2110 -2980 2490 1960
use cell_unit  cell_unit_8
timestamp 1654419664
transform 1 0 2110 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_9
timestamp 1654419664
transform 1 0 2110 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_10
timestamp 1654419664
transform 1 0 2110 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_11
timestamp 1654419664
transform 1 0 6710 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_12
timestamp 1654419664
transform 1 0 11310 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_13
timestamp 1654419664
transform 1 0 15910 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_14
timestamp 1654419664
transform 1 0 20510 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_15
timestamp 1654419664
transform 1 0 25110 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_16
timestamp 1654419664
transform 1 0 29710 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_17
timestamp 1654419664
transform 1 0 34310 0 1 7915
box -2110 -2980 2490 1960
use cell_unit  cell_unit_18
timestamp 1654419664
transform 1 0 6710 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_19
timestamp 1654419664
transform 1 0 11310 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_20
timestamp 1654419664
transform 1 0 15910 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_21
timestamp 1654419664
transform 1 0 20510 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_22
timestamp 1654419664
transform 1 0 25110 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_23
timestamp 1654419664
transform 1 0 29710 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_24
timestamp 1654419664
transform 1 0 34310 0 1 12855
box -2110 -2980 2490 1960
use cell_unit  cell_unit_25
timestamp 1654419664
transform 1 0 6710 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_26
timestamp 1654419664
transform 1 0 11310 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_27
timestamp 1654419664
transform 1 0 15910 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_28
timestamp 1654419664
transform 1 0 20510 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_29
timestamp 1654419664
transform 1 0 25110 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_30
timestamp 1654419664
transform 1 0 29710 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_31
timestamp 1654419664
transform 1 0 34310 0 1 17795
box -2110 -2980 2490 1960
use cell_unit  cell_unit_32
timestamp 1654419664
transform 1 0 2110 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_33
timestamp 1654419664
transform 1 0 2110 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_34
timestamp 1654419664
transform 1 0 6710 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_35
timestamp 1654419664
transform 1 0 11310 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_36
timestamp 1654419664
transform 1 0 15910 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_37
timestamp 1654419664
transform 1 0 20510 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_38
timestamp 1654419664
transform 1 0 25110 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_39
timestamp 1654419664
transform 1 0 29710 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_40
timestamp 1654419664
transform 1 0 34310 0 1 22735
box -2110 -2980 2490 1960
use cell_unit  cell_unit_41
timestamp 1654419664
transform 1 0 6710 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_42
timestamp 1654419664
transform 1 0 11310 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_43
timestamp 1654419664
transform 1 0 15910 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_44
timestamp 1654419664
transform 1 0 20510 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_45
timestamp 1654419664
transform 1 0 25110 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_46
timestamp 1654419664
transform 1 0 29710 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_47
timestamp 1654419664
transform 1 0 34310 0 1 27675
box -2110 -2980 2490 1960
use cell_unit  cell_unit_48
timestamp 1654419664
transform 1 0 2110 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_49
timestamp 1654419664
transform 1 0 6710 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_50
timestamp 1654419664
transform 1 0 11310 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_51
timestamp 1654419664
transform 1 0 15910 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_52
timestamp 1654419664
transform 1 0 20510 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_53
timestamp 1654419664
transform 1 0 25110 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_54
timestamp 1654419664
transform 1 0 29710 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_55
timestamp 1654419664
transform 1 0 34310 0 1 32615
box -2110 -2980 2490 1960
use cell_unit  cell_unit_56
timestamp 1654419664
transform 1 0 2110 0 1 37555
box -2110 -2980 2490 1960
use cell_unit  cell_unit_57
timestamp 1654419664
transform 1 0 6710 0 1 37555
box -2110 -2980 2490 1960
use cell_unit  cell_unit_58
timestamp 1654419664
transform 1 0 11310 0 1 37555
box -2110 -2980 2490 1960
use cell_unit  cell_unit_59
timestamp 1654419664
transform 1 0 15910 0 1 37555
box -2110 -2980 2490 1960
use cell_unit  cell_unit_60
timestamp 1654419664
transform 1 0 2110 0 1 42495
box -2110 -2980 2490 1960
use cell_unit  cell_unit_61
timestamp 1654419664
transform 1 0 6710 0 1 42495
box -2110 -2980 2490 1960
use cell_unit  cell_unit_62
timestamp 1654419664
transform 1 0 2110 0 1 47435
box -2110 -2980 2490 1960
use inv_1  inv_1_0
timestamp 1654380766
transform 1 0 -230 0 1 55
box -3210 -60 230 4880
use inv_1  inv_1_1
timestamp 1654380766
transform 1 0 -230 0 1 19815
box -3210 -60 230 4880
use inv_1  inv_1_2
timestamp 1654380766
transform 1 0 -230 0 1 29695
box -3210 -60 230 4880
use inv_1  inv_1_3
timestamp 1654380766
transform 1 0 -230 0 1 34635
box -3210 -60 230 4880
use inv_1  inv_1_4
timestamp 1654380766
transform 1 0 -230 0 1 39575
box -3210 -60 230 4880
use inv_1  inv_1_5
timestamp 1654380766
transform 1 0 -230 0 1 44515
box -3210 -60 230 4880
<< labels >>
flabel metal3 -4880 51360 -4880 51360 3 FreeSans 1200 0 0 0 OUT_P
port 1 e
flabel metal3 41300 54400 41300 54400 7 FreeSans 1200 0 0 0 OUT_N
port 2 w
flabel metal2 41300 46730 41300 46730 7 FreeSans 1200 0 0 0 bit0
port 3 w
flabel metal2 41300 41750 41300 41750 7 FreeSans 1200 0 0 0 bit1
port 4 w
flabel metal2 41300 36795 41300 36795 7 FreeSans 1200 0 0 0 bit2
port 5 w
flabel metal2 41300 31875 41300 31875 7 FreeSans 1200 0 0 0 bit3
port 6 w
flabel metal2 41300 21965 41300 21965 7 FreeSans 1200 0 0 0 bit4
port 7 w
flabel metal2 41300 2195 41300 2195 7 FreeSans 1200 0 0 0 bit5
port 8 w
flabel metal2 -2990 55395 -2990 55395 5 FreeSans 1200 0 0 0 VDD
port 9 s
flabel metal1 -1445 55395 -1445 55395 5 FreeSans 1200 0 0 0 GND
port 10 s
<< end >>
