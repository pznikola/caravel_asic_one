* NGSPICE file created from vco_pair_pex.ext - technology: sky130B

.subckt vco_pair_pex OUT_P OUT_N GND
X0 OUT_N.t13 OUT_P.t14 GND.t77 GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X1 OUT_N.t12 OUT_P.t15 GND.t75 GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X2 GND.t73 OUT_P.t16 OUT_N.t11 GND.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X3 GND GND.t39 GND GND.t40 sky130_fd_pr__nfet_01v8 ad=5.656e+13p pd=4.264e+08u as=0p ps=0u w=5.05e+06u l=150000u
X4 GND.t71 OUT_P.t17 OUT_N.t10 GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X5 GND.t69 OUT_P.t18 OUT_N.t9 GND.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X6 OUT_P.t6 OUT_N.t14 GND.t49 GND.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X7 GND GND.t34 GND GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X8 OUT_N.t8 OUT_P.t19 GND.t67 GND.t66 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X9 GND GND.t29 GND GND.t30 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X10 GND.t91 OUT_N.t15 OUT_P.t13 GND.t90 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X11 OUT_N.t7 OUT_P.t20 GND.t65 GND.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X12 GND.t83 OUT_N.t16 OUT_P.t9 GND.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X13 GND.t28 GND.t25 GND.t27 GND.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X14 GND.t81 OUT_N.t17 OUT_P.t8 GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X15 GND.t63 OUT_P.t21 OUT_N.t6 GND.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X16 OUT_P.t7 OUT_N.t18 GND.t79 GND.t78 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X17 OUT_N.t5 OUT_P.t22 GND.t61 GND.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X18 GND.t87 OUT_N.t19 OUT_P.t11 GND.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X19 GND.t7 OUT_N.t20 OUT_P.t3 GND.t6 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X20 GND.t24 GND.t21 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X21 OUT_P.t10 OUT_N.t21 GND.t85 GND.t84 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X22 GND.t47 OUT_N.t22 OUT_P.t5 GND.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X23 OUT_P.t4 OUT_N.t23 GND.t45 GND.t44 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X24 OUT_P.t1 OUT_N.t24 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X25 OUT_P.t2 OUT_N.t25 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X26 OUT_N.t4 OUT_P.t23 GND.t59 GND.t58 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X27 OUT_P.t0 OUT_N.t26 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X28 GND.t57 OUT_P.t24 OUT_N.t3 GND.t56 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X29 GND.t89 OUT_N.t27 OUT_P.t12 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X30 GND.t55 OUT_P.t25 OUT_N.t2 GND.t54 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X31 GND.t20 GND.t17 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X32 GND.t16 GND.t13 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X33 GND.t53 OUT_P.t26 OUT_N.t1 GND.t52 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X34 GND GND.t8 GND GND.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
X35 OUT_N.t0 OUT_P.t27 GND.t51 GND.t50 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.05e+06u l=150000u
R0 OUT_P.n1266 OUT_P.t24 846.712
R1 OUT_P.n1269 OUT_P.t14 846.712
R2 OUT_P.n1195 OUT_P.t20 846.712
R3 OUT_P.n1209 OUT_P.t26 846.712
R4 OUT_P.n1294 OUT_P.t25 846.712
R5 OUT_P.n1297 OUT_P.t23 846.712
R6 OUT_P.n1158 OUT_P.t15 846.712
R7 OUT_P.n1172 OUT_P.t18 846.712
R8 OUT_P.n1246 OUT_P.t17 846.712
R9 OUT_P.n1233 OUT_P.t22 846.712
R10 OUT_P.n1128 OUT_P.t19 846.712
R11 OUT_P.n1125 OUT_P.t21 846.712
R12 OUT_P.n0 OUT_P.t27 846.712
R13 OUT_P.n1323 OUT_P.t16 846.712
R14 OUT_P.n1267 OUT_P.n1266 24.127
R15 OUT_P.n1270 OUT_P.n1269 24.127
R16 OUT_P.n457 OUT_P.n456 24.127
R17 OUT_P.n440 OUT_P.n439 24.127
R18 OUT_P.n1210 OUT_P.n1209 24.127
R19 OUT_P.n1196 OUT_P.n1195 24.127
R20 OUT_P.n487 OUT_P.n486 24.127
R21 OUT_P.n498 OUT_P.n497 24.127
R22 OUT_P.n1295 OUT_P.n1294 24.127
R23 OUT_P.n1298 OUT_P.n1297 24.127
R24 OUT_P.n538 OUT_P.n537 24.127
R25 OUT_P.n521 OUT_P.n520 24.127
R26 OUT_P.n1173 OUT_P.n1172 24.127
R27 OUT_P.n1159 OUT_P.n1158 24.127
R28 OUT_P.n568 OUT_P.n567 24.127
R29 OUT_P.n580 OUT_P.n579 24.127
R30 OUT_P.n773 OUT_P.n772 24.127
R31 OUT_P.n780 OUT_P.n779 24.127
R32 OUT_P.n1247 OUT_P.n1246 24.127
R33 OUT_P.n1234 OUT_P.n1233 24.127
R34 OUT_P.n1126 OUT_P.n1125 24.127
R35 OUT_P.n1129 OUT_P.n1128 24.127
R36 OUT_P.n614 OUT_P.n613 24.127
R37 OUT_P.n626 OUT_P.n625 24.127
R38 OUT_P.n667 OUT_P.n666 24.127
R39 OUT_P.n675 OUT_P.n674 24.127
R40 OUT_P.n1324 OUT_P.n1323 24.127
R41 OUT_P.n1 OUT_P.n0 24.127
R42 OUT_P.n874 OUT_P.n873 9.31
R43 OUT_P.n975 OUT_P.n974 9.31
R44 OUT_P.n1076 OUT_P.n1075 9.31
R45 OUT_P.n42 OUT_P.n41 9.3
R46 OUT_P.n40 OUT_P.n39 9.3
R47 OUT_P.n52 OUT_P.n51 9.3
R48 OUT_P.n82 OUT_P.n81 9.3
R49 OUT_P.n72 OUT_P.n71 9.3
R50 OUT_P.n80 OUT_P.n79 9.3
R51 OUT_P.n77 OUT_P.n76 9.3
R52 OUT_P.n70 OUT_P.n69 9.3
R53 OUT_P.n66 OUT_P.n65 9.3
R54 OUT_P.n60 OUT_P.n59 9.3
R55 OUT_P.n56 OUT_P.n55 9.3
R56 OUT_P.n20 OUT_P.n19 9.3
R57 OUT_P.n47 OUT_P.n46 9.3
R58 OUT_P.n87 OUT_P.n86 9.3
R59 OUT_P.n209 OUT_P.n208 9.3
R60 OUT_P.n198 OUT_P.n197 9.3
R61 OUT_P.n204 OUT_P.n203 9.3
R62 OUT_P.n162 OUT_P.n161 9.3
R63 OUT_P.n164 OUT_P.n163 9.3
R64 OUT_P.n202 OUT_P.n201 9.3
R65 OUT_P.n182 OUT_P.n181 9.3
R66 OUT_P.n178 OUT_P.n177 9.3
R67 OUT_P.n174 OUT_P.n173 9.3
R68 OUT_P.n170 OUT_P.n169 9.3
R69 OUT_P.n188 OUT_P.n187 9.3
R70 OUT_P.n191 OUT_P.n190 9.3
R71 OUT_P.n193 OUT_P.n192 9.3
R72 OUT_P.n125 OUT_P.n124 9.3
R73 OUT_P.n314 OUT_P.n313 9.3
R74 OUT_P.n303 OUT_P.n302 9.3
R75 OUT_P.n309 OUT_P.n308 9.3
R76 OUT_P.n267 OUT_P.n266 9.3
R77 OUT_P.n269 OUT_P.n268 9.3
R78 OUT_P.n307 OUT_P.n306 9.3
R79 OUT_P.n287 OUT_P.n286 9.3
R80 OUT_P.n283 OUT_P.n282 9.3
R81 OUT_P.n279 OUT_P.n278 9.3
R82 OUT_P.n275 OUT_P.n274 9.3
R83 OUT_P.n293 OUT_P.n292 9.3
R84 OUT_P.n296 OUT_P.n295 9.3
R85 OUT_P.n298 OUT_P.n297 9.3
R86 OUT_P.n230 OUT_P.n229 9.3
R87 OUT_P.n419 OUT_P.n418 9.3
R88 OUT_P.n408 OUT_P.n407 9.3
R89 OUT_P.n414 OUT_P.n413 9.3
R90 OUT_P.n372 OUT_P.n371 9.3
R91 OUT_P.n374 OUT_P.n373 9.3
R92 OUT_P.n412 OUT_P.n411 9.3
R93 OUT_P.n392 OUT_P.n391 9.3
R94 OUT_P.n388 OUT_P.n387 9.3
R95 OUT_P.n384 OUT_P.n383 9.3
R96 OUT_P.n380 OUT_P.n379 9.3
R97 OUT_P.n398 OUT_P.n397 9.3
R98 OUT_P.n401 OUT_P.n400 9.3
R99 OUT_P.n403 OUT_P.n402 9.3
R100 OUT_P.n335 OUT_P.n334 9.3
R101 OUT_P.n848 OUT_P.n847 9.3
R102 OUT_P.n854 OUT_P.n853 9.3
R103 OUT_P.n844 OUT_P.n843 9.3
R104 OUT_P.n870 OUT_P.n869 9.3
R105 OUT_P.n864 OUT_P.n863 9.3
R106 OUT_P.n860 OUT_P.n859 9.3
R107 OUT_P.n838 OUT_P.n837 9.3
R108 OUT_P.n827 OUT_P.n826 9.3
R109 OUT_P.n829 OUT_P.n828 9.3
R110 OUT_P.n820 OUT_P.n819 9.3
R111 OUT_P.n834 OUT_P.n833 9.3
R112 OUT_P.n840 OUT_P.n839 9.3
R113 OUT_P.n850 OUT_P.n849 9.3
R114 OUT_P.n966 OUT_P.n965 9.3
R115 OUT_P.n956 OUT_P.n955 9.3
R116 OUT_P.n972 OUT_P.n971 9.3
R117 OUT_P.n950 OUT_P.n949 9.3
R118 OUT_P.n941 OUT_P.n940 9.3
R119 OUT_P.n939 OUT_P.n938 9.3
R120 OUT_P.n931 OUT_P.n930 9.3
R121 OUT_P.n935 OUT_P.n934 9.3
R122 OUT_P.n929 OUT_P.n928 9.3
R123 OUT_P.n922 OUT_P.n921 9.3
R124 OUT_P.n946 OUT_P.n945 9.3
R125 OUT_P.n952 OUT_P.n951 9.3
R126 OUT_P.n962 OUT_P.n961 9.3
R127 OUT_P.n1067 OUT_P.n1066 9.3
R128 OUT_P.n1057 OUT_P.n1056 9.3
R129 OUT_P.n1073 OUT_P.n1072 9.3
R130 OUT_P.n1051 OUT_P.n1050 9.3
R131 OUT_P.n1042 OUT_P.n1041 9.3
R132 OUT_P.n1040 OUT_P.n1039 9.3
R133 OUT_P.n1032 OUT_P.n1031 9.3
R134 OUT_P.n1036 OUT_P.n1035 9.3
R135 OUT_P.n1030 OUT_P.n1029 9.3
R136 OUT_P.n1023 OUT_P.n1022 9.3
R137 OUT_P.n1047 OUT_P.n1046 9.3
R138 OUT_P.n1053 OUT_P.n1052 9.3
R139 OUT_P.n1063 OUT_P.n1062 9.3
R140 OUT_P.n442 OUT_P.n441 9.3
R141 OUT_P.n489 OUT_P.n488 9.3
R142 OUT_P.n500 OUT_P.n499 9.3
R143 OUT_P.n523 OUT_P.n522 9.3
R144 OUT_P.n570 OUT_P.n569 9.3
R145 OUT_P.n582 OUT_P.n581 9.3
R146 OUT_P.n782 OUT_P.n781 9.3
R147 OUT_P.n616 OUT_P.n615 9.3
R148 OUT_P.n628 OUT_P.n627 9.3
R149 OUT_P.n677 OUT_P.n676 9.3
R150 OUT_P.n78 OUT_P.n44 9
R151 OUT_P.n68 OUT_P.n67 9
R152 OUT_P.n58 OUT_P.n45 9
R153 OUT_P.n21 OUT_P.n18 9
R154 OUT_P.n36 OUT_P.n35 9
R155 OUT_P.n49 OUT_P.n48 9
R156 OUT_P.n88 OUT_P.n43 9
R157 OUT_P.n171 OUT_P.n168 9
R158 OUT_P.n180 OUT_P.n167 9
R159 OUT_P.n189 OUT_P.n166 9
R160 OUT_P.n210 OUT_P.n165 9
R161 OUT_P.n141 OUT_P.n140 9
R162 OUT_P.n200 OUT_P.n199 9
R163 OUT_P.n126 OUT_P.n123 9
R164 OUT_P.n276 OUT_P.n273 9
R165 OUT_P.n285 OUT_P.n272 9
R166 OUT_P.n294 OUT_P.n271 9
R167 OUT_P.n315 OUT_P.n270 9
R168 OUT_P.n246 OUT_P.n245 9
R169 OUT_P.n305 OUT_P.n304 9
R170 OUT_P.n231 OUT_P.n228 9
R171 OUT_P.n381 OUT_P.n378 9
R172 OUT_P.n390 OUT_P.n377 9
R173 OUT_P.n399 OUT_P.n376 9
R174 OUT_P.n420 OUT_P.n375 9
R175 OUT_P.n351 OUT_P.n350 9
R176 OUT_P.n410 OUT_P.n409 9
R177 OUT_P.n336 OUT_P.n333 9
R178 OUT_P.n861 OUT_P.n807 9
R179 OUT_P.n872 OUT_P.n871 9
R180 OUT_P.n818 OUT_P.n813 9
R181 OUT_P.n825 OUT_P.n824 9
R182 OUT_P.n831 OUT_P.n830 9
R183 OUT_P.n841 OUT_P.n809 9
R184 OUT_P.n851 OUT_P.n808 9
R185 OUT_P.n920 OUT_P.n915 9
R186 OUT_P.n973 OUT_P.n908 9
R187 OUT_P.n932 OUT_P.n911 9
R188 OUT_P.n927 OUT_P.n926 9
R189 OUT_P.n943 OUT_P.n942 9
R190 OUT_P.n953 OUT_P.n910 9
R191 OUT_P.n963 OUT_P.n909 9
R192 OUT_P.n1021 OUT_P.n1016 9
R193 OUT_P.n1074 OUT_P.n1009 9
R194 OUT_P.n1033 OUT_P.n1012 9
R195 OUT_P.n1028 OUT_P.n1027 9
R196 OUT_P.n1044 OUT_P.n1043 9
R197 OUT_P.n1054 OUT_P.n1011 9
R198 OUT_P.n1064 OUT_P.n1010 9
R199 OUT_P.n566 OUT_P.n565 9
R200 OUT_P.n578 OUT_P.n577 9
R201 OUT_P.n519 OUT_P.n518 9
R202 OUT_P.n485 OUT_P.n484 9
R203 OUT_P.n496 OUT_P.n495 9
R204 OUT_P.n438 OUT_P.n437 9
R205 OUT_P.n778 OUT_P.n777 9
R206 OUT_P.n612 OUT_P.n611 9
R207 OUT_P.n624 OUT_P.n623 9
R208 OUT_P.n673 OUT_P.n672 9
R209 OUT_P.n1278 OUT_P.n1277 8.764
R210 OUT_P.n449 OUT_P.n448 8.764
R211 OUT_P.n1205 OUT_P.n1204 8.764
R212 OUT_P.n507 OUT_P.n506 8.764
R213 OUT_P.n1306 OUT_P.n1305 8.764
R214 OUT_P.n530 OUT_P.n529 8.764
R215 OUT_P.n1168 OUT_P.n1167 8.764
R216 OUT_P.n589 OUT_P.n588 8.764
R217 OUT_P.n789 OUT_P.n788 8.764
R218 OUT_P.n1232 OUT_P.n1231 8.764
R219 OUT_P.n1138 OUT_P.n1137 8.764
R220 OUT_P.n635 OUT_P.n634 8.764
R221 OUT_P.n684 OUT_P.n683 8.764
R222 OUT_P.n1329 OUT_P.n1328 8.764
R223 OUT_P.n15 OUT_P.n14 8.097
R224 OUT_P.n120 OUT_P.n119 8.097
R225 OUT_P.n225 OUT_P.n224 8.097
R226 OUT_P.n330 OUT_P.n329 8.097
R227 OUT_P.n1272 OUT_P.n1271 6.364
R228 OUT_P.n1198 OUT_P.n1197 6.364
R229 OUT_P.n1300 OUT_P.n1299 6.364
R230 OUT_P.n1161 OUT_P.n1160 6.364
R231 OUT_P.n1237 OUT_P.n1235 6.364
R232 OUT_P.n1131 OUT_P.n1130 6.364
R233 OUT_P.n1335 OUT_P.n2 6.364
R234 OUT_P.n32 OUT_P.n31 4.574
R235 OUT_P.n137 OUT_P.n136 4.574
R236 OUT_P.n242 OUT_P.n241 4.574
R237 OUT_P.n347 OUT_P.n346 4.574
R238 OUT_P.n822 OUT_P.n812 4.574
R239 OUT_P.n924 OUT_P.n914 4.574
R240 OUT_P.n1025 OUT_P.n1015 4.574
R241 OUT_P.n1279 OUT_P.n1278 4.574
R242 OUT_P.n1206 OUT_P.n1205 4.574
R243 OUT_P.n1307 OUT_P.n1306 4.574
R244 OUT_P.n1169 OUT_P.n1168 4.574
R245 OUT_P.n590 OUT_P.n589 4.574
R246 OUT_P.n531 OUT_P.n530 4.574
R247 OUT_P.n508 OUT_P.n507 4.574
R248 OUT_P.n450 OUT_P.n449 4.574
R249 OUT_P.n790 OUT_P.n789 4.574
R250 OUT_P.n1243 OUT_P.n1232 4.574
R251 OUT_P.n1139 OUT_P.n1138 4.574
R252 OUT_P.n636 OUT_P.n635 4.574
R253 OUT_P.n685 OUT_P.n684 4.574
R254 OUT_P.n1330 OUT_P.n1329 4.574
R255 OUT_P.n458 OUT_P.n457 4.559
R256 OUT_P.n539 OUT_P.n538 4.559
R257 OUT_P.n691 OUT_P.n667 4.559
R258 OUT_P.n795 OUT_P.n773 4.557
R259 OUT_P.n1325 OUT_P.n1324 4.554
R260 OUT_P.n1248 OUT_P.n1247 4.553
R261 OUT_P.n1211 OUT_P.n1210 4.553
R262 OUT_P.n1174 OUT_P.n1173 4.553
R263 OUT_P.n1142 OUT_P.n1126 4.553
R264 OUT_P.n1282 OUT_P.n1267 4.552
R265 OUT_P.n1310 OUT_P.n1295 4.552
R266 OUT_P.n774 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE 4.156
R267 OUT_P.n31 OUT_P.n29 3.388
R268 OUT_P.n136 OUT_P.n134 3.388
R269 OUT_P.n241 OUT_P.n239 3.388
R270 OUT_P.n346 OUT_P.n344 3.388
R271 OUT_P.n812 OUT_P.n811 3.388
R272 OUT_P.n914 OUT_P.n913 3.388
R273 OUT_P.n1015 OUT_P.n1014 3.388
R274 OUT_P.n15 OUT_P.t3 3.326
R275 OUT_P.n15 OUT_P.t1 3.326
R276 OUT_P.n120 OUT_P.t8 3.326
R277 OUT_P.n120 OUT_P.t10 3.326
R278 OUT_P.n225 OUT_P.t13 3.326
R279 OUT_P.n225 OUT_P.t6 3.326
R280 OUT_P.n330 OUT_P.t11 3.326
R281 OUT_P.n330 OUT_P.t7 3.326
R282 OUT_P.n814 OUT_P.t5 3.326
R283 OUT_P.n814 OUT_P.t0 3.326
R284 OUT_P.n916 OUT_P.t9 3.326
R285 OUT_P.n916 OUT_P.t4 3.326
R286 OUT_P.n1017 OUT_P.t12 3.326
R287 OUT_P.n1017 OUT_P.t2 3.326
R288 OUT_P.n593 OUT_P.n592 2.473
R289 OUT_P.n512 OUT_P.n511 2.473
R290 OUT_P.n639 OUT_P.n638 2.473
R291 OUT_P.n107 OUT_P.n89 2.473
R292 OUT_P.n338 OUT_P.n337 2.473
R293 OUT_P.n353 OUT_P.n352 2.473
R294 OUT_P.n422 OUT_P.n421 2.473
R295 OUT_P.n233 OUT_P.n232 2.473
R296 OUT_P.n248 OUT_P.n247 2.473
R297 OUT_P.n317 OUT_P.n316 2.473
R298 OUT_P.n128 OUT_P.n127 2.473
R299 OUT_P.n143 OUT_P.n142 2.473
R300 OUT_P.n212 OUT_P.n211 2.473
R301 OUT_P.n23 OUT_P.n22 2.473
R302 OUT_P.n38 OUT_P.n37 2.473
R303 OUT_P.n875 OUT_P.n874 1.813
R304 OUT_P.n976 OUT_P.n975 1.813
R305 OUT_P.n1077 OUT_P.n1076 1.813
R306 OUT_P.n1283 OUT_P.n1282 1.805
R307 OUT_P.n1311 OUT_P.n1310 1.805
R308 OUT_P.n1325 OUT_P.n1322 1.805
R309 OUT_P.n729 OUT_P.n548 1.705
R310 OUT_P.n724 OUT_P.n723 1.705
R311 OUT_P.n757 OUT_P.n467 1.705
R312 OUT_P.n752 OUT_P.n751 1.705
R313 OUT_P.n661 OUT_P.n660 1.705
R314 OUT_P.n701 OUT_P.n700 1.705
R315 OUT_P.n1322 OUT_P.n1321 1.705
R316 OUT_P.n1292 OUT_P.n1291 1.705
R317 OUT_P.n1320 OUT_P.n1319 1.705
R318 OUT_P.n668 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE 1.375
R319 OUT_P.n433 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/GATE 1.375
R320 OUT_P.n514 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/GATE 1.375
R321 OUT_P.n1265 OUT_P.n1264 1.329
R322 OUT_P.n796 OUT_P.n795 1.188
R323 OUT_P.n540 OUT_P.n539 1.187
R324 OUT_P.n459 OUT_P.n458 1.187
R325 OUT_P.n692 OUT_P.n691 1.187
R326 OUT_P.n1212 OUT_P.n1211 1.183
R327 OUT_P.n1175 OUT_P.n1174 1.183
R328 OUT_P.n1143 OUT_P.n1142 1.183
R329 OUT_P.n1249 OUT_P.n1248 1.183
R330 OUT_P.n16 OUT_P.n15 1.155
R331 OUT_P.n121 OUT_P.n120 1.155
R332 OUT_P.n226 OUT_P.n225 1.155
R333 OUT_P.n331 OUT_P.n330 1.155
R334 OUT_P.n815 OUT_P.n814 1.155
R335 OUT_P.n917 OUT_P.n916 1.155
R336 OUT_P.n1018 OUT_P.n1017 1.155
R337 OUT_P.n710 OUT_P.n709 1.137
R338 OUT_P.n738 OUT_P.n737 1.137
R339 OUT_P.n767 OUT_P.n766 1.137
R340 OUT_P.n804 OUT_P.n803 1.137
R341 OUT_P.n1256 OUT_P.n1255 1.137
R342 OUT_P.n1228 OUT_P.n1227 1.137
R343 OUT_P.n1219 OUT_P.n1218 1.137
R344 OUT_P.n1191 OUT_P.n1190 1.137
R345 OUT_P.n1182 OUT_P.n1181 1.137
R346 OUT_P.n1154 OUT_P.n1153 1.137
R347 OUT_P.n1145 OUT_P.n1144 1.137
R348 OUT_P.n647 OUT_P.n646 1.137
R349 OUT_P.n1104 OUT_P.n1103 1.133
R350 OUT_P.n1003 OUT_P.n1002 1.133
R351 OUT_P.n902 OUT_P.n901 1.133
R352 OUT_P.n1262 OUT_P.n432 1.133
R353 OUT_P.n426 OUT_P.n425 1.133
R354 OUT_P.n321 OUT_P.n320 1.133
R355 OUT_P.n216 OUT_P.n215 1.133
R356 OUT_P.n111 OUT_P.n110 1.133
R357 OUT_P.n1263 OUT_P.n11 1.133
R358 OUT_P.n1258 OUT_P.n1257 1.059
R359 OUT_P.n774 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE 1
R360 OUT_P.n17 OUT_P.n16 0.893
R361 OUT_P.n122 OUT_P.n121 0.893
R362 OUT_P.n227 OUT_P.n226 0.893
R363 OUT_P.n332 OUT_P.n331 0.893
R364 OUT_P.n816 OUT_P.n815 0.893
R365 OUT_P.n918 OUT_P.n917 0.893
R366 OUT_P.n1019 OUT_P.n1018 0.893
R367 OUT_P.n1123 OUT_P.n1122 0.868
R368 OUT_P.n1261 OUT_P.n1111 0.853
R369 OUT_P.n1271 OUT_P.n1270 0.77
R370 OUT_P.n441 OUT_P.n440 0.77
R371 OUT_P.n1197 OUT_P.n1196 0.77
R372 OUT_P.n488 OUT_P.n487 0.77
R373 OUT_P.n499 OUT_P.n498 0.77
R374 OUT_P.n1299 OUT_P.n1298 0.77
R375 OUT_P.n522 OUT_P.n521 0.77
R376 OUT_P.n1160 OUT_P.n1159 0.77
R377 OUT_P.n569 OUT_P.n568 0.77
R378 OUT_P.n581 OUT_P.n580 0.77
R379 OUT_P.n781 OUT_P.n780 0.77
R380 OUT_P.n1235 OUT_P.n1234 0.77
R381 OUT_P.n1130 OUT_P.n1129 0.77
R382 OUT_P.n615 OUT_P.n614 0.77
R383 OUT_P.n627 OUT_P.n626 0.77
R384 OUT_P.n676 OUT_P.n675 0.77
R385 OUT_P.n2 OUT_P.n1 0.77
R386 OUT_P.n492 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/GATE 0.666
R387 OUT_P.n717 OUT_P.n716 0.65
R388 OUT_P.n654 OUT_P.n653 0.65
R389 OUT_P.n745 OUT_P.n744 0.645
R390 OUT_P.n31 OUT_P.n30 0.506
R391 OUT_P.n136 OUT_P.n135 0.506
R392 OUT_P.n241 OUT_P.n240 0.506
R393 OUT_P.n346 OUT_P.n345 0.506
R394 OUT_P.n812 OUT_P.n810 0.506
R395 OUT_P.n914 OUT_P.n912 0.506
R396 OUT_P.n1015 OUT_P.n1013 0.506
R397 OUT_P.n86 OUT_P.n85 0.476
R398 OUT_P.n208 OUT_P.n207 0.476
R399 OUT_P.n313 OUT_P.n312 0.476
R400 OUT_P.n418 OUT_P.n417 0.476
R401 OUT_P.n833 OUT_P.n832 0.476
R402 OUT_P.n934 OUT_P.n933 0.476
R403 OUT_P.n1035 OUT_P.n1034 0.476
R404 OUT_P.n1293 OUT_P.n1292 0.456
R405 OUT_P.n1321 OUT_P.n1320 0.456
R406 OUT_P.n1221 OUT_P.n1220 0.45
R407 OUT_P.n1184 OUT_P.n1183 0.45
R408 OUT_P.n1147 OUT_P.n1146 0.45
R409 OUT_P.n76 OUT_P.n75 0.445
R410 OUT_P.n197 OUT_P.n196 0.445
R411 OUT_P.n302 OUT_P.n301 0.445
R412 OUT_P.n407 OUT_P.n406 0.445
R413 OUT_P.n843 OUT_P.n842 0.445
R414 OUT_P.n945 OUT_P.n944 0.445
R415 OUT_P.n1046 OUT_P.n1045 0.445
R416 OUT_P.n1111 OUT_P.n805 0.43
R417 OUT_P.n65 OUT_P.n64 0.414
R418 OUT_P.n187 OUT_P.n186 0.414
R419 OUT_P.n292 OUT_P.n291 0.414
R420 OUT_P.n397 OUT_P.n396 0.414
R421 OUT_P.n853 OUT_P.n852 0.414
R422 OUT_P.n955 OUT_P.n954 0.414
R423 OUT_P.n1056 OUT_P.n1055 0.414
R424 OUT_P.n863 OUT_P.n862 0.382
R425 OUT_P.n965 OUT_P.n964 0.382
R426 OUT_P.n1066 OUT_P.n1065 0.382
R427 OUT_P.n731 OUT_P.n730 0.294
R428 OUT_P.n759 OUT_P.n758 0.294
R429 OUT_P.n703 OUT_P.n702 0.292
R430 OUT_P.n1109 OUT_P.n1108 0.262
R431 OUT_P.n1262 OUT_P.n1261 0.175
R432 OUT_P.n1008 OUT_P.n1007 0.163
R433 OUT_P.n907 OUT_P.n906 0.163
R434 OUT_P.n326 OUT_P.n325 0.163
R435 OUT_P.n221 OUT_P.n220 0.163
R436 OUT_P.n116 OUT_P.n115 0.163
R437 OUT_P.n431 OUT_P.n430 0.159
R438 OUT_P.n1292 OUT_P.n1265 0.088
R439 OUT_P.n1320 OUT_P.n1293 0.088
R440 OUT_P.n11 OUT_P 0.065
R441 OUT_P.n83 OUT_P.n82 0.06
R442 OUT_P.n73 OUT_P.n72 0.06
R443 OUT_P.n62 OUT_P.n61 0.06
R444 OUT_P.n54 OUT_P.n53 0.06
R445 OUT_P.n205 OUT_P.n204 0.06
R446 OUT_P.n194 OUT_P.n193 0.06
R447 OUT_P.n184 OUT_P.n183 0.06
R448 OUT_P.n176 OUT_P.n175 0.06
R449 OUT_P.n310 OUT_P.n309 0.06
R450 OUT_P.n299 OUT_P.n298 0.06
R451 OUT_P.n289 OUT_P.n288 0.06
R452 OUT_P.n281 OUT_P.n280 0.06
R453 OUT_P.n415 OUT_P.n414 0.06
R454 OUT_P.n404 OUT_P.n403 0.06
R455 OUT_P.n394 OUT_P.n393 0.06
R456 OUT_P.n386 OUT_P.n385 0.06
R457 OUT_P.n857 OUT_P.n856 0.06
R458 OUT_P.n848 OUT_P.n846 0.06
R459 OUT_P.n838 OUT_P.n836 0.06
R460 OUT_P.n959 OUT_P.n958 0.06
R461 OUT_P.n950 OUT_P.n948 0.06
R462 OUT_P.n939 OUT_P.n937 0.06
R463 OUT_P.n1060 OUT_P.n1059 0.06
R464 OUT_P.n1051 OUT_P.n1049 0.06
R465 OUT_P.n1040 OUT_P.n1038 0.06
R466 OUT_P.n1230 OUT_P.n1229 0.055
R467 OUT_P.n1193 OUT_P.n1192 0.055
R468 OUT_P.n1156 OUT_P.n1155 0.055
R469 OUT_P.n1124 OUT_P.n1123 0.055
R470 OUT_P.n825 OUT_P.n823 0.053
R471 OUT_P.n823 OUT_P.n822 0.053
R472 OUT_P.n927 OUT_P.n925 0.053
R473 OUT_P.n925 OUT_P.n924 0.053
R474 OUT_P.n1028 OUT_P.n1026 0.053
R475 OUT_P.n1026 OUT_P.n1025 0.053
R476 OUT_P.n867 OUT_P.n866 0.052
R477 OUT_P.n969 OUT_P.n968 0.052
R478 OUT_P.n1070 OUT_P.n1069 0.052
R479 OUT_P.n1141 OUT_P.n1140 0.051
R480 OUT_P.n1136 OUT_P.n1135 0.051
R481 OUT_P.n1281 OUT_P.n1280 0.051
R482 OUT_P.n1276 OUT_P.n1275 0.051
R483 OUT_P.n1208 OUT_P.n1207 0.051
R484 OUT_P.n1203 OUT_P.n1202 0.051
R485 OUT_P.n1309 OUT_P.n1308 0.051
R486 OUT_P.n1304 OUT_P.n1303 0.051
R487 OUT_P.n1171 OUT_P.n1170 0.051
R488 OUT_P.n1166 OUT_P.n1165 0.051
R489 OUT_P.n1245 OUT_P.n1244 0.051
R490 OUT_P.n1242 OUT_P.n1241 0.051
R491 OUT_P.n1327 OUT_P.n1326 0.051
R492 OUT_P.n1332 OUT_P.n1331 0.051
R493 OUT_P.n690 OUT_P.n689 0.048
R494 OUT_P.n681 OUT_P.n680 0.048
R495 OUT_P.n794 OUT_P.n793 0.048
R496 OUT_P.n786 OUT_P.n785 0.048
R497 OUT_P.n455 OUT_P.n454 0.048
R498 OUT_P.n446 OUT_P.n445 0.048
R499 OUT_P.n511 OUT_P.n491 0.048
R500 OUT_P.n504 OUT_P.n503 0.048
R501 OUT_P.n536 OUT_P.n535 0.048
R502 OUT_P.n527 OUT_P.n526 0.048
R503 OUT_P.n592 OUT_P.n573 0.048
R504 OUT_P.n586 OUT_P.n585 0.048
R505 OUT_P.n638 OUT_P.n619 0.048
R506 OUT_P.n632 OUT_P.n631 0.048
R507 OUT_P.n34 OUT_P.n33 0.045
R508 OUT_P.n87 OUT_P.n84 0.045
R509 OUT_P.n139 OUT_P.n138 0.045
R510 OUT_P.n209 OUT_P.n206 0.045
R511 OUT_P.n244 OUT_P.n243 0.045
R512 OUT_P.n314 OUT_P.n311 0.045
R513 OUT_P.n349 OUT_P.n348 0.045
R514 OUT_P.n419 OUT_P.n416 0.045
R515 OUT_P.n22 OUT_P.n21 0.043
R516 OUT_P.n56 OUT_P.n54 0.043
R517 OUT_P.n127 OUT_P.n126 0.043
R518 OUT_P.n178 OUT_P.n176 0.043
R519 OUT_P.n232 OUT_P.n231 0.043
R520 OUT_P.n283 OUT_P.n281 0.043
R521 OUT_P.n337 OUT_P.n336 0.043
R522 OUT_P.n388 OUT_P.n386 0.043
R523 OUT_P.n818 OUT_P.n817 0.043
R524 OUT_P.n920 OUT_P.n919 0.043
R525 OUT_P.n1021 OUT_P.n1020 0.043
R526 OUT_P.n1326 OUT_P.n1325 0.041
R527 OUT_P.n1282 OUT_P.n1281 0.041
R528 OUT_P.n1310 OUT_P.n1309 0.041
R529 OUT_P.n1139 OUT_P.n1136 0.04
R530 OUT_P.n835 OUT_P.n834 0.04
R531 OUT_P.n936 OUT_P.n935 0.04
R532 OUT_P.n1037 OUT_P.n1036 0.04
R533 OUT_P.n1279 OUT_P.n1276 0.04
R534 OUT_P.n1214 OUT_P.n1213 0.04
R535 OUT_P.n1206 OUT_P.n1203 0.04
R536 OUT_P.n1307 OUT_P.n1304 0.04
R537 OUT_P.n1177 OUT_P.n1176 0.04
R538 OUT_P.n1169 OUT_P.n1166 0.04
R539 OUT_P.n1243 OUT_P.n1242 0.04
R540 OUT_P.n1251 OUT_P.n1250 0.04
R541 OUT_P.n1119 OUT_P.n1118 0.04
R542 OUT_P.n1331 OUT_P.n1330 0.04
R543 OUT_P.n1248 OUT_P.n1245 0.039
R544 OUT_P.n1142 OUT_P.n1141 0.039
R545 OUT_P.n1211 OUT_P.n1208 0.039
R546 OUT_P.n1174 OUT_P.n1171 0.039
R547 OUT_P.n37 OUT_P.n36 0.038
R548 OUT_P.n142 OUT_P.n141 0.038
R549 OUT_P.n247 OUT_P.n246 0.038
R550 OUT_P.n352 OUT_P.n351 0.038
R551 OUT_P.n1140 OUT_P.n1139 0.038
R552 OUT_P.n1280 OUT_P.n1279 0.038
R553 OUT_P.n1215 OUT_P.n1214 0.038
R554 OUT_P.n1207 OUT_P.n1206 0.038
R555 OUT_P.n1308 OUT_P.n1307 0.038
R556 OUT_P.n1178 OUT_P.n1177 0.038
R557 OUT_P.n1170 OUT_P.n1169 0.038
R558 OUT_P.n1244 OUT_P.n1243 0.038
R559 OUT_P.n1252 OUT_P.n1251 0.038
R560 OUT_P.n1118 OUT_P.n1117 0.038
R561 OUT_P.n1330 OUT_P.n1327 0.038
R562 OUT_P.n63 OUT_P.n62 0.036
R563 OUT_P.n185 OUT_P.n184 0.036
R564 OUT_P.n290 OUT_P.n289 0.036
R565 OUT_P.n395 OUT_P.n394 0.036
R566 OUT_P.n856 OUT_P.n855 0.036
R567 OUT_P.n958 OUT_P.n957 0.036
R568 OUT_P.n1059 OUT_P.n1058 0.036
R569 OUT_P.n1275 OUT_P.n1274 0.036
R570 OUT_P.n1303 OUT_P.n1302 0.036
R571 OUT_P.n1333 OUT_P.n1332 0.036
R572 OUT_P.n1216 OUT_P.n1215 0.034
R573 OUT_P.n1179 OUT_P.n1178 0.034
R574 OUT_P.n1253 OUT_P.n1252 0.034
R575 OUT_P.n1117 OUT_P.n1116 0.034
R576 OUT_P.n1135 OUT_P.n1134 0.033
R577 OUT_P.n1202 OUT_P.n1201 0.033
R578 OUT_P.n1165 OUT_P.n1164 0.033
R579 OUT_P.n1241 OUT_P.n1240 0.033
R580 OUT_P.n1120 OUT_P.n1119 0.033
R581 OUT_P.n688 OUT_P.n687 0.032
R582 OUT_P.n793 OUT_P.n792 0.032
R583 OUT_P.n453 OUT_P.n452 0.032
R584 OUT_P.n511 OUT_P.n510 0.032
R585 OUT_P.n534 OUT_P.n533 0.032
R586 OUT_P.n545 OUT_P.n544 0.032
R587 OUT_P.n512 OUT_P.n480 0.032
R588 OUT_P.n464 OUT_P.n463 0.032
R589 OUT_P.n801 OUT_P.n800 0.032
R590 OUT_P.n697 OUT_P.n696 0.032
R591 OUT_P.n691 OUT_P.n690 0.031
R592 OUT_P.n458 OUT_P.n455 0.031
R593 OUT_P.n539 OUT_P.n536 0.031
R594 OUT_P.n80 OUT_P.n78 0.031
R595 OUT_P.n202 OUT_P.n200 0.031
R596 OUT_P.n307 OUT_P.n305 0.031
R597 OUT_P.n412 OUT_P.n410 0.031
R598 OUT_P.n872 OUT_P.n870 0.031
R599 OUT_P.n841 OUT_P.n840 0.031
R600 OUT_P.n831 OUT_P.n829 0.031
R601 OUT_P.n973 OUT_P.n972 0.031
R602 OUT_P.n943 OUT_P.n941 0.031
R603 OUT_P.n932 OUT_P.n931 0.031
R604 OUT_P.n1074 OUT_P.n1073 0.031
R605 OUT_P.n1044 OUT_P.n1042 0.031
R606 OUT_P.n1033 OUT_P.n1032 0.031
R607 OUT_P.n795 OUT_P.n794 0.031
R608 OUT_P.n592 OUT_P.n591 0.03
R609 OUT_P.n590 OUT_P.n587 0.03
R610 OUT_P.n593 OUT_P.n562 0.03
R611 OUT_P.n561 OUT_P.n560 0.03
R612 OUT_P.n638 OUT_P.n637 0.03
R613 OUT_P.n636 OUT_P.n633 0.03
R614 OUT_P.n639 OUT_P.n608 0.03
R615 OUT_P.n607 OUT_P.n606 0.03
R616 OUT_P.n1131 OUT_P.n1127 0.029
R617 OUT_P.n1198 OUT_P.n1194 0.029
R618 OUT_P.n1161 OUT_P.n1157 0.029
R619 OUT_P.n1237 OUT_P.n1236 0.029
R620 OUT_P.n1272 OUT_P.n1268 0.028
R621 OUT_P.n1300 OUT_P.n1296 0.028
R622 OUT_P.n1336 OUT_P.n1335 0.028
R623 OUT_P.n685 OUT_P.n682 0.028
R624 OUT_P.n866 OUT_P.n865 0.028
R625 OUT_P.n968 OUT_P.n967 0.028
R626 OUT_P.n1069 OUT_P.n1068 0.028
R627 OUT_P.n450 OUT_P.n447 0.028
R628 OUT_P.n531 OUT_P.n528 0.028
R629 OUT_P.n513 OUT_P.n512 0.028
R630 OUT_P.n802 OUT_P.n801 0.028
R631 OUT_P.n1122 OUT_P.n1121 0.027
R632 OUT_P.n1218 OUT_P.n1217 0.027
R633 OUT_P.n1181 OUT_P.n1180 0.027
R634 OUT_P.n1255 OUT_P.n1254 0.027
R635 OUT_P.n77 OUT_P.n74 0.026
R636 OUT_P.n74 OUT_P.n73 0.026
R637 OUT_P.n70 OUT_P.n68 0.026
R638 OUT_P.n60 OUT_P.n58 0.026
R639 OUT_P.n198 OUT_P.n195 0.026
R640 OUT_P.n195 OUT_P.n194 0.026
R641 OUT_P.n191 OUT_P.n189 0.026
R642 OUT_P.n182 OUT_P.n180 0.026
R643 OUT_P.n303 OUT_P.n300 0.026
R644 OUT_P.n300 OUT_P.n299 0.026
R645 OUT_P.n296 OUT_P.n294 0.026
R646 OUT_P.n287 OUT_P.n285 0.026
R647 OUT_P.n408 OUT_P.n405 0.026
R648 OUT_P.n405 OUT_P.n404 0.026
R649 OUT_P.n401 OUT_P.n399 0.026
R650 OUT_P.n392 OUT_P.n390 0.026
R651 OUT_P.n644 OUT_P.n643 0.026
R652 OUT_P.n861 OUT_P.n860 0.026
R653 OUT_P.n851 OUT_P.n850 0.026
R654 OUT_P.n846 OUT_P.n845 0.026
R655 OUT_P.n845 OUT_P.n844 0.026
R656 OUT_P.n887 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/DRAIN 0.026
R657 OUT_P.n963 OUT_P.n962 0.026
R658 OUT_P.n953 OUT_P.n952 0.026
R659 OUT_P.n948 OUT_P.n947 0.026
R660 OUT_P.n947 OUT_P.n946 0.026
R661 OUT_P.n988 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/DRAIN 0.026
R662 OUT_P.n1064 OUT_P.n1063 0.026
R663 OUT_P.n1054 OUT_P.n1053 0.026
R664 OUT_P.n1049 OUT_P.n1048 0.026
R665 OUT_P.n1048 OUT_P.n1047 0.026
R666 OUT_P.n1089 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/DRAIN 0.026
R667 OUT_P.n584 OUT_P.n583 0.026
R668 OUT_P.n664 OUT_P.n663 0.026
R669 OUT_P.n707 OUT_P.n706 0.026
R670 OUT_P.n555 OUT_P.n554 0.026
R671 OUT_P.n547 OUT_P.n546 0.026
R672 OUT_P.n727 OUT_P.n726 0.026
R673 OUT_P.n735 OUT_P.n734 0.026
R674 OUT_P.n466 OUT_P.n465 0.026
R675 OUT_P.n755 OUT_P.n754 0.026
R676 OUT_P.n770 OUT_P.n769 0.026
R677 OUT_P.n630 OUT_P.n629 0.026
R678 OUT_P.n601 OUT_P.n600 0.026
R679 OUT_P.n699 OUT_P.n698 0.026
R680 OUT_P.n790 OUT_P.n787 0.025
R681 OUT_P.n1190 OUT_P.n1186 0.025
R682 OUT_P.n508 OUT_P.n505 0.025
R683 OUT_P.n1153 OUT_P.n1149 0.025
R684 OUT_P.n478 OUT_P.n477 0.025
R685 OUT_P.n1227 OUT_P.n1223 0.025
R686 OUT_P.n776 OUT_P.n775 0.025
R687 OUT_P.n494 OUT_P.n493 0.025
R688 OUT_P.n53 OUT_P.n52 0.024
R689 OUT_P.n52 OUT_P.n50 0.024
R690 OUT_P.n175 OUT_P.n174 0.024
R691 OUT_P.n174 OUT_P.n172 0.024
R692 OUT_P.n280 OUT_P.n279 0.024
R693 OUT_P.n279 OUT_P.n277 0.024
R694 OUT_P.n385 OUT_P.n384 0.024
R695 OUT_P.n384 OUT_P.n382 0.024
R696 OUT_P.n870 OUT_P.n868 0.024
R697 OUT_P.n972 OUT_P.n970 0.024
R698 OUT_P.n1073 OUT_P.n1071 0.024
R699 OUT_P.n104 OUT_P.n103 0.023
R700 OUT_P.n101 OUT_P.n100 0.023
R701 OUT_P.n158 OUT_P.n157 0.023
R702 OUT_P.n155 OUT_P.n154 0.023
R703 OUT_P.n263 OUT_P.n262 0.023
R704 OUT_P.n260 OUT_P.n259 0.023
R705 OUT_P.n368 OUT_P.n367 0.023
R706 OUT_P.n365 OUT_P.n364 0.023
R707 OUT_P.n896 OUT_P.n895 0.023
R708 OUT_P.n997 OUT_P.n996 0.023
R709 OUT_P.n1098 OUT_P.n1097 0.023
R710 OUT_P.n594 OUT_P.n593 0.023
R711 OUT_P.n557 OUT_P.n556 0.023
R712 OUT_P.n640 OUT_P.n639 0.023
R713 OUT_P.n603 OUT_P.n602 0.023
R714 OUT_P.n32 OUT_P.n28 0.021
R715 OUT_P.n137 OUT_P.n133 0.021
R716 OUT_P.n242 OUT_P.n238 0.021
R717 OUT_P.n347 OUT_P.n343 0.021
R718 OUT_P.n679 OUT_P.n678 0.021
R719 OUT_P.n784 OUT_P.n783 0.021
R720 OUT_P.n822 OUT_P.n821 0.021
R721 OUT_P.n924 OUT_P.n923 0.021
R722 OUT_P.n1025 OUT_P.n1024 0.021
R723 OUT_P.n444 OUT_P.n443 0.021
R724 OUT_P.n483 OUT_P.n482 0.021
R725 OUT_P.n502 OUT_P.n501 0.021
R726 OUT_P.n525 OUT_P.n524 0.021
R727 OUT_P.n559 OUT_P.n558 0.021
R728 OUT_P.n721 OUT_P.n720 0.021
R729 OUT_P.n718 OUT_P.n717 0.021
R730 OUT_P.n743 OUT_P.n742 0.021
R731 OUT_P.n741 OUT_P.n740 0.021
R732 OUT_P.n472 OUT_P.n471 0.021
R733 OUT_P.n749 OUT_P.n748 0.021
R734 OUT_P.n746 OUT_P.n745 0.021
R735 OUT_P.n764 OUT_P.n763 0.021
R736 OUT_P.n605 OUT_P.n604 0.021
R737 OUT_P.n658 OUT_P.n657 0.021
R738 OUT_P.n655 OUT_P.n654 0.021
R739 OUT_P.n1261 OUT_P.n1260 0.02
R740 OUT_P.n22 OUT_P.n17 0.019
R741 OUT_P.n89 OUT_P.n42 0.019
R742 OUT_P.n61 OUT_P.n60 0.019
R743 OUT_P.n127 OUT_P.n122 0.019
R744 OUT_P.n211 OUT_P.n164 0.019
R745 OUT_P.n183 OUT_P.n182 0.019
R746 OUT_P.n232 OUT_P.n227 0.019
R747 OUT_P.n316 OUT_P.n269 0.019
R748 OUT_P.n288 OUT_P.n287 0.019
R749 OUT_P.n337 OUT_P.n332 0.019
R750 OUT_P.n421 OUT_P.n374 0.019
R751 OUT_P.n393 OUT_P.n392 0.019
R752 OUT_P.n827 OUT_P.n825 0.019
R753 OUT_P.n821 OUT_P.n820 0.019
R754 OUT_P.n817 OUT_P.n816 0.019
R755 OUT_P.n929 OUT_P.n927 0.019
R756 OUT_P.n923 OUT_P.n922 0.019
R757 OUT_P.n919 OUT_P.n918 0.019
R758 OUT_P.n1030 OUT_P.n1028 0.019
R759 OUT_P.n1024 OUT_P.n1023 0.019
R760 OUT_P.n1020 OUT_P.n1019 0.019
R761 OUT_P.n566 OUT_P.n564 0.019
R762 OUT_P.n572 OUT_P.n571 0.019
R763 OUT_P.n715 OUT_P.n714 0.019
R764 OUT_P.n713 OUT_P.n712 0.019
R765 OUT_P.n612 OUT_P.n610 0.019
R766 OUT_P.n618 OUT_P.n617 0.019
R767 OUT_P.n652 OUT_P.n651 0.019
R768 OUT_P.n650 OUT_P.n649 0.019
R769 OUT_P.n1186 OUT_P.n1185 0.018
R770 OUT_P.n1149 OUT_P.n1148 0.018
R771 OUT_P.n1223 OUT_P.n1222 0.018
R772 OUT_P.n1121 OUT_P.n1120 0.018
R773 OUT_P.n1285 OUT_P.n1284 0.017
R774 OUT_P.n1288 OUT_P.n1287 0.017
R775 OUT_P.n490 OUT_P.n489 0.017
R776 OUT_P.n1313 OUT_P.n1312 0.017
R777 OUT_P.n1316 OUT_P.n1315 0.017
R778 OUT_P.n710 OUT_P.n594 0.017
R779 OUT_P.n551 OUT_P.n550 0.017
R780 OUT_P.n474 OUT_P.n473 0.017
R781 OUT_P.n470 OUT_P.n469 0.017
R782 OUT_P.n766 OUT_P.n765 0.017
R783 OUT_P.n647 OUT_P.n640 0.017
R784 OUT_P.n597 OUT_P.n596 0.017
R785 OUT_P.n10 OUT_P.n9 0.017
R786 OUT_P.n7 OUT_P.n6 0.017
R787 OUT_P.n37 OUT_P.n34 0.016
R788 OUT_P.n142 OUT_P.n139 0.016
R789 OUT_P.n247 OUT_P.n244 0.016
R790 OUT_P.n352 OUT_P.n349 0.016
R791 OUT_P.n671 OUT_P.n670 0.016
R792 OUT_P.n836 OUT_P.n835 0.016
R793 OUT_P.n937 OUT_P.n936 0.016
R794 OUT_P.n1038 OUT_P.n1037 0.016
R795 OUT_P.n436 OUT_P.n435 0.016
R796 OUT_P.n1217 OUT_P.n1216 0.016
R797 OUT_P.n491 OUT_P.n490 0.016
R798 OUT_P.n517 OUT_P.n516 0.016
R799 OUT_P.n1180 OUT_P.n1179 0.016
R800 OUT_P.n573 OUT_P.n572 0.016
R801 OUT_P.n574 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/GATE 0.016
R802 OUT_P.n712 OUT_P.n711 0.016
R803 OUT_P.n723 OUT_P.n722 0.016
R804 OUT_P.n740 OUT_P.n739 0.016
R805 OUT_P.n476 OUT_P.n475 0.016
R806 OUT_P.n751 OUT_P.n750 0.016
R807 OUT_P.n797 OUT_P.n796 0.016
R808 OUT_P.n762 OUT_P.n761 0.016
R809 OUT_P.n1254 OUT_P.n1253 0.016
R810 OUT_P.n1256 OUT_P.n1230 0.016
R811 OUT_P.n1229 OUT_P.n1228 0.016
R812 OUT_P.n1219 OUT_P.n1193 0.016
R813 OUT_P.n1192 OUT_P.n1191 0.016
R814 OUT_P.n1182 OUT_P.n1156 0.016
R815 OUT_P.n1155 OUT_P.n1154 0.016
R816 OUT_P.n1145 OUT_P.n1124 0.016
R817 OUT_P.n1116 OUT_P.n1115 0.016
R818 OUT_P.n619 OUT_P.n618 0.016
R819 OUT_P.n620 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/GATE 0.016
R820 OUT_P.n649 OUT_P.n648 0.016
R821 OUT_P.n660 OUT_P.n659 0.016
R822 OUT_P.n775 OUT_P.n774 0.014
R823 OUT_P.n493 OUT_P.n492 0.014
R824 OUT_P.n21 OUT_P.n20 0.014
R825 OUT_P.n72 OUT_P.n70 0.014
R826 OUT_P.n68 OUT_P.n66 0.014
R827 OUT_P.n126 OUT_P.n125 0.014
R828 OUT_P.n193 OUT_P.n191 0.014
R829 OUT_P.n189 OUT_P.n188 0.014
R830 OUT_P.n231 OUT_P.n230 0.014
R831 OUT_P.n298 OUT_P.n296 0.014
R832 OUT_P.n294 OUT_P.n293 0.014
R833 OUT_P.n336 OUT_P.n335 0.014
R834 OUT_P.n403 OUT_P.n401 0.014
R835 OUT_P.n399 OUT_P.n398 0.014
R836 OUT_P.n669 OUT_P.n668 0.014
R837 OUT_P.n783 OUT_P.n782 0.014
R838 OUT_P.n865 OUT_P.n864 0.014
R839 OUT_P.n864 OUT_P.n861 0.014
R840 OUT_P.n854 OUT_P.n851 0.014
R841 OUT_P.n850 OUT_P.n848 0.014
R842 OUT_P.n820 OUT_P.n818 0.014
R843 OUT_P.n899 OUT_P.n898 0.014
R844 OUT_P.n967 OUT_P.n966 0.014
R845 OUT_P.n966 OUT_P.n963 0.014
R846 OUT_P.n956 OUT_P.n953 0.014
R847 OUT_P.n952 OUT_P.n950 0.014
R848 OUT_P.n922 OUT_P.n920 0.014
R849 OUT_P.n1000 OUT_P.n999 0.014
R850 OUT_P.n1068 OUT_P.n1067 0.014
R851 OUT_P.n1067 OUT_P.n1064 0.014
R852 OUT_P.n1057 OUT_P.n1054 0.014
R853 OUT_P.n1053 OUT_P.n1051 0.014
R854 OUT_P.n1023 OUT_P.n1021 0.014
R855 OUT_P.n1101 OUT_P.n1100 0.014
R856 OUT_P.n1108 OUT_P.n1107 0.014
R857 OUT_P.n1007 OUT_P.n1006 0.014
R858 OUT_P.n906 OUT_P.n905 0.014
R859 OUT_P.n1287 OUT_P.n1286 0.014
R860 OUT_P.n1268 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/GATE 0.014
R861 OUT_P.n434 OUT_P.n433 0.014
R862 OUT_P.n501 OUT_P.n500 0.014
R863 OUT_P.n1315 OUT_P.n1314 0.014
R864 OUT_P.n1296 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/GATE 0.014
R865 OUT_P.n515 OUT_P.n514 0.014
R866 OUT_P.n576 OUT_P.n575 0.014
R867 OUT_P.n716 OUT_P.n715 0.014
R868 OUT_P.n541 OUT_P.n540 0.014
R869 OUT_P.n548 OUT_P.n541 0.014
R870 OUT_P.n723 OUT_P.n551 0.014
R871 OUT_P.n720 OUT_P.n719 0.014
R872 OUT_P.n744 OUT_P.n743 0.014
R873 OUT_P.n475 OUT_P.n474 0.014
R874 OUT_P.n460 OUT_P.n459 0.014
R875 OUT_P.n467 OUT_P.n460 0.014
R876 OUT_P.n751 OUT_P.n470 0.014
R877 OUT_P.n748 OUT_P.n747 0.014
R878 OUT_P.n766 OUT_P.n762 0.014
R879 OUT_P.n622 OUT_P.n621 0.014
R880 OUT_P.n653 OUT_P.n652 0.014
R881 OUT_P.n693 OUT_P.n692 0.014
R882 OUT_P.n700 OUT_P.n693 0.014
R883 OUT_P.n660 OUT_P.n597 0.014
R884 OUT_P.n657 OUT_P.n656 0.014
R885 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE OUT_P.n1336 0.014
R886 OUT_P.n8 OUT_P.n7 0.014
R887 OUT_P.n430 OUT_P.n429 0.014
R888 OUT_P.n325 OUT_P.n324 0.014
R889 OUT_P.n220 OUT_P.n219 0.014
R890 OUT_P.n115 OUT_P.n114 0.014
R891 OUT_P.n1105 OUT_P.n1104 0.014
R892 OUT_P.n1004 OUT_P.n1003 0.014
R893 OUT_P.n903 OUT_P.n902 0.014
R894 OUT_P.n1263 OUT_P.n1262 0.014
R895 OUT_P.n427 OUT_P.n426 0.014
R896 OUT_P.n322 OUT_P.n321 0.014
R897 OUT_P.n217 OUT_P.n216 0.014
R898 OUT_P.n112 OUT_P.n111 0.014
R899 OUT_P.n98 OUT_P.n97 0.013
R900 OUT_P.n94 OUT_P.n93 0.013
R901 OUT_P.n152 OUT_P.n151 0.013
R902 OUT_P.n148 OUT_P.n147 0.013
R903 OUT_P.n257 OUT_P.n256 0.013
R904 OUT_P.n253 OUT_P.n252 0.013
R905 OUT_P.n362 OUT_P.n361 0.013
R906 OUT_P.n358 OUT_P.n357 0.013
R907 OUT_P.n1127 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/GATE 0.013
R908 OUT_P.n1286 OUT_P.n1285 0.013
R909 OUT_P.n1194 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/GATE 0.013
R910 OUT_P.n1314 OUT_P.n1313 0.013
R911 OUT_P.n1157 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/GATE 0.013
R912 OUT_P.n1236 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE 0.013
R913 OUT_P.n9 OUT_P.n8 0.013
R914 OUT_P.n89 OUT_P.n88 0.012
R915 OUT_P.n84 OUT_P.n83 0.012
R916 OUT_P.n66 OUT_P.n63 0.012
R917 OUT_P.n58 OUT_P.n57 0.012
R918 OUT_P.n211 OUT_P.n210 0.012
R919 OUT_P.n206 OUT_P.n205 0.012
R920 OUT_P.n188 OUT_P.n185 0.012
R921 OUT_P.n180 OUT_P.n179 0.012
R922 OUT_P.n316 OUT_P.n315 0.012
R923 OUT_P.n311 OUT_P.n310 0.012
R924 OUT_P.n293 OUT_P.n290 0.012
R925 OUT_P.n285 OUT_P.n284 0.012
R926 OUT_P.n421 OUT_P.n420 0.012
R927 OUT_P.n416 OUT_P.n415 0.012
R928 OUT_P.n398 OUT_P.n395 0.012
R929 OUT_P.n390 OUT_P.n389 0.012
R930 OUT_P.n858 OUT_P.n857 0.012
R931 OUT_P.n855 OUT_P.n854 0.012
R932 OUT_P.n893 OUT_P.n892 0.012
R933 OUT_P.n892 OUT_P.n891 0.012
R934 OUT_P.n891 OUT_P.n890 0.012
R935 OUT_P.n890 OUT_P.n889 0.012
R936 OUT_P.n960 OUT_P.n959 0.012
R937 OUT_P.n957 OUT_P.n956 0.012
R938 OUT_P.n994 OUT_P.n993 0.012
R939 OUT_P.n993 OUT_P.n992 0.012
R940 OUT_P.n992 OUT_P.n991 0.012
R941 OUT_P.n991 OUT_P.n990 0.012
R942 OUT_P.n1061 OUT_P.n1060 0.012
R943 OUT_P.n1058 OUT_P.n1057 0.012
R944 OUT_P.n1095 OUT_P.n1094 0.012
R945 OUT_P.n1094 OUT_P.n1093 0.012
R946 OUT_P.n1093 OUT_P.n1092 0.012
R947 OUT_P.n1092 OUT_P.n1091 0.012
R948 OUT_P.n578 OUT_P.n576 0.012
R949 OUT_P.n553 OUT_P.n552 0.012
R950 OUT_P.n739 OUT_P.n738 0.012
R951 OUT_P.n803 OUT_P.n797 0.012
R952 OUT_P.n624 OUT_P.n622 0.012
R953 OUT_P.n599 OUT_P.n598 0.012
R954 OUT_P.n1260 OUT_P.n1259 0.011
R955 OUT_P.n25 OUT_P.n24 0.011
R956 OUT_P.n106 OUT_P.n105 0.011
R957 OUT_P.n130 OUT_P.n129 0.011
R958 OUT_P.n160 OUT_P.n159 0.011
R959 OUT_P.n235 OUT_P.n234 0.011
R960 OUT_P.n265 OUT_P.n264 0.011
R961 OUT_P.n340 OUT_P.n339 0.011
R962 OUT_P.n370 OUT_P.n369 0.011
R963 OUT_P.n643 OUT_P.n642 0.011
R964 OUT_P.n702 OUT_P.n701 0.011
R965 OUT_P.n665 OUT_P.n664 0.011
R966 OUT_P.n706 OUT_P.n705 0.011
R967 OUT_P.n704 OUT_P.n703 0.011
R968 OUT_P.n730 OUT_P.n729 0.011
R969 OUT_P.n728 OUT_P.n727 0.011
R970 OUT_P.n736 OUT_P.n735 0.011
R971 OUT_P.n758 OUT_P.n757 0.011
R972 OUT_P.n756 OUT_P.n755 0.011
R973 OUT_P.n805 OUT_P.n804 0.011
R974 OUT_P.n771 OUT_P.n770 0.011
R975 OUT_P.n1259 OUT_P.n1258 0.011
R976 OUT_P.n1132 OUT_P.n1131 0.011
R977 OUT_P.n1273 OUT_P.n1272 0.011
R978 OUT_P.n1199 OUT_P.n1198 0.011
R979 OUT_P.n1301 OUT_P.n1300 0.011
R980 OUT_P.n1162 OUT_P.n1161 0.011
R981 OUT_P.n1238 OUT_P.n1237 0.011
R982 OUT_P.n1335 OUT_P.n1334 0.011
R983 OUT_P.n27 OUT_P.n26 0.01
R984 OUT_P.n97 OUT_P.n96 0.01
R985 OUT_P.n95 OUT_P.n94 0.01
R986 OUT_P.n93 OUT_P.n92 0.01
R987 OUT_P.n91 OUT_P.n90 0.01
R988 OUT_P.n132 OUT_P.n131 0.01
R989 OUT_P.n151 OUT_P.n150 0.01
R990 OUT_P.n149 OUT_P.n148 0.01
R991 OUT_P.n147 OUT_P.n146 0.01
R992 OUT_P.n145 OUT_P.n144 0.01
R993 OUT_P.n237 OUT_P.n236 0.01
R994 OUT_P.n256 OUT_P.n255 0.01
R995 OUT_P.n254 OUT_P.n253 0.01
R996 OUT_P.n252 OUT_P.n251 0.01
R997 OUT_P.n250 OUT_P.n249 0.01
R998 OUT_P.n342 OUT_P.n341 0.01
R999 OUT_P.n361 OUT_P.n360 0.01
R1000 OUT_P.n359 OUT_P.n358 0.01
R1001 OUT_P.n357 OUT_P.n356 0.01
R1002 OUT_P.n355 OUT_P.n354 0.01
R1003 OUT_P.n678 OUT_P.n677 0.01
R1004 OUT_P.n673 OUT_P.n671 0.01
R1005 OUT_P.n894 OUT_P.n893 0.01
R1006 OUT_P.n995 OUT_P.n994 0.01
R1007 OUT_P.n1096 OUT_P.n1095 0.01
R1008 OUT_P.n1110 OUT_P.n1109 0.01
R1009 OUT_P.n443 OUT_P.n442 0.01
R1010 OUT_P.n438 OUT_P.n436 0.01
R1011 OUT_P.n524 OUT_P.n523 0.01
R1012 OUT_P.n519 OUT_P.n517 0.01
R1013 OUT_P.n719 OUT_P.n718 0.01
R1014 OUT_P.n747 OUT_P.n746 0.01
R1015 OUT_P.n656 OUT_P.n655 0.01
R1016 OUT_P.n878 OUT_P.n877 0.009
R1017 OUT_P.n979 OUT_P.n978 0.009
R1018 OUT_P.n1080 OUT_P.n1079 0.009
R1019 OUT_P.n82 OUT_P.n80 0.009
R1020 OUT_P.n78 OUT_P.n77 0.009
R1021 OUT_P.n49 OUT_P.n47 0.009
R1022 OUT_P.n24 OUT_P.n23 0.009
R1023 OUT_P.n204 OUT_P.n202 0.009
R1024 OUT_P.n200 OUT_P.n198 0.009
R1025 OUT_P.n171 OUT_P.n170 0.009
R1026 OUT_P.n129 OUT_P.n128 0.009
R1027 OUT_P.n309 OUT_P.n307 0.009
R1028 OUT_P.n305 OUT_P.n303 0.009
R1029 OUT_P.n276 OUT_P.n275 0.009
R1030 OUT_P.n234 OUT_P.n233 0.009
R1031 OUT_P.n414 OUT_P.n412 0.009
R1032 OUT_P.n410 OUT_P.n408 0.009
R1033 OUT_P.n381 OUT_P.n380 0.009
R1034 OUT_P.n339 OUT_P.n338 0.009
R1035 OUT_P.n844 OUT_P.n841 0.009
R1036 OUT_P.n840 OUT_P.n838 0.009
R1037 OUT_P.n889 OUT_P.n888 0.009
R1038 OUT_P.n946 OUT_P.n943 0.009
R1039 OUT_P.n941 OUT_P.n939 0.009
R1040 OUT_P.n990 OUT_P.n989 0.009
R1041 OUT_P.n1047 OUT_P.n1044 0.009
R1042 OUT_P.n1042 OUT_P.n1040 0.009
R1043 OUT_P.n1091 OUT_P.n1090 0.009
R1044 OUT_P.n1110 OUT_P.n806 0.009
R1045 OUT_P.n1284 OUT_P.n1283 0.009
R1046 OUT_P.n1312 OUT_P.n1311 0.009
R1047 OUT_P.n663 OUT_P.n662 0.009
R1048 OUT_P.n726 OUT_P.n725 0.009
R1049 OUT_P.n734 OUT_P.n733 0.009
R1050 OUT_P.n732 OUT_P.n731 0.009
R1051 OUT_P.n754 OUT_P.n753 0.009
R1052 OUT_P.n769 OUT_P.n768 0.009
R1053 OUT_P.n767 OUT_P.n759 0.009
R1054 OUT_P.n1322 OUT_P.n10 0.009
R1055 OUT_P.n103 OUT_P.n102 0.008
R1056 OUT_P.n99 OUT_P.n98 0.008
R1057 OUT_P.n157 OUT_P.n156 0.008
R1058 OUT_P.n153 OUT_P.n152 0.008
R1059 OUT_P.n262 OUT_P.n261 0.008
R1060 OUT_P.n258 OUT_P.n257 0.008
R1061 OUT_P.n367 OUT_P.n366 0.008
R1062 OUT_P.n363 OUT_P.n362 0.008
R1063 OUT_P.n680 OUT_P.n679 0.008
R1064 OUT_P.n645 OUT_P.n644 0.008
R1065 OUT_P.n787 OUT_P.n786 0.008
R1066 OUT_P.n774 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE 0.008
R1067 OUT_P.n901 OUT_P.n886 0.008
R1068 OUT_P.n900 OUT_P.n899 0.008
R1069 OUT_P.n897 OUT_P.n896 0.008
R1070 OUT_P.n1002 OUT_P.n987 0.008
R1071 OUT_P.n1001 OUT_P.n1000 0.008
R1072 OUT_P.n998 OUT_P.n997 0.008
R1073 OUT_P.n1103 OUT_P.n1088 0.008
R1074 OUT_P.n1102 OUT_P.n1101 0.008
R1075 OUT_P.n1099 OUT_P.n1098 0.008
R1076 OUT_P.n1291 OUT_P.n1288 0.008
R1077 OUT_P.n445 OUT_P.n444 0.008
R1078 OUT_P.n505 OUT_P.n504 0.008
R1079 OUT_P.n492 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/GATE 0.008
R1080 OUT_P.n1319 OUT_P.n1316 0.008
R1081 OUT_P.n526 OUT_P.n525 0.008
R1082 OUT_P.n587 OUT_P.n586 0.008
R1083 OUT_P.n575 OUT_P.n574 0.008
R1084 OUT_P.n708 OUT_P.n707 0.008
R1085 OUT_P.n560 OUT_P.n559 0.008
R1086 OUT_P.n722 OUT_P.n721 0.008
R1087 OUT_P.n477 OUT_P.n476 0.008
R1088 OUT_P.n750 OUT_P.n749 0.008
R1089 OUT_P.n761 OUT_P.n760 0.008
R1090 OUT_P.n633 OUT_P.n632 0.008
R1091 OUT_P.n621 OUT_P.n620 0.008
R1092 OUT_P.n606 OUT_P.n605 0.008
R1093 OUT_P.n659 OUT_P.n658 0.008
R1094 OUT_P.n6 OUT_P.n5 0.008
R1095 OUT_P.n1111 OUT_P.n1110 0.008
R1096 OUT_P.n109 OUT_P.n108 0.007
R1097 OUT_P.n214 OUT_P.n213 0.007
R1098 OUT_P.n319 OUT_P.n318 0.007
R1099 OUT_P.n424 OUT_P.n423 0.007
R1100 OUT_P.n1104 OUT_P.n1008 0.007
R1101 OUT_P.n1003 OUT_P.n907 0.007
R1102 OUT_P.n432 OUT_P.n431 0.007
R1103 OUT_P.n1264 OUT_P.n1263 0.007
R1104 OUT_P.n426 OUT_P.n326 0.007
R1105 OUT_P.n321 OUT_P.n221 0.007
R1106 OUT_P.n216 OUT_P.n116 0.007
R1107 OUT_P.n33 OUT_P.n32 0.007
R1108 OUT_P.n50 OUT_P.n49 0.007
R1109 OUT_P.n138 OUT_P.n137 0.007
R1110 OUT_P.n172 OUT_P.n171 0.007
R1111 OUT_P.n243 OUT_P.n242 0.007
R1112 OUT_P.n277 OUT_P.n276 0.007
R1113 OUT_P.n348 OUT_P.n347 0.007
R1114 OUT_P.n382 OUT_P.n381 0.007
R1115 OUT_P.n682 OUT_P.n681 0.007
R1116 OUT_P.n791 OUT_P.n790 0.007
R1117 OUT_P.n785 OUT_P.n784 0.007
R1118 OUT_P.n868 OUT_P.n867 0.007
R1119 OUT_P.n860 OUT_P.n858 0.007
R1120 OUT_P.n883 OUT_P.n882 0.007
R1121 OUT_P.n885 OUT_P.n884 0.007
R1122 OUT_P.n970 OUT_P.n969 0.007
R1123 OUT_P.n962 OUT_P.n960 0.007
R1124 OUT_P.n984 OUT_P.n983 0.007
R1125 OUT_P.n986 OUT_P.n985 0.007
R1126 OUT_P.n1071 OUT_P.n1070 0.007
R1127 OUT_P.n1063 OUT_P.n1061 0.007
R1128 OUT_P.n1085 OUT_P.n1084 0.007
R1129 OUT_P.n1087 OUT_P.n1086 0.007
R1130 OUT_P.n447 OUT_P.n446 0.007
R1131 OUT_P.n1218 OUT_P.n1212 0.007
R1132 OUT_P.n1190 OUT_P.n1189 0.007
R1133 OUT_P.n509 OUT_P.n508 0.007
R1134 OUT_P.n503 OUT_P.n502 0.007
R1135 OUT_P.n528 OUT_P.n527 0.007
R1136 OUT_P.n1181 OUT_P.n1175 0.007
R1137 OUT_P.n1153 OUT_P.n1152 0.007
R1138 OUT_P.n564 OUT_P.n563 0.007
R1139 OUT_P.n591 OUT_P.n590 0.007
R1140 OUT_P.n585 OUT_P.n584 0.007
R1141 OUT_P.n714 OUT_P.n713 0.007
R1142 OUT_P.n711 OUT_P.n710 0.007
R1143 OUT_P.n562 OUT_P.n561 0.007
R1144 OUT_P.n556 OUT_P.n555 0.007
R1145 OUT_P.n554 OUT_P.n553 0.007
R1146 OUT_P.n548 OUT_P.n547 0.007
R1147 OUT_P.n550 OUT_P.n549 0.007
R1148 OUT_P.n738 OUT_P.n513 0.007
R1149 OUT_P.n479 OUT_P.n478 0.007
R1150 OUT_P.n473 OUT_P.n472 0.007
R1151 OUT_P.n467 OUT_P.n466 0.007
R1152 OUT_P.n469 OUT_P.n468 0.007
R1153 OUT_P.n803 OUT_P.n802 0.007
R1154 OUT_P.n799 OUT_P.n798 0.007
R1155 OUT_P.n765 OUT_P.n764 0.007
R1156 OUT_P.n1255 OUT_P.n1249 0.007
R1157 OUT_P.n1227 OUT_P.n1226 0.007
R1158 OUT_P.n1144 OUT_P.n1143 0.007
R1159 OUT_P.n610 OUT_P.n609 0.007
R1160 OUT_P.n637 OUT_P.n636 0.007
R1161 OUT_P.n631 OUT_P.n630 0.007
R1162 OUT_P.n651 OUT_P.n650 0.007
R1163 OUT_P.n648 OUT_P.n647 0.007
R1164 OUT_P.n608 OUT_P.n607 0.007
R1165 OUT_P.n602 OUT_P.n601 0.007
R1166 OUT_P.n600 OUT_P.n599 0.007
R1167 OUT_P.n700 OUT_P.n699 0.007
R1168 OUT_P.n596 OUT_P.n595 0.007
R1169 OUT_P.n1122 OUT_P.n1114 0.006
R1170 OUT_P.n102 OUT_P.n101 0.006
R1171 OUT_P.n100 OUT_P.n99 0.006
R1172 OUT_P.n156 OUT_P.n155 0.006
R1173 OUT_P.n154 OUT_P.n153 0.006
R1174 OUT_P.n261 OUT_P.n260 0.006
R1175 OUT_P.n259 OUT_P.n258 0.006
R1176 OUT_P.n366 OUT_P.n365 0.006
R1177 OUT_P.n364 OUT_P.n363 0.006
R1178 OUT_P.n646 OUT_P.n645 0.006
R1179 OUT_P.n882 OUT_P.n881 0.006
R1180 OUT_P.n886 OUT_P.n885 0.006
R1181 OUT_P.n901 OUT_P.n900 0.006
R1182 OUT_P.n898 OUT_P.n897 0.006
R1183 OUT_P.n983 OUT_P.n982 0.006
R1184 OUT_P.n987 OUT_P.n986 0.006
R1185 OUT_P.n1002 OUT_P.n1001 0.006
R1186 OUT_P.n999 OUT_P.n998 0.006
R1187 OUT_P.n1084 OUT_P.n1083 0.006
R1188 OUT_P.n1088 OUT_P.n1087 0.006
R1189 OUT_P.n1103 OUT_P.n1102 0.006
R1190 OUT_P.n1100 OUT_P.n1099 0.006
R1191 OUT_P.n709 OUT_P.n708 0.006
R1192 OUT_P.n670 OUT_P.n669 0.005
R1193 OUT_P.n668 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE 0.005
R1194 OUT_P.n435 OUT_P.n434 0.005
R1195 OUT_P.n433 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/GATE 0.005
R1196 OUT_P.n516 OUT_P.n515 0.005
R1197 OUT_P.n514 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/GATE 0.005
R1198 OUT_P.n662 OUT_P.n661 0.005
R1199 OUT_P.n725 OUT_P.n724 0.005
R1200 OUT_P.n733 OUT_P.n732 0.005
R1201 OUT_P.n753 OUT_P.n752 0.005
R1202 OUT_P.n768 OUT_P.n767 0.005
R1203 OUT_P.n42 OUT_P.n40 0.004
R1204 OUT_P.n88 OUT_P.n87 0.004
R1205 OUT_P.n110 OUT_P.n38 0.004
R1206 OUT_P.n110 OUT_P.n109 0.004
R1207 OUT_P.n90 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN 0.004
R1208 OUT_P.n164 OUT_P.n162 0.004
R1209 OUT_P.n210 OUT_P.n209 0.004
R1210 OUT_P.n215 OUT_P.n143 0.004
R1211 OUT_P.n215 OUT_P.n214 0.004
R1212 OUT_P.n144 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/DRAIN 0.004
R1213 OUT_P.n269 OUT_P.n267 0.004
R1214 OUT_P.n315 OUT_P.n314 0.004
R1215 OUT_P.n320 OUT_P.n248 0.004
R1216 OUT_P.n320 OUT_P.n319 0.004
R1217 OUT_P.n249 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/DRAIN 0.004
R1218 OUT_P.n374 OUT_P.n372 0.004
R1219 OUT_P.n420 OUT_P.n419 0.004
R1220 OUT_P.n425 OUT_P.n353 0.004
R1221 OUT_P.n425 OUT_P.n424 0.004
R1222 OUT_P.n354 OUT_P 0.004
R1223 OUT_P.n834 OUT_P.n831 0.004
R1224 OUT_P.n829 OUT_P.n827 0.004
R1225 OUT_P.n888 OUT_P.n887 0.004
R1226 OUT_P.n935 OUT_P.n932 0.004
R1227 OUT_P.n931 OUT_P.n929 0.004
R1228 OUT_P.n989 OUT_P.n988 0.004
R1229 OUT_P.n1036 OUT_P.n1033 0.004
R1230 OUT_P.n1032 OUT_P.n1030 0.004
R1231 OUT_P.n1090 OUT_P.n1089 0.004
R1232 OUT_P.n496 OUT_P.n494 0.004
R1233 OUT_P.n778 OUT_P.n776 0.004
R1234 OUT_P.n1107 OUT_P.n1106 0.003
R1235 OUT_P.n1006 OUT_P.n1005 0.003
R1236 OUT_P.n905 OUT_P.n904 0.003
R1237 OUT_P.n1106 OUT_P.n1105 0.003
R1238 OUT_P.n1005 OUT_P.n1004 0.003
R1239 OUT_P.n904 OUT_P.n903 0.003
R1240 OUT_P.n429 OUT_P.n428 0.003
R1241 OUT_P.n324 OUT_P.n323 0.003
R1242 OUT_P.n219 OUT_P.n218 0.003
R1243 OUT_P.n114 OUT_P.n113 0.003
R1244 OUT_P.n428 OUT_P.n427 0.003
R1245 OUT_P.n323 OUT_P.n322 0.003
R1246 OUT_P.n218 OUT_P.n217 0.003
R1247 OUT_P.n113 OUT_P.n112 0.003
R1248 OUT_P.n874 OUT_P.n872 0.003
R1249 OUT_P.n975 OUT_P.n973 0.003
R1250 OUT_P.n1076 OUT_P.n1074 0.003
R1251 OUT_P.n38 OUT_P.n27 0.003
R1252 OUT_P.n143 OUT_P.n132 0.003
R1253 OUT_P.n248 OUT_P.n237 0.003
R1254 OUT_P.n353 OUT_P.n342 0.003
R1255 OUT_P.n687 OUT_P.n686 0.003
R1256 OUT_P.n686 OUT_P.n685 0.003
R1257 OUT_P.n677 OUT_P.n673 0.003
R1258 OUT_P.n1134 OUT_P.n1133 0.003
R1259 OUT_P.n1133 OUT_P.n1132 0.003
R1260 OUT_P.n792 OUT_P.n791 0.003
R1261 OUT_P.n782 OUT_P.n778 0.003
R1262 OUT_P.n895 OUT_P.n894 0.003
R1263 OUT_P.n996 OUT_P.n995 0.003
R1264 OUT_P.n1097 OUT_P.n1096 0.003
R1265 OUT_P.n1291 OUT_P.n1290 0.003
R1266 OUT_P.n1274 OUT_P.n1273 0.003
R1267 OUT_P.n452 OUT_P.n451 0.003
R1268 OUT_P.n451 OUT_P.n450 0.003
R1269 OUT_P.n442 OUT_P.n438 0.003
R1270 OUT_P.n1189 OUT_P.n1188 0.003
R1271 OUT_P.n1188 OUT_P.n1187 0.003
R1272 OUT_P.n1201 OUT_P.n1200 0.003
R1273 OUT_P.n1200 OUT_P.n1199 0.003
R1274 OUT_P.n485 OUT_P.n483 0.003
R1275 OUT_P.n489 OUT_P.n485 0.003
R1276 OUT_P.n510 OUT_P.n509 0.003
R1277 OUT_P.n500 OUT_P.n496 0.003
R1278 OUT_P.n1319 OUT_P.n1318 0.003
R1279 OUT_P.n1302 OUT_P.n1301 0.003
R1280 OUT_P.n533 OUT_P.n532 0.003
R1281 OUT_P.n532 OUT_P.n531 0.003
R1282 OUT_P.n523 OUT_P.n519 0.003
R1283 OUT_P.n1152 OUT_P.n1151 0.003
R1284 OUT_P.n1151 OUT_P.n1150 0.003
R1285 OUT_P.n1164 OUT_P.n1163 0.003
R1286 OUT_P.n1163 OUT_P.n1162 0.003
R1287 OUT_P.n570 OUT_P.n566 0.003
R1288 OUT_P.n571 OUT_P.n570 0.003
R1289 OUT_P.n583 OUT_P.n582 0.003
R1290 OUT_P.n582 OUT_P.n578 0.003
R1291 OUT_P.n558 OUT_P.n557 0.003
R1292 OUT_P.n544 OUT_P.n543 0.003
R1293 OUT_P.n543 OUT_P.n542 0.003
R1294 OUT_P.n742 OUT_P.n741 0.003
R1295 OUT_P.n480 OUT_P.n479 0.003
R1296 OUT_P.n463 OUT_P.n462 0.003
R1297 OUT_P.n462 OUT_P.n461 0.003
R1298 OUT_P.n800 OUT_P.n799 0.003
R1299 OUT_P.n1240 OUT_P.n1239 0.003
R1300 OUT_P.n1239 OUT_P.n1238 0.003
R1301 OUT_P.n1226 OUT_P.n1225 0.003
R1302 OUT_P.n1225 OUT_P.n1224 0.003
R1303 OUT_P.n1114 OUT_P.n1113 0.003
R1304 OUT_P.n1113 OUT_P.n1112 0.003
R1305 OUT_P.n616 OUT_P.n612 0.003
R1306 OUT_P.n617 OUT_P.n616 0.003
R1307 OUT_P.n629 OUT_P.n628 0.003
R1308 OUT_P.n628 OUT_P.n624 0.003
R1309 OUT_P.n604 OUT_P.n603 0.003
R1310 OUT_P.n696 OUT_P.n695 0.003
R1311 OUT_P.n695 OUT_P.n694 0.003
R1312 OUT_P.n1334 OUT_P.n1333 0.003
R1313 OUT_P.n5 OUT_P.n4 0.003
R1314 OUT_P.n108 OUT_P.n107 0.002
R1315 OUT_P.n213 OUT_P.n212 0.002
R1316 OUT_P.n318 OUT_P.n317 0.002
R1317 OUT_P.n423 OUT_P.n422 0.002
R1318 OUT_P.n877 OUT_P.n876 0.002
R1319 OUT_P.n881 OUT_P.n880 0.002
R1320 OUT_P.n978 OUT_P.n977 0.002
R1321 OUT_P.n982 OUT_P.n981 0.002
R1322 OUT_P.n1079 OUT_P.n1078 0.002
R1323 OUT_P.n1083 OUT_P.n1082 0.002
R1324 OUT_P.n1082 OUT_P.n1081 0.002
R1325 OUT_P.n981 OUT_P.n980 0.002
R1326 OUT_P.n880 OUT_P.n879 0.002
R1327 OUT_P.n57 OUT_P.n56 0.002
R1328 OUT_P.n107 OUT_P.n106 0.002
R1329 OUT_P.n105 OUT_P.n104 0.002
R1330 OUT_P.n96 OUT_P.n95 0.002
R1331 OUT_P.n179 OUT_P.n178 0.002
R1332 OUT_P.n212 OUT_P.n160 0.002
R1333 OUT_P.n159 OUT_P.n158 0.002
R1334 OUT_P.n150 OUT_P.n149 0.002
R1335 OUT_P.n284 OUT_P.n283 0.002
R1336 OUT_P.n317 OUT_P.n265 0.002
R1337 OUT_P.n264 OUT_P.n263 0.002
R1338 OUT_P.n255 OUT_P.n254 0.002
R1339 OUT_P.n389 OUT_P.n388 0.002
R1340 OUT_P.n422 OUT_P.n370 0.002
R1341 OUT_P.n369 OUT_P.n368 0.002
R1342 OUT_P.n360 OUT_P.n359 0.002
R1343 OUT_P.n884 OUT_P.n883 0.002
R1344 OUT_P.n985 OUT_P.n984 0.002
R1345 OUT_P.n1086 OUT_P.n1085 0.002
R1346 OUT_P.n701 OUT_P.n665 0.002
R1347 OUT_P.n729 OUT_P.n728 0.002
R1348 OUT_P.n737 OUT_P.n736 0.002
R1349 OUT_P.n757 OUT_P.n756 0.002
R1350 OUT_P.n804 OUT_P.n771 0.002
R1351 OUT_P.n1257 OUT_P.n1256 0.002
R1352 OUT_P.n1228 OUT_P.n1221 0.002
R1353 OUT_P.n1220 OUT_P.n1219 0.002
R1354 OUT_P.n1191 OUT_P.n1184 0.002
R1355 OUT_P.n1183 OUT_P.n1182 0.002
R1356 OUT_P.n1154 OUT_P.n1147 0.002
R1357 OUT_P.n1146 OUT_P.n1145 0.002
R1358 OUT_P.n13 OUT_P.n12 0.002
R1359 OUT_P.n118 OUT_P.n117 0.002
R1360 OUT_P.n223 OUT_P.n222 0.002
R1361 OUT_P.n328 OUT_P.n327 0.002
R1362 OUT_P.n23 OUT_P.n13 0.001
R1363 OUT_P.n26 OUT_P.n25 0.001
R1364 OUT_P.n92 OUT_P.n91 0.001
R1365 OUT_P.n128 OUT_P.n118 0.001
R1366 OUT_P.n131 OUT_P.n130 0.001
R1367 OUT_P.n146 OUT_P.n145 0.001
R1368 OUT_P.n233 OUT_P.n223 0.001
R1369 OUT_P.n236 OUT_P.n235 0.001
R1370 OUT_P.n251 OUT_P.n250 0.001
R1371 OUT_P.n338 OUT_P.n328 0.001
R1372 OUT_P.n341 OUT_P.n340 0.001
R1373 OUT_P.n356 OUT_P.n355 0.001
R1374 OUT_P.n689 OUT_P.n688 0.001
R1375 OUT_P.n642 OUT_P.n641 0.001
R1376 OUT_P.n876 OUT_P.n875 0.001
R1377 OUT_P.n879 OUT_P.n878 0.001
R1378 OUT_P.n977 OUT_P.n976 0.001
R1379 OUT_P.n980 OUT_P.n979 0.001
R1380 OUT_P.n1078 OUT_P.n1077 0.001
R1381 OUT_P.n1081 OUT_P.n1080 0.001
R1382 OUT_P.n1290 OUT_P.n1289 0.001
R1383 OUT_P.n454 OUT_P.n453 0.001
R1384 OUT_P.n482 OUT_P.n481 0.001
R1385 OUT_P.n1318 OUT_P.n1317 0.001
R1386 OUT_P.n535 OUT_P.n534 0.001
R1387 OUT_P.n705 OUT_P.n704 0.001
R1388 OUT_P.n546 OUT_P.n545 0.001
R1389 OUT_P.n465 OUT_P.n464 0.001
R1390 OUT_P.n698 OUT_P.n697 0.001
R1391 OUT_P.n4 OUT_P.n3 0.001
R1392 GND.n658 GND.t17 846.712
R1393 GND.n652 GND.t34 846.712
R1394 GND.n6125 GND.t29 846.712
R1395 GND.n6132 GND.t25 846.712
R1396 GND.n3800 GND.t39 846.712
R1397 GND.n3788 GND.t13 846.712
R1398 GND.n4301 GND.t21 846.712
R1399 GND.n2418 GND.t8 846.712
R1400 GND.n2728 GND.t9 638.041
R1401 GND.n4133 GND.t22 638.041
R1402 GND.n4133 GND.t70 638.041
R1403 GND.n3202 GND.t60 638.041
R1404 GND.n3202 GND.t88 638.041
R1405 GND.n1828 GND.t4 638.041
R1406 GND.n1828 GND.t52 638.041
R1407 GND.n1844 GND.t64 638.041
R1408 GND.n1844 GND.t82 638.041
R1409 GND.n5154 GND.t44 638.041
R1410 GND.n5154 GND.t68 638.041
R1411 GND.n4403 GND.t74 638.041
R1412 GND.n4403 GND.t46 638.041
R1413 GND.n4775 GND.t0 638.041
R1414 GND.n4775 GND.t62 638.041
R1415 GND.n1300 GND.t66 638.041
R1416 GND.n1300 GND.t35 638.041
R1417 GND.n667 GND.t18 638.041
R1418 GND.n3034 GND.t40 638.041
R1419 GND.n3611 GND.t14 638.041
R1420 GND.n3611 GND.t86 638.041
R1421 GND.n3574 GND.t78 638.041
R1422 GND.n3574 GND.t56 638.041
R1423 GND.n5867 GND.t76 638.041
R1424 GND.n5867 GND.t90 638.041
R1425 GND.n1813 GND.t48 638.041
R1426 GND.n1813 GND.t54 638.041
R1427 GND.n1800 GND.t58 638.041
R1428 GND.n1800 GND.t80 638.041
R1429 GND.n1787 GND.t84 638.041
R1430 GND.n1787 GND.t72 638.041
R1431 GND.n1774 GND.t50 638.041
R1432 GND.n1774 GND.t6 638.041
R1433 GND.n1611 GND.t2 638.041
R1434 GND.n1611 GND.t30 638.041
R1435 GND.n1093 GND.t26 638.041
R1436 GND.n5972 GND.n5971 135.862
R1437 GND.n4750 GND.n4749 135.862
R1438 GND.n5952 GND.n5951 115.482
R1439 GND.n4767 GND.n4766 115.482
R1440 GND.n5934 GND.n5933 95.103
R1441 GND.n5128 GND.n5127 95.103
R1442 GND.n5916 GND.n5915 74.724
R1443 GND.n5146 GND.n5145 74.724
R1444 GND.n4668 GND.n4667 55.353
R1445 GND.n3485 GND.n3484 55.353
R1446 GND.n1690 GND.n1689 54.344
R1447 GND.n1374 GND.n1373 54.344
R1448 GND.n5792 GND.n5791 54.344
R1449 GND.n5612 GND.n5611 54.344
R1450 GND.n1918 GND.n1917 54.344
R1451 GND.n2098 GND.n2097 54.344
R1452 GND.n5228 GND.n5227 54.344
R1453 GND.n5408 GND.n5407 54.344
R1454 GND.n4478 GND.n4477 54.344
R1455 GND.n4660 GND.n4659 54.344
R1456 GND.n4669 GND.n4668 54.344
R1457 GND.n4849 GND.n4848 54.344
R1458 GND.n5029 GND.n5028 54.344
R1459 GND.n3494 GND.n3493 54.344
R1460 GND.n3486 GND.n3485 54.344
R1461 GND.n3310 GND.n3309 54.344
R1462 GND.n3703 GND.n3702 54.344
R1463 GND.n4207 GND.n4206 54.344
R1464 GND.n5898 GND.n5897 54.344
R1465 GND.n1185 GND.n1184 54.344
R1466 GND.n740 GND.n739 54.344
R1467 GND.n5508 GND.n5507 54.344
R1468 GND.n3113 GND.n3112 54.344
R1469 GND.n2802 GND.n2801 54.344
R1470 GND.n1702 GND.n1701 47.551
R1471 GND.n1362 GND.n1361 47.551
R1472 GND.n5804 GND.n5803 47.551
R1473 GND.n5624 GND.n5623 47.551
R1474 GND.n1906 GND.n1905 47.551
R1475 GND.n2086 GND.n2085 47.551
R1476 GND.n5216 GND.n5215 47.551
R1477 GND.n5396 GND.n5395 47.551
R1478 GND.n4466 GND.n4465 47.551
R1479 GND.n4837 GND.n4836 47.551
R1480 GND.n5017 GND.n5016 47.551
R1481 GND.n3322 GND.n3321 47.551
R1482 GND.n3715 GND.n3714 47.551
R1483 GND.n4195 GND.n4194 47.551
R1484 GND.n1197 GND.n1196 47.551
R1485 GND.n728 GND.n727 47.551
R1486 GND.n3125 GND.n3124 47.551
R1487 GND.n2790 GND.n2789 47.551
R1488 GND.n6319 GND.n6317 46.305
R1489 GND.n1612 GND.n1610 44.155
R1490 GND.n5714 GND.n5713 44.155
R1491 GND.n2000 GND.n1999 44.155
R1492 GND.n1845 GND.n1843 44.155
R1493 GND.n5310 GND.n5309 44.155
R1494 GND.n5155 GND.n5153 44.155
R1495 GND.n4560 GND.n4559 44.155
R1496 GND.n4931 GND.n4930 44.155
R1497 GND.n4776 GND.n4774 44.155
R1498 GND.n3625 GND.n3624 44.155
R1499 GND.n4289 GND.n4288 44.155
R1500 GND.n1107 GND.n1106 44.155
R1501 GND.n668 GND.n666 44.155
R1502 GND.n3035 GND.n3033 44.155
R1503 GND.n2884 GND.n2883 44.155
R1504 GND.n1714 GND.n1713 40.758
R1505 GND.n1350 GND.n1349 40.758
R1506 GND.n5816 GND.n5815 40.758
R1507 GND.n5636 GND.n5635 40.758
R1508 GND.n1894 GND.n1893 40.758
R1509 GND.n2074 GND.n2073 40.758
R1510 GND.n5204 GND.n5203 40.758
R1511 GND.n5384 GND.n5383 40.758
R1512 GND.n4454 GND.n4453 40.758
R1513 GND.n4635 GND.n4634 40.758
R1514 GND.n4694 GND.n4693 40.758
R1515 GND.n4825 GND.n4824 40.758
R1516 GND.n5005 GND.n5004 40.758
R1517 GND.n3519 GND.n3518 40.758
R1518 GND.n3460 GND.n3459 40.758
R1519 GND.n3334 GND.n3333 40.758
R1520 GND.n3727 GND.n3726 40.758
R1521 GND.n4183 GND.n4182 40.758
R1522 GND.n1209 GND.n1208 40.758
R1523 GND.n716 GND.n715 40.758
R1524 GND.n3137 GND.n3136 40.758
R1525 GND.n2778 GND.n2777 40.758
R1526 GND.n1763 GND.n1762 40.459
R1527 GND.n1303 GND.n1302 40.459
R1528 GND.n5870 GND.n5869 40.459
R1529 GND.n5685 GND.n5684 40.459
R1530 GND.n1831 GND.n1830 40.459
R1531 GND.n1816 GND.n1815 40.459
R1532 GND.n2027 GND.n2026 40.459
R1533 GND.n1803 GND.n1802 40.459
R1534 GND.n5337 GND.n5336 40.459
R1535 GND.n1790 GND.n1789 40.459
R1536 GND.n4404 GND.n4401 40.459
R1537 GND.n4587 GND.n4586 40.459
R1538 GND.n1777 GND.n1776 40.459
R1539 GND.n4958 GND.n4957 40.459
R1540 GND.n3411 GND.n3410 40.459
R1541 GND.n3383 GND.n3382 40.459
R1542 GND.n3205 GND.n3204 40.459
R1543 GND.n3575 GND.n3573 40.459
R1544 GND.n3614 GND.n3613 40.459
R1545 GND.n4136 GND.n4135 40.459
R1546 GND.n1096 GND.n1095 40.459
R1547 GND.n6153 GND.n6152 40.459
R1548 GND.n2731 GND.n2730 40.459
R1549 GND.n3186 GND.n3185 40.459
R1550 GND.n1456 GND.n1455 40.459
R1551 GND.n1624 GND.n1623 37.362
R1552 GND.n1445 GND.n1443 37.362
R1553 GND.n5726 GND.n5725 37.362
R1554 GND.n5546 GND.n5544 37.362
R1555 GND.n1988 GND.n1987 37.362
R1556 GND.n2168 GND.n2167 37.362
R1557 GND.n5298 GND.n5297 37.362
R1558 GND.n5478 GND.n5477 37.362
R1559 GND.n4548 GND.n4547 37.362
R1560 GND.n4600 GND.n4599 37.362
R1561 GND.n4734 GND.n4732 37.362
R1562 GND.n4919 GND.n4918 37.362
R1563 GND.n5099 GND.n5098 37.362
R1564 GND.n3559 GND.n3557 37.362
R1565 GND.n3425 GND.n3423 37.362
R1566 GND.n3244 GND.n3242 37.362
R1567 GND.n3637 GND.n3636 37.362
R1568 GND.n4277 GND.n4276 37.362
R1569 GND.n1119 GND.n1118 37.362
R1570 GND.n810 GND.n809 37.362
R1571 GND.n3047 GND.n3046 37.362
R1572 GND.n2872 GND.n2871 37.362
R1573 GND.n1751 GND.n1750 34.603
R1574 GND.n1315 GND.n1314 34.603
R1575 GND.n5853 GND.n5852 34.603
R1576 GND.n5673 GND.n5672 34.603
R1577 GND.n1859 GND.n1858 34.603
R1578 GND.n2039 GND.n2038 34.603
R1579 GND.n5169 GND.n5168 34.603
R1580 GND.n5349 GND.n5348 34.603
R1581 GND.n4419 GND.n4418 34.603
R1582 GND.n4790 GND.n4789 34.603
R1583 GND.n4970 GND.n4969 34.603
R1584 GND.n3371 GND.n3370 34.603
R1585 GND.n3764 GND.n3763 34.603
R1586 GND.n4148 GND.n4147 34.603
R1587 GND.n1246 GND.n1245 34.603
R1588 GND.n681 GND.n680 34.603
R1589 GND.n3174 GND.n3173 34.603
R1590 GND.n2743 GND.n2742 34.603
R1591 GND.n1726 GND.n1725 33.965
R1592 GND.n1338 GND.n1337 33.965
R1593 GND.n5828 GND.n5827 33.965
R1594 GND.n5648 GND.n5647 33.965
R1595 GND.n1882 GND.n1881 33.965
R1596 GND.n2062 GND.n2061 33.965
R1597 GND.n5192 GND.n5191 33.965
R1598 GND.n5372 GND.n5371 33.965
R1599 GND.n4442 GND.n4441 33.965
R1600 GND.n4813 GND.n4812 33.965
R1601 GND.n4993 GND.n4992 33.965
R1602 GND.n3346 GND.n3345 33.965
R1603 GND.n3739 GND.n3738 33.965
R1604 GND.n4171 GND.n4170 33.965
R1605 GND.n5880 GND.n5879 33.965
R1606 GND.n1221 GND.n1220 33.965
R1607 GND.n704 GND.n703 33.965
R1608 GND.n5526 GND.n5525 33.965
R1609 GND.n3149 GND.n3148 33.965
R1610 GND.n2766 GND.n2765 33.965
R1611 GND.n2441 GND.n2439 33.505
R1612 GND.n1636 GND.n1635 30.568
R1613 GND.n1432 GND.n1431 30.568
R1614 GND.n5738 GND.n5737 30.568
R1615 GND.n5558 GND.n5557 30.568
R1616 GND.n1976 GND.n1975 30.568
R1617 GND.n2156 GND.n2155 30.568
R1618 GND.n5286 GND.n5285 30.568
R1619 GND.n5466 GND.n5465 30.568
R1620 GND.n4536 GND.n4535 30.568
R1621 GND.n4907 GND.n4906 30.568
R1622 GND.n5087 GND.n5086 30.568
R1623 GND.n3256 GND.n3255 30.568
R1624 GND.n3649 GND.n3648 30.568
R1625 GND.n4265 GND.n4264 30.568
R1626 GND.n1131 GND.n1130 30.568
R1627 GND.n798 GND.n797 30.568
R1628 GND.n3059 GND.n3058 30.568
R1629 GND.n2860 GND.n2859 30.568
R1630 GND.n1264 GND.n1263 30.117
R1631 GND.n1739 GND.n1738 28.618
R1632 GND.n1327 GND.n1326 28.618
R1633 GND.n5841 GND.n5840 28.618
R1634 GND.n5661 GND.n5660 28.618
R1635 GND.n1871 GND.n1870 28.618
R1636 GND.n2051 GND.n2050 28.618
R1637 GND.n5181 GND.n5180 28.618
R1638 GND.n5361 GND.n5360 28.618
R1639 GND.n4431 GND.n4430 28.618
R1640 GND.n4720 GND.n4719 28.618
R1641 GND.n4611 GND.n4610 28.618
R1642 GND.n4802 GND.n4801 28.618
R1643 GND.n4982 GND.n4981 28.618
R1644 GND.n3436 GND.n3435 28.618
R1645 GND.n3359 GND.n3358 28.618
R1646 GND.n3545 GND.n3544 28.618
R1647 GND.n3752 GND.n3751 28.618
R1648 GND.n4160 GND.n4159 28.618
R1649 GND.n1234 GND.n1233 28.618
R1650 GND.n693 GND.n692 28.618
R1651 GND.n3162 GND.n3161 28.618
R1652 GND.n2755 GND.n2754 28.618
R1653 GND.n5875 GND.n5874 28.611
R1654 GND.n5532 GND.n5531 28.611
R1655 GND.n1821 GND.n1820 28.611
R1656 GND.n2180 GND.n2178 28.611
R1657 GND.n1808 GND.n1807 28.611
R1658 GND.n5490 GND.n5488 28.611
R1659 GND.n1795 GND.n1794 28.611
R1660 GND.n4746 GND.n4744 28.611
R1661 GND.n1782 GND.n1781 28.611
R1662 GND.n5111 GND.n5109 28.611
R1663 GND.n3580 GND.n3579 28.611
R1664 GND.n3230 GND.n3229 28.611
R1665 GND.n3777 GND.n3775 28.611
R1666 GND.n1259 GND.n1257 28.611
R1667 GND.n6317 GND.n671 28.611
R1668 GND.n1738 GND.n1737 27.172
R1669 GND.n1326 GND.n1325 27.172
R1670 GND.n5840 GND.n5839 27.172
R1671 GND.n5660 GND.n5659 27.172
R1672 GND.n1870 GND.n1869 27.172
R1673 GND.n2050 GND.n2049 27.172
R1674 GND.n5180 GND.n5179 27.172
R1675 GND.n5360 GND.n5359 27.172
R1676 GND.n4430 GND.n4429 27.172
R1677 GND.n4610 GND.n4609 27.172
R1678 GND.n4719 GND.n4718 27.172
R1679 GND.n4801 GND.n4800 27.172
R1680 GND.n4981 GND.n4980 27.172
R1681 GND.n3544 GND.n3543 27.172
R1682 GND.n3435 GND.n3434 27.172
R1683 GND.n3358 GND.n3357 27.172
R1684 GND.n3751 GND.n3750 27.172
R1685 GND.n4159 GND.n4158 27.172
R1686 GND.n1233 GND.n1232 27.172
R1687 GND.n692 GND.n691 27.172
R1688 GND.n3161 GND.n3160 27.172
R1689 GND.n2754 GND.n2753 27.172
R1690 GND.n1683 GND.n1682 25.966
R1691 GND.n1383 GND.n1382 25.966
R1692 GND.n5785 GND.n5784 25.966
R1693 GND.n5605 GND.n5604 25.966
R1694 GND.n1927 GND.n1926 25.966
R1695 GND.n2107 GND.n2106 25.966
R1696 GND.n5237 GND.n5236 25.966
R1697 GND.n5417 GND.n5416 25.966
R1698 GND.n5416 GND.n5415 25.966
R1699 GND.n2106 GND.n2105 25.966
R1700 GND.n5604 GND.n5603 25.966
R1701 GND.n4487 GND.n4486 25.966
R1702 GND.n4858 GND.n4857 25.966
R1703 GND.n5038 GND.n5037 25.966
R1704 GND.n5037 GND.n5036 25.966
R1705 GND.n4857 GND.n4856 25.966
R1706 GND.n4486 GND.n4485 25.966
R1707 GND.n5236 GND.n5235 25.966
R1708 GND.n1926 GND.n1925 25.966
R1709 GND.n5784 GND.n5783 25.966
R1710 GND.n3303 GND.n3302 25.966
R1711 GND.n3302 GND.n3301 25.966
R1712 GND.n3696 GND.n3695 25.966
R1713 GND.n4216 GND.n4215 25.966
R1714 GND.n3695 GND.n3694 25.966
R1715 GND.n4215 GND.n4214 25.966
R1716 GND.n1178 GND.n1177 25.966
R1717 GND.n749 GND.n748 25.966
R1718 GND.n3106 GND.n3105 25.966
R1719 GND.n2811 GND.n2810 25.966
R1720 GND.n2810 GND.n2809 25.966
R1721 GND.n3105 GND.n3104 25.966
R1722 GND.n1177 GND.n1176 25.966
R1723 GND.n748 GND.n747 25.966
R1724 GND.n1682 GND.n1681 25.966
R1725 GND.n1382 GND.n1381 25.966
R1726 GND.n653 GND.n652 24.127
R1727 GND.n659 GND.n658 24.127
R1728 GND.n495 GND.n494 24.127
R1729 GND.n501 GND.n500 24.127
R1730 GND.n1279 GND.n1278 24.127
R1731 GND.n1269 GND.n1268 24.127
R1732 GND.n6126 GND.n6125 24.127
R1733 GND.n6133 GND.n6132 24.127
R1734 GND.n3801 GND.n3800 24.127
R1735 GND.n3789 GND.n3788 24.127
R1736 GND.n3954 GND.n3953 24.127
R1737 GND.n3961 GND.n3960 24.127
R1738 GND.n2419 GND.n2418 24.127
R1739 GND.n4302 GND.n4301 24.127
R1740 GND.n2261 GND.n2260 24.127
R1741 GND.n2267 GND.n2266 24.127
R1742 GND.n1648 GND.n1647 23.775
R1743 GND.n1420 GND.n1419 23.775
R1744 GND.n5750 GND.n5749 23.775
R1745 GND.n5570 GND.n5569 23.775
R1746 GND.n1964 GND.n1963 23.775
R1747 GND.n2144 GND.n2143 23.775
R1748 GND.n5274 GND.n5273 23.775
R1749 GND.n5454 GND.n5453 23.775
R1750 GND.n4524 GND.n4523 23.775
R1751 GND.n4625 GND.n4623 23.775
R1752 GND.n4709 GND.n4707 23.775
R1753 GND.n4895 GND.n4894 23.775
R1754 GND.n5075 GND.n5074 23.775
R1755 GND.n3534 GND.n3532 23.775
R1756 GND.n3450 GND.n3448 23.775
R1757 GND.n3268 GND.n3267 23.775
R1758 GND.n3661 GND.n3660 23.775
R1759 GND.n4253 GND.n4252 23.775
R1760 GND.n1143 GND.n1142 23.775
R1761 GND.n786 GND.n785 23.775
R1762 GND.n3071 GND.n3070 23.775
R1763 GND.n2848 GND.n2847 23.775
R1764 GND.n1671 GND.n1670 22.848
R1765 GND.n1395 GND.n1394 22.848
R1766 GND.n5773 GND.n5772 22.848
R1767 GND.n5593 GND.n5592 22.848
R1768 GND.n1939 GND.n1938 22.848
R1769 GND.n2119 GND.n2118 22.848
R1770 GND.n5249 GND.n5248 22.848
R1771 GND.n5429 GND.n5428 22.848
R1772 GND.n5428 GND.n5427 22.848
R1773 GND.n2118 GND.n2117 22.848
R1774 GND.n5592 GND.n5591 22.848
R1775 GND.n4499 GND.n4498 22.848
R1776 GND.n4648 GND.n4647 22.848
R1777 GND.n4681 GND.n4680 22.848
R1778 GND.n4682 GND.n4681 22.848
R1779 GND.n4647 GND.n4646 22.848
R1780 GND.n4870 GND.n4869 22.848
R1781 GND.n5050 GND.n5049 22.848
R1782 GND.n5049 GND.n5048 22.848
R1783 GND.n4869 GND.n4868 22.848
R1784 GND.n4498 GND.n4497 22.848
R1785 GND.n5248 GND.n5247 22.848
R1786 GND.n1938 GND.n1937 22.848
R1787 GND.n5772 GND.n5771 22.848
R1788 GND.n3507 GND.n3506 22.848
R1789 GND.n3472 GND.n3471 22.848
R1790 GND.n3291 GND.n3290 22.848
R1791 GND.n3473 GND.n3472 22.848
R1792 GND.n3506 GND.n3505 22.848
R1793 GND.n3290 GND.n3289 22.848
R1794 GND.n3684 GND.n3683 22.848
R1795 GND.n4228 GND.n4227 22.848
R1796 GND.n3683 GND.n3682 22.848
R1797 GND.n4227 GND.n4226 22.848
R1798 GND.n1166 GND.n1165 22.848
R1799 GND.n761 GND.n760 22.848
R1800 GND.n3094 GND.n3093 22.848
R1801 GND.n2823 GND.n2822 22.848
R1802 GND.n2822 GND.n2821 22.848
R1803 GND.n3093 GND.n3092 22.848
R1804 GND.n1165 GND.n1164 22.848
R1805 GND.n760 GND.n759 22.848
R1806 GND.n1670 GND.n1669 22.848
R1807 GND.n1394 GND.n1393 22.848
R1808 GND.n1727 GND.n1726 22.503
R1809 GND.n1339 GND.n1338 22.503
R1810 GND.n5829 GND.n5828 22.503
R1811 GND.n5649 GND.n5648 22.503
R1812 GND.n1883 GND.n1882 22.503
R1813 GND.n2063 GND.n2062 22.503
R1814 GND.n5193 GND.n5192 22.503
R1815 GND.n5373 GND.n5372 22.503
R1816 GND.n4443 GND.n4442 22.503
R1817 GND.n4814 GND.n4813 22.503
R1818 GND.n4994 GND.n4993 22.503
R1819 GND.n3347 GND.n3346 22.503
R1820 GND.n3740 GND.n3739 22.503
R1821 GND.n4172 GND.n4171 22.503
R1822 GND.n1222 GND.n1221 22.503
R1823 GND.n705 GND.n704 22.503
R1824 GND.n3150 GND.n3149 22.503
R1825 GND.n2767 GND.n2766 22.503
R1826 GND.n1750 GND.n1749 20.379
R1827 GND.n1314 GND.n1313 20.379
R1828 GND.n5852 GND.n5851 20.379
R1829 GND.n5672 GND.n5671 20.379
R1830 GND.n1858 GND.n1857 20.379
R1831 GND.n2038 GND.n2037 20.379
R1832 GND.n5168 GND.n5167 20.379
R1833 GND.n5348 GND.n5347 20.379
R1834 GND.n4418 GND.n4417 20.379
R1835 GND.n4789 GND.n4788 20.379
R1836 GND.n4969 GND.n4968 20.379
R1837 GND.n3370 GND.n3369 20.379
R1838 GND.n3763 GND.n3762 20.379
R1839 GND.n4147 GND.n4146 20.379
R1840 GND.n1245 GND.n1244 20.379
R1841 GND.n680 GND.n679 20.379
R1842 GND.n3173 GND.n3172 20.379
R1843 GND.n2742 GND.n2741 20.379
R1844 GND.n1659 GND.n1658 19.694
R1845 GND.n1407 GND.n1406 19.694
R1846 GND.n5761 GND.n5760 19.694
R1847 GND.n5581 GND.n5580 19.694
R1848 GND.n1951 GND.n1950 19.694
R1849 GND.n2131 GND.n2130 19.694
R1850 GND.n5261 GND.n5260 19.694
R1851 GND.n5441 GND.n5440 19.694
R1852 GND.n5440 GND.n5439 19.694
R1853 GND.n2130 GND.n2129 19.694
R1854 GND.n5580 GND.n5579 19.694
R1855 GND.n4511 GND.n4510 19.694
R1856 GND.n4882 GND.n4881 19.694
R1857 GND.n5062 GND.n5061 19.694
R1858 GND.n5061 GND.n5060 19.694
R1859 GND.n4881 GND.n4880 19.694
R1860 GND.n4510 GND.n4509 19.694
R1861 GND.n5260 GND.n5259 19.694
R1862 GND.n1950 GND.n1949 19.694
R1863 GND.n5760 GND.n5759 19.694
R1864 GND.n3279 GND.n3278 19.694
R1865 GND.n3278 GND.n3277 19.694
R1866 GND.n3672 GND.n3671 19.694
R1867 GND.n4240 GND.n4239 19.694
R1868 GND.n3671 GND.n3670 19.694
R1869 GND.n4239 GND.n4238 19.694
R1870 GND.n1154 GND.n1153 19.694
R1871 GND.n773 GND.n772 19.694
R1872 GND.n3082 GND.n3081 19.694
R1873 GND.n2835 GND.n2834 19.694
R1874 GND.n2834 GND.n2833 19.694
R1875 GND.n3081 GND.n3080 19.694
R1876 GND.n1153 GND.n1152 19.694
R1877 GND.n772 GND.n771 19.694
R1878 GND.n1658 GND.n1657 19.694
R1879 GND.n1406 GND.n1405 19.694
R1880 GND.n1660 GND.n1659 16.982
R1881 GND.n1408 GND.n1407 16.982
R1882 GND.n5762 GND.n5761 16.982
R1883 GND.n5582 GND.n5581 16.982
R1884 GND.n1952 GND.n1951 16.982
R1885 GND.n2132 GND.n2131 16.982
R1886 GND.n5262 GND.n5261 16.982
R1887 GND.n5442 GND.n5441 16.982
R1888 GND.n4512 GND.n4511 16.982
R1889 GND.n4883 GND.n4882 16.982
R1890 GND.n5063 GND.n5062 16.982
R1891 GND.n3280 GND.n3279 16.982
R1892 GND.n3673 GND.n3672 16.982
R1893 GND.n4241 GND.n4240 16.982
R1894 GND.n1155 GND.n1154 16.982
R1895 GND.n774 GND.n773 16.982
R1896 GND.n3083 GND.n3082 16.982
R1897 GND.n2836 GND.n2835 16.982
R1898 GND.n1647 GND.n1646 16.504
R1899 GND.n1419 GND.n1418 16.504
R1900 GND.n5749 GND.n5748 16.504
R1901 GND.n5569 GND.n5568 16.504
R1902 GND.n1963 GND.n1962 16.504
R1903 GND.n2143 GND.n2142 16.504
R1904 GND.n5273 GND.n5272 16.504
R1905 GND.n5453 GND.n5452 16.504
R1906 GND.n5452 GND.n5451 16.504
R1907 GND.n2142 GND.n2141 16.504
R1908 GND.n5568 GND.n5567 16.504
R1909 GND.n4523 GND.n4522 16.504
R1910 GND.n4623 GND.n4622 16.504
R1911 GND.n4706 GND.n4705 16.504
R1912 GND.n4707 GND.n4706 16.504
R1913 GND.n4622 GND.n4621 16.504
R1914 GND.n4894 GND.n4893 16.504
R1915 GND.n5074 GND.n5073 16.504
R1916 GND.n5073 GND.n5072 16.504
R1917 GND.n4893 GND.n4892 16.504
R1918 GND.n4522 GND.n4521 16.504
R1919 GND.n5272 GND.n5271 16.504
R1920 GND.n1962 GND.n1961 16.504
R1921 GND.n5748 GND.n5747 16.504
R1922 GND.n3532 GND.n3531 16.504
R1923 GND.n3447 GND.n3446 16.504
R1924 GND.n3267 GND.n3266 16.504
R1925 GND.n3448 GND.n3447 16.504
R1926 GND.n3531 GND.n3530 16.504
R1927 GND.n3266 GND.n3265 16.504
R1928 GND.n3660 GND.n3659 16.504
R1929 GND.n4252 GND.n4251 16.504
R1930 GND.n3659 GND.n3658 16.504
R1931 GND.n4251 GND.n4250 16.504
R1932 GND.n1142 GND.n1141 16.504
R1933 GND.n785 GND.n784 16.504
R1934 GND.n3070 GND.n3069 16.504
R1935 GND.n2847 GND.n2846 16.504
R1936 GND.n2846 GND.n2845 16.504
R1937 GND.n3069 GND.n3068 16.504
R1938 GND.n1141 GND.n1140 16.504
R1939 GND.n784 GND.n783 16.504
R1940 GND.n1646 GND.n1645 16.504
R1941 GND.n1418 GND.n1417 16.504
R1942 GND.n1715 GND.n1714 16.252
R1943 GND.n1351 GND.n1350 16.252
R1944 GND.n5817 GND.n5816 16.252
R1945 GND.n5637 GND.n5636 16.252
R1946 GND.n1895 GND.n1894 16.252
R1947 GND.n2075 GND.n2074 16.252
R1948 GND.n5205 GND.n5204 16.252
R1949 GND.n5385 GND.n5384 16.252
R1950 GND.n4455 GND.n4454 16.252
R1951 GND.n4695 GND.n4694 16.252
R1952 GND.n4636 GND.n4635 16.252
R1953 GND.n4826 GND.n4825 16.252
R1954 GND.n5006 GND.n5005 16.252
R1955 GND.n3461 GND.n3460 16.252
R1956 GND.n3335 GND.n3334 16.252
R1957 GND.n3520 GND.n3519 16.252
R1958 GND.n3728 GND.n3727 16.252
R1959 GND.n4184 GND.n4183 16.252
R1960 GND.n1210 GND.n1209 16.252
R1961 GND.n717 GND.n716 16.252
R1962 GND.n3138 GND.n3137 16.252
R1963 GND.n2779 GND.n2778 16.252
R1964 GND.n5973 GND.n5970 15.058
R1965 GND.n4751 GND.n4748 15.058
R1966 GND.n1762 GND.n1761 13.586
R1967 GND.n1302 GND.n1301 13.586
R1968 GND.n1455 GND.n1454 13.586
R1969 GND.n5869 GND.n5868 13.586
R1970 GND.n5684 GND.n5683 13.586
R1971 GND.n1830 GND.n1829 13.586
R1972 GND.n1815 GND.n1814 13.586
R1973 GND.n2026 GND.n2025 13.586
R1974 GND.n1802 GND.n1801 13.586
R1975 GND.n5336 GND.n5335 13.586
R1976 GND.n1789 GND.n1788 13.586
R1977 GND.n4586 GND.n4585 13.586
R1978 GND.n4401 GND.n4400 13.586
R1979 GND.n1776 GND.n1775 13.586
R1980 GND.n4957 GND.n4956 13.586
R1981 GND.n3573 GND.n3572 13.586
R1982 GND.n3410 GND.n3409 13.586
R1983 GND.n3382 GND.n3381 13.586
R1984 GND.n3204 GND.n3203 13.586
R1985 GND.n3613 GND.n3612 13.586
R1986 GND.n4135 GND.n4134 13.586
R1987 GND.n3593 GND.n3592 13.586
R1988 GND.n1095 GND.n1094 13.586
R1989 GND.n6152 GND.n6151 13.586
R1990 GND.n3224 GND.n3223 13.586
R1991 GND.n3185 GND.n3184 13.586
R1992 GND.n2730 GND.n2729 13.586
R1993 GND.n1635 GND.n1634 13.278
R1994 GND.n1431 GND.n1430 13.278
R1995 GND.n5737 GND.n5736 13.278
R1996 GND.n5557 GND.n5556 13.278
R1997 GND.n1975 GND.n1974 13.278
R1998 GND.n2155 GND.n2154 13.278
R1999 GND.n5285 GND.n5284 13.278
R2000 GND.n5465 GND.n5464 13.278
R2001 GND.n5464 GND.n5463 13.278
R2002 GND.n2154 GND.n2153 13.278
R2003 GND.n5556 GND.n5555 13.278
R2004 GND.n4535 GND.n4534 13.278
R2005 GND.n4906 GND.n4905 13.278
R2006 GND.n5086 GND.n5085 13.278
R2007 GND.n5085 GND.n5084 13.278
R2008 GND.n4905 GND.n4904 13.278
R2009 GND.n4534 GND.n4533 13.278
R2010 GND.n5284 GND.n5283 13.278
R2011 GND.n1974 GND.n1973 13.278
R2012 GND.n5736 GND.n5735 13.278
R2013 GND.n3255 GND.n3254 13.278
R2014 GND.n3254 GND.n3253 13.278
R2015 GND.n3648 GND.n3647 13.278
R2016 GND.n4264 GND.n4263 13.278
R2017 GND.n3647 GND.n3646 13.278
R2018 GND.n4263 GND.n4262 13.278
R2019 GND.n1130 GND.n1129 13.278
R2020 GND.n797 GND.n796 13.278
R2021 GND.n3058 GND.n3057 13.278
R2022 GND.n2859 GND.n2858 13.278
R2023 GND.n2858 GND.n2857 13.278
R2024 GND.n3057 GND.n3056 13.278
R2025 GND.n1129 GND.n1128 13.278
R2026 GND.n796 GND.n795 13.278
R2027 GND.n1634 GND.n1633 13.278
R2028 GND.n1430 GND.n1429 13.278
R2029 GND.n6215 GND.n6214 13.176
R2030 GND.n604 GND.n603 13.176
R2031 GND.n6074 GND.n6073 13.176
R2032 GND.n994 GND.n993 13.176
R2033 GND.n897 GND.n896 13.176
R2034 GND.n3902 GND.n3901 13.176
R2035 GND.n2616 GND.n2615 13.176
R2036 GND.n2519 GND.n2518 13.176
R2037 GND.n4072 GND.n4071 13.176
R2038 GND.n2370 GND.n2369 13.176
R2039 GND.n2961 GND.n2960 13.176
R2040 GND.n1540 GND.n1539 13.176
R2041 GND.n5953 GND.n5950 12.8
R2042 GND.n4768 GND.n4765 12.8
R2043 GND.n5935 GND.n5932 10.541
R2044 GND.n5129 GND.n5126 10.541
R2045 GND.n1672 GND.n1671 10.189
R2046 GND.n1396 GND.n1395 10.189
R2047 GND.n5774 GND.n5773 10.189
R2048 GND.n5594 GND.n5593 10.189
R2049 GND.n1940 GND.n1939 10.189
R2050 GND.n2120 GND.n2119 10.189
R2051 GND.n5250 GND.n5249 10.189
R2052 GND.n5430 GND.n5429 10.189
R2053 GND.n4500 GND.n4499 10.189
R2054 GND.n4650 GND.n4648 10.189
R2055 GND.n4684 GND.n4682 10.189
R2056 GND.n4871 GND.n4870 10.189
R2057 GND.n5051 GND.n5050 10.189
R2058 GND.n3509 GND.n3507 10.189
R2059 GND.n3475 GND.n3473 10.189
R2060 GND.n3292 GND.n3291 10.189
R2061 GND.n3685 GND.n3684 10.189
R2062 GND.n4229 GND.n4228 10.189
R2063 GND.n1167 GND.n1166 10.189
R2064 GND.n762 GND.n761 10.189
R2065 GND.n3095 GND.n3094 10.189
R2066 GND.n2824 GND.n2823 10.189
R2067 GND.n1623 GND.n1622 10.016
R2068 GND.n1443 GND.n1442 10.016
R2069 GND.n5725 GND.n5724 10.016
R2070 GND.n5544 GND.n5543 10.016
R2071 GND.n1987 GND.n1986 10.016
R2072 GND.n2167 GND.n2166 10.016
R2073 GND.n5297 GND.n5296 10.016
R2074 GND.n5477 GND.n5476 10.016
R2075 GND.n5476 GND.n5475 10.016
R2076 GND.n2166 GND.n2165 10.016
R2077 GND.n5543 GND.n5542 10.016
R2078 GND.n4547 GND.n4546 10.016
R2079 GND.n4599 GND.n4598 10.016
R2080 GND.n4731 GND.n4730 10.016
R2081 GND.n4732 GND.n4731 10.016
R2082 GND.n4598 GND.n4597 10.016
R2083 GND.n4918 GND.n4917 10.016
R2084 GND.n5098 GND.n5097 10.016
R2085 GND.n5097 GND.n5096 10.016
R2086 GND.n4917 GND.n4916 10.016
R2087 GND.n4546 GND.n4545 10.016
R2088 GND.n5296 GND.n5295 10.016
R2089 GND.n1986 GND.n1985 10.016
R2090 GND.n5724 GND.n5723 10.016
R2091 GND.n3557 GND.n3556 10.016
R2092 GND.n3422 GND.n3421 10.016
R2093 GND.n3242 GND.n3241 10.016
R2094 GND.n3423 GND.n3422 10.016
R2095 GND.n3556 GND.n3555 10.016
R2096 GND.n3241 GND.n3240 10.016
R2097 GND.n3636 GND.n3635 10.016
R2098 GND.n4276 GND.n4275 10.016
R2099 GND.n3635 GND.n3634 10.016
R2100 GND.n4275 GND.n4274 10.016
R2101 GND.n1118 GND.n1117 10.016
R2102 GND.n809 GND.n808 10.016
R2103 GND.n3046 GND.n3045 10.016
R2104 GND.n2871 GND.n2870 10.016
R2105 GND.n2870 GND.n2869 10.016
R2106 GND.n3045 GND.n3044 10.016
R2107 GND.n1117 GND.n1116 10.016
R2108 GND.n808 GND.n807 10.016
R2109 GND.n1622 GND.n1621 10.016
R2110 GND.n1442 GND.n1441 10.016
R2111 GND.n1703 GND.n1702 9.861
R2112 GND.n1363 GND.n1362 9.861
R2113 GND.n5805 GND.n5804 9.861
R2114 GND.n5625 GND.n5624 9.861
R2115 GND.n1907 GND.n1906 9.861
R2116 GND.n2087 GND.n2086 9.861
R2117 GND.n5217 GND.n5216 9.861
R2118 GND.n5397 GND.n5396 9.861
R2119 GND.n4467 GND.n4466 9.861
R2120 GND.n4838 GND.n4837 9.861
R2121 GND.n5018 GND.n5017 9.861
R2122 GND.n3323 GND.n3322 9.861
R2123 GND.n3716 GND.n3715 9.861
R2124 GND.n4196 GND.n4195 9.861
R2125 GND.n1198 GND.n1197 9.861
R2126 GND.n729 GND.n728 9.861
R2127 GND.n3126 GND.n3125 9.861
R2128 GND.n2791 GND.n2790 9.861
R2129 GND.n7883 GND.n7882 9.3
R2130 GND.n7979 GND.n7978 9.3
R2131 GND.n7841 GND.n7840 9.3
R2132 GND.n7943 GND.n7942 9.3
R2133 GND.n7981 GND.n7980 9.3
R2134 GND.n8009 GND.n8008 9.3
R2135 GND.n7843 GND.n7842 9.3
R2136 GND.n7848 GND.n7847 9.3
R2137 GND.n7909 GND.n7908 9.3
R2138 GND.n7850 GND.n7849 9.3
R2139 GND.n7914 GND.n7913 9.3
R2140 GND.n7855 GND.n7854 9.3
R2141 GND.n7861 GND.n7860 9.3
R2142 GND.n7880 GND.n7879 9.3
R2143 GND.n8019 GND.n8018 9.3
R2144 GND.n7920 GND.n7919 9.3
R2145 GND.n7922 GND.n7921 9.3
R2146 GND.n7954 GND.n7953 9.3
R2147 GND.n8027 GND.n8026 9.3
R2148 GND.n8021 GND.n8020 9.3
R2149 GND.n8002 GND.n8001 9.3
R2150 GND.n7990 GND.n7989 9.3
R2151 GND.n7996 GND.n7995 9.3
R2152 GND.n7870 GND.n7869 9.3
R2153 GND.n7893 GND.n7892 9.3
R2154 GND.n7900 GND.n7899 9.3
R2155 GND.n7873 GND.n7872 9.3
R2156 GND.n7928 GND.n7927 9.3
R2157 GND.n7656 GND.n7655 9.3
R2158 GND.n7752 GND.n7751 9.3
R2159 GND.n7614 GND.n7613 9.3
R2160 GND.n7716 GND.n7715 9.3
R2161 GND.n7754 GND.n7753 9.3
R2162 GND.n7782 GND.n7781 9.3
R2163 GND.n7616 GND.n7615 9.3
R2164 GND.n7621 GND.n7620 9.3
R2165 GND.n7682 GND.n7681 9.3
R2166 GND.n7623 GND.n7622 9.3
R2167 GND.n7687 GND.n7686 9.3
R2168 GND.n7628 GND.n7627 9.3
R2169 GND.n7634 GND.n7633 9.3
R2170 GND.n7653 GND.n7652 9.3
R2171 GND.n7792 GND.n7791 9.3
R2172 GND.n7693 GND.n7692 9.3
R2173 GND.n7695 GND.n7694 9.3
R2174 GND.n7727 GND.n7726 9.3
R2175 GND.n7800 GND.n7799 9.3
R2176 GND.n7794 GND.n7793 9.3
R2177 GND.n7775 GND.n7774 9.3
R2178 GND.n7763 GND.n7762 9.3
R2179 GND.n7769 GND.n7768 9.3
R2180 GND.n7643 GND.n7642 9.3
R2181 GND.n7666 GND.n7665 9.3
R2182 GND.n7673 GND.n7672 9.3
R2183 GND.n7646 GND.n7645 9.3
R2184 GND.n7701 GND.n7700 9.3
R2185 GND.n7429 GND.n7428 9.3
R2186 GND.n7525 GND.n7524 9.3
R2187 GND.n7387 GND.n7386 9.3
R2188 GND.n7489 GND.n7488 9.3
R2189 GND.n7527 GND.n7526 9.3
R2190 GND.n7555 GND.n7554 9.3
R2191 GND.n7389 GND.n7388 9.3
R2192 GND.n7394 GND.n7393 9.3
R2193 GND.n7455 GND.n7454 9.3
R2194 GND.n7396 GND.n7395 9.3
R2195 GND.n7460 GND.n7459 9.3
R2196 GND.n7401 GND.n7400 9.3
R2197 GND.n7407 GND.n7406 9.3
R2198 GND.n7426 GND.n7425 9.3
R2199 GND.n7565 GND.n7564 9.3
R2200 GND.n7466 GND.n7465 9.3
R2201 GND.n7468 GND.n7467 9.3
R2202 GND.n7500 GND.n7499 9.3
R2203 GND.n7573 GND.n7572 9.3
R2204 GND.n7567 GND.n7566 9.3
R2205 GND.n7548 GND.n7547 9.3
R2206 GND.n7536 GND.n7535 9.3
R2207 GND.n7542 GND.n7541 9.3
R2208 GND.n7416 GND.n7415 9.3
R2209 GND.n7439 GND.n7438 9.3
R2210 GND.n7446 GND.n7445 9.3
R2211 GND.n7419 GND.n7418 9.3
R2212 GND.n7474 GND.n7473 9.3
R2213 GND.n7202 GND.n7201 9.3
R2214 GND.n7298 GND.n7297 9.3
R2215 GND.n7160 GND.n7159 9.3
R2216 GND.n7262 GND.n7261 9.3
R2217 GND.n7300 GND.n7299 9.3
R2218 GND.n7328 GND.n7327 9.3
R2219 GND.n7162 GND.n7161 9.3
R2220 GND.n7167 GND.n7166 9.3
R2221 GND.n7228 GND.n7227 9.3
R2222 GND.n7169 GND.n7168 9.3
R2223 GND.n7233 GND.n7232 9.3
R2224 GND.n7174 GND.n7173 9.3
R2225 GND.n7180 GND.n7179 9.3
R2226 GND.n7199 GND.n7198 9.3
R2227 GND.n7338 GND.n7337 9.3
R2228 GND.n7239 GND.n7238 9.3
R2229 GND.n7241 GND.n7240 9.3
R2230 GND.n7273 GND.n7272 9.3
R2231 GND.n7346 GND.n7345 9.3
R2232 GND.n7340 GND.n7339 9.3
R2233 GND.n7321 GND.n7320 9.3
R2234 GND.n7309 GND.n7308 9.3
R2235 GND.n7315 GND.n7314 9.3
R2236 GND.n7189 GND.n7188 9.3
R2237 GND.n7212 GND.n7211 9.3
R2238 GND.n7219 GND.n7218 9.3
R2239 GND.n7192 GND.n7191 9.3
R2240 GND.n7247 GND.n7246 9.3
R2241 GND.n6975 GND.n6974 9.3
R2242 GND.n7071 GND.n7070 9.3
R2243 GND.n6933 GND.n6932 9.3
R2244 GND.n7035 GND.n7034 9.3
R2245 GND.n7073 GND.n7072 9.3
R2246 GND.n7101 GND.n7100 9.3
R2247 GND.n6935 GND.n6934 9.3
R2248 GND.n6940 GND.n6939 9.3
R2249 GND.n7001 GND.n7000 9.3
R2250 GND.n6942 GND.n6941 9.3
R2251 GND.n7006 GND.n7005 9.3
R2252 GND.n6947 GND.n6946 9.3
R2253 GND.n6953 GND.n6952 9.3
R2254 GND.n6972 GND.n6971 9.3
R2255 GND.n7111 GND.n7110 9.3
R2256 GND.n7012 GND.n7011 9.3
R2257 GND.n7014 GND.n7013 9.3
R2258 GND.n7046 GND.n7045 9.3
R2259 GND.n7119 GND.n7118 9.3
R2260 GND.n7113 GND.n7112 9.3
R2261 GND.n7094 GND.n7093 9.3
R2262 GND.n7082 GND.n7081 9.3
R2263 GND.n7088 GND.n7087 9.3
R2264 GND.n6962 GND.n6961 9.3
R2265 GND.n6985 GND.n6984 9.3
R2266 GND.n6992 GND.n6991 9.3
R2267 GND.n6965 GND.n6964 9.3
R2268 GND.n7020 GND.n7019 9.3
R2269 GND.n6748 GND.n6747 9.3
R2270 GND.n6844 GND.n6843 9.3
R2271 GND.n6706 GND.n6705 9.3
R2272 GND.n6808 GND.n6807 9.3
R2273 GND.n6846 GND.n6845 9.3
R2274 GND.n6874 GND.n6873 9.3
R2275 GND.n6708 GND.n6707 9.3
R2276 GND.n6713 GND.n6712 9.3
R2277 GND.n6774 GND.n6773 9.3
R2278 GND.n6715 GND.n6714 9.3
R2279 GND.n6779 GND.n6778 9.3
R2280 GND.n6720 GND.n6719 9.3
R2281 GND.n6726 GND.n6725 9.3
R2282 GND.n6745 GND.n6744 9.3
R2283 GND.n6884 GND.n6883 9.3
R2284 GND.n6785 GND.n6784 9.3
R2285 GND.n6787 GND.n6786 9.3
R2286 GND.n6819 GND.n6818 9.3
R2287 GND.n6892 GND.n6891 9.3
R2288 GND.n6886 GND.n6885 9.3
R2289 GND.n6867 GND.n6866 9.3
R2290 GND.n6855 GND.n6854 9.3
R2291 GND.n6861 GND.n6860 9.3
R2292 GND.n6735 GND.n6734 9.3
R2293 GND.n6758 GND.n6757 9.3
R2294 GND.n6765 GND.n6764 9.3
R2295 GND.n6738 GND.n6737 9.3
R2296 GND.n6793 GND.n6792 9.3
R2297 GND.n6428 GND.n6427 9.3
R2298 GND.n6512 GND.n6511 9.3
R2299 GND.n6374 GND.n6373 9.3
R2300 GND.n6476 GND.n6475 9.3
R2301 GND.n6514 GND.n6513 9.3
R2302 GND.n6542 GND.n6541 9.3
R2303 GND.n6376 GND.n6375 9.3
R2304 GND.n6381 GND.n6380 9.3
R2305 GND.n6453 GND.n6452 9.3
R2306 GND.n6383 GND.n6382 9.3
R2307 GND.n6458 GND.n6457 9.3
R2308 GND.n6436 GND.n6435 9.3
R2309 GND.n6442 GND.n6441 9.3
R2310 GND.n6425 GND.n6424 9.3
R2311 GND.n6552 GND.n6551 9.3
R2312 GND.n6388 GND.n6387 9.3
R2313 GND.n6415 GND.n6414 9.3
R2314 GND.n6487 GND.n6486 9.3
R2315 GND.n6407 GND.n6406 9.3
R2316 GND.n6400 GND.n6399 9.3
R2317 GND.n6396 GND.n6395 9.3
R2318 GND.n6390 GND.n6389 9.3
R2319 GND.n6560 GND.n6559 9.3
R2320 GND.n6554 GND.n6553 9.3
R2321 GND.n6535 GND.n6534 9.3
R2322 GND.n6523 GND.n6522 9.3
R2323 GND.n6529 GND.n6528 9.3
R2324 GND.n6419 GND.n6418 9.3
R2325 GND.n600 GND.n599 9.3
R2326 GND.n607 GND.n606 9.3
R2327 GND.n614 GND.n613 9.3
R2328 GND.n621 GND.n620 9.3
R2329 GND.n628 GND.n627 9.3
R2330 GND.n635 GND.n634 9.3
R2331 GND.n642 GND.n641 9.3
R2332 GND.n647 GND.n646 9.3
R2333 GND.n547 GND.n546 9.3
R2334 GND.n556 GND.n555 9.3
R2335 GND.n541 GND.n540 9.3
R2336 GND.n545 GND.n544 9.3
R2337 GND.n552 GND.n551 9.3
R2338 GND.n558 GND.n557 9.3
R2339 GND.n645 GND.n644 9.3
R2340 GND.n640 GND.n639 9.3
R2341 GND.n638 GND.n637 9.3
R2342 GND.n633 GND.n632 9.3
R2343 GND.n631 GND.n630 9.3
R2344 GND.n626 GND.n625 9.3
R2345 GND.n624 GND.n623 9.3
R2346 GND.n619 GND.n618 9.3
R2347 GND.n617 GND.n616 9.3
R2348 GND.n612 GND.n611 9.3
R2349 GND.n610 GND.n609 9.3
R2350 GND.n605 GND.n604 9.3
R2351 GND.n602 GND.n601 9.3
R2352 GND.n598 GND.n597 9.3
R2353 GND.n569 GND.n568 9.3
R2354 GND.n536 GND.n535 9.3
R2355 GND.n534 GND.n533 9.3
R2356 GND.n530 GND.n529 9.3
R2357 GND.n524 GND.n523 9.3
R2358 GND.n519 GND.n518 9.3
R2359 GND.n514 GND.n513 9.3
R2360 GND.n509 GND.n508 9.3
R2361 GND.n651 GND.n650 9.3
R2362 GND.n649 GND.n648 9.3
R2363 GND.n1039 GND.n1038 9.3
R2364 GND.n1048 GND.n1047 9.3
R2365 GND.n1059 GND.n1058 9.3
R2366 GND.n1071 GND.n1070 9.3
R2367 GND.n1037 GND.n1036 9.3
R2368 GND.n1044 GND.n1043 9.3
R2369 GND.n1066 GND.n1065 9.3
R2370 GND.n1061 GND.n1060 9.3
R2371 GND.n1055 GND.n1054 9.3
R2372 GND.n1050 GND.n1049 9.3
R2373 GND.n950 GND.n949 9.3
R2374 GND.n955 GND.n954 9.3
R2375 GND.n962 GND.n961 9.3
R2376 GND.n969 GND.n968 9.3
R2377 GND.n976 GND.n975 9.3
R2378 GND.n983 GND.n982 9.3
R2379 GND.n990 GND.n989 9.3
R2380 GND.n953 GND.n952 9.3
R2381 GND.n957 GND.n956 9.3
R2382 GND.n960 GND.n959 9.3
R2383 GND.n964 GND.n963 9.3
R2384 GND.n967 GND.n966 9.3
R2385 GND.n971 GND.n970 9.3
R2386 GND.n974 GND.n973 9.3
R2387 GND.n978 GND.n977 9.3
R2388 GND.n981 GND.n980 9.3
R2389 GND.n985 GND.n984 9.3
R2390 GND.n988 GND.n987 9.3
R2391 GND.n992 GND.n991 9.3
R2392 GND.n995 GND.n994 9.3
R2393 GND.n1000 GND.n999 9.3
R2394 GND.n997 GND.n996 9.3
R2395 GND.n948 GND.n947 9.3
R2396 GND.n946 GND.n945 9.3
R2397 GND.n1081 GND.n1080 9.3
R2398 GND.n1086 GND.n1085 9.3
R2399 GND.n1077 GND.n1076 9.3
R2400 GND.n1025 GND.n1024 9.3
R2401 GND.n942 GND.n941 9.3
R2402 GND.n935 GND.n934 9.3
R2403 GND.n928 GND.n927 9.3
R2404 GND.n921 GND.n920 9.3
R2405 GND.n914 GND.n913 9.3
R2406 GND.n907 GND.n906 9.3
R2407 GND.n900 GND.n899 9.3
R2408 GND.n893 GND.n892 9.3
R2409 GND.n884 GND.n883 9.3
R2410 GND.n829 GND.n828 9.3
R2411 GND.n851 GND.n850 9.3
R2412 GND.n862 GND.n861 9.3
R2413 GND.n871 GND.n870 9.3
R2414 GND.n834 GND.n833 9.3
R2415 GND.n839 GND.n838 9.3
R2416 GND.n845 GND.n844 9.3
R2417 GND.n849 GND.n848 9.3
R2418 GND.n856 GND.n855 9.3
R2419 GND.n860 GND.n859 9.3
R2420 GND.n867 GND.n866 9.3
R2421 GND.n873 GND.n872 9.3
R2422 GND.n824 GND.n823 9.3
R2423 GND.n891 GND.n890 9.3
R2424 GND.n895 GND.n894 9.3
R2425 GND.n898 GND.n897 9.3
R2426 GND.n903 GND.n902 9.3
R2427 GND.n905 GND.n904 9.3
R2428 GND.n910 GND.n909 9.3
R2429 GND.n912 GND.n911 9.3
R2430 GND.n917 GND.n916 9.3
R2431 GND.n919 GND.n918 9.3
R2432 GND.n924 GND.n923 9.3
R2433 GND.n926 GND.n925 9.3
R2434 GND.n931 GND.n930 9.3
R2435 GND.n933 GND.n932 9.3
R2436 GND.n938 GND.n937 9.3
R2437 GND.n940 GND.n939 9.3
R2438 GND.n944 GND.n943 9.3
R2439 GND.n6124 GND.n6123 9.3
R2440 GND.n6137 GND.n6136 9.3
R2441 GND.n6135 GND.n6134 9.3
R2442 GND.n6128 GND.n6127 9.3
R2443 GND.n6070 GND.n6069 9.3
R2444 GND.n6077 GND.n6076 9.3
R2445 GND.n6084 GND.n6083 9.3
R2446 GND.n6091 GND.n6090 9.3
R2447 GND.n6098 GND.n6097 9.3
R2448 GND.n6105 GND.n6104 9.3
R2449 GND.n6112 GND.n6111 9.3
R2450 GND.n6117 GND.n6116 9.3
R2451 GND.n5983 GND.n5982 9.3
R2452 GND.n6021 GND.n6020 9.3
R2453 GND.n6025 GND.n6024 9.3
R2454 GND.n6016 GND.n6015 9.3
R2455 GND.n5999 GND.n5998 9.3
R2456 GND.n5988 GND.n5987 9.3
R2457 GND.n5993 GND.n5992 9.3
R2458 GND.n6005 GND.n6004 9.3
R2459 GND.n6003 GND.n6002 9.3
R2460 GND.n6010 GND.n6009 9.3
R2461 GND.n6014 GND.n6013 9.3
R2462 GND.n6027 GND.n6026 9.3
R2463 GND.n6115 GND.n6114 9.3
R2464 GND.n6110 GND.n6109 9.3
R2465 GND.n6108 GND.n6107 9.3
R2466 GND.n6103 GND.n6102 9.3
R2467 GND.n6101 GND.n6100 9.3
R2468 GND.n6096 GND.n6095 9.3
R2469 GND.n6094 GND.n6093 9.3
R2470 GND.n6089 GND.n6088 9.3
R2471 GND.n6087 GND.n6086 9.3
R2472 GND.n6082 GND.n6081 9.3
R2473 GND.n6080 GND.n6079 9.3
R2474 GND.n6075 GND.n6074 9.3
R2475 GND.n6072 GND.n6071 9.3
R2476 GND.n6068 GND.n6067 9.3
R2477 GND.n6038 GND.n6037 9.3
R2478 GND.n5978 GND.n5977 9.3
R2479 GND.n6121 GND.n6120 9.3
R2480 GND.n6119 GND.n6118 9.3
R2481 GND.n1283 GND.n1282 9.3
R2482 GND.n1267 GND.n1266 9.3
R2483 GND.n1281 GND.n1280 9.3
R2484 GND.n1271 GND.n1270 9.3
R2485 GND.n2661 GND.n2660 9.3
R2486 GND.n2670 GND.n2669 9.3
R2487 GND.n2681 GND.n2680 9.3
R2488 GND.n2693 GND.n2692 9.3
R2489 GND.n2659 GND.n2658 9.3
R2490 GND.n2666 GND.n2665 9.3
R2491 GND.n2688 GND.n2687 9.3
R2492 GND.n2683 GND.n2682 9.3
R2493 GND.n2677 GND.n2676 9.3
R2494 GND.n2672 GND.n2671 9.3
R2495 GND.n2572 GND.n2571 9.3
R2496 GND.n2577 GND.n2576 9.3
R2497 GND.n2584 GND.n2583 9.3
R2498 GND.n2591 GND.n2590 9.3
R2499 GND.n2598 GND.n2597 9.3
R2500 GND.n2605 GND.n2604 9.3
R2501 GND.n2612 GND.n2611 9.3
R2502 GND.n2575 GND.n2574 9.3
R2503 GND.n2579 GND.n2578 9.3
R2504 GND.n2582 GND.n2581 9.3
R2505 GND.n2586 GND.n2585 9.3
R2506 GND.n2589 GND.n2588 9.3
R2507 GND.n2593 GND.n2592 9.3
R2508 GND.n2596 GND.n2595 9.3
R2509 GND.n2600 GND.n2599 9.3
R2510 GND.n2603 GND.n2602 9.3
R2511 GND.n2607 GND.n2606 9.3
R2512 GND.n2610 GND.n2609 9.3
R2513 GND.n2614 GND.n2613 9.3
R2514 GND.n2617 GND.n2616 9.3
R2515 GND.n2622 GND.n2621 9.3
R2516 GND.n2619 GND.n2618 9.3
R2517 GND.n2570 GND.n2569 9.3
R2518 GND.n2568 GND.n2567 9.3
R2519 GND.n2703 GND.n2702 9.3
R2520 GND.n2708 GND.n2707 9.3
R2521 GND.n2699 GND.n2698 9.3
R2522 GND.n2647 GND.n2646 9.3
R2523 GND.n2564 GND.n2563 9.3
R2524 GND.n2557 GND.n2556 9.3
R2525 GND.n2550 GND.n2549 9.3
R2526 GND.n2543 GND.n2542 9.3
R2527 GND.n2536 GND.n2535 9.3
R2528 GND.n2529 GND.n2528 9.3
R2529 GND.n2522 GND.n2521 9.3
R2530 GND.n2515 GND.n2514 9.3
R2531 GND.n2506 GND.n2505 9.3
R2532 GND.n2451 GND.n2450 9.3
R2533 GND.n2473 GND.n2472 9.3
R2534 GND.n2484 GND.n2483 9.3
R2535 GND.n2493 GND.n2492 9.3
R2536 GND.n2456 GND.n2455 9.3
R2537 GND.n2461 GND.n2460 9.3
R2538 GND.n2467 GND.n2466 9.3
R2539 GND.n2471 GND.n2470 9.3
R2540 GND.n2478 GND.n2477 9.3
R2541 GND.n2482 GND.n2481 9.3
R2542 GND.n2489 GND.n2488 9.3
R2543 GND.n2495 GND.n2494 9.3
R2544 GND.n2446 GND.n2445 9.3
R2545 GND.n2513 GND.n2512 9.3
R2546 GND.n2517 GND.n2516 9.3
R2547 GND.n2520 GND.n2519 9.3
R2548 GND.n2525 GND.n2524 9.3
R2549 GND.n2527 GND.n2526 9.3
R2550 GND.n2532 GND.n2531 9.3
R2551 GND.n2534 GND.n2533 9.3
R2552 GND.n2539 GND.n2538 9.3
R2553 GND.n2541 GND.n2540 9.3
R2554 GND.n2546 GND.n2545 9.3
R2555 GND.n2548 GND.n2547 9.3
R2556 GND.n2553 GND.n2552 9.3
R2557 GND.n2555 GND.n2554 9.3
R2558 GND.n2560 GND.n2559 9.3
R2559 GND.n2562 GND.n2561 9.3
R2560 GND.n2566 GND.n2565 9.3
R2561 GND.n3952 GND.n3951 9.3
R2562 GND.n3965 GND.n3964 9.3
R2563 GND.n3963 GND.n3962 9.3
R2564 GND.n3956 GND.n3955 9.3
R2565 GND.n3898 GND.n3897 9.3
R2566 GND.n3905 GND.n3904 9.3
R2567 GND.n3912 GND.n3911 9.3
R2568 GND.n3919 GND.n3918 9.3
R2569 GND.n3926 GND.n3925 9.3
R2570 GND.n3933 GND.n3932 9.3
R2571 GND.n3940 GND.n3939 9.3
R2572 GND.n3945 GND.n3944 9.3
R2573 GND.n3811 GND.n3810 9.3
R2574 GND.n3849 GND.n3848 9.3
R2575 GND.n3853 GND.n3852 9.3
R2576 GND.n3844 GND.n3843 9.3
R2577 GND.n3827 GND.n3826 9.3
R2578 GND.n3816 GND.n3815 9.3
R2579 GND.n3821 GND.n3820 9.3
R2580 GND.n3833 GND.n3832 9.3
R2581 GND.n3831 GND.n3830 9.3
R2582 GND.n3838 GND.n3837 9.3
R2583 GND.n3842 GND.n3841 9.3
R2584 GND.n3855 GND.n3854 9.3
R2585 GND.n3943 GND.n3942 9.3
R2586 GND.n3938 GND.n3937 9.3
R2587 GND.n3936 GND.n3935 9.3
R2588 GND.n3931 GND.n3930 9.3
R2589 GND.n3929 GND.n3928 9.3
R2590 GND.n3924 GND.n3923 9.3
R2591 GND.n3922 GND.n3921 9.3
R2592 GND.n3917 GND.n3916 9.3
R2593 GND.n3915 GND.n3914 9.3
R2594 GND.n3910 GND.n3909 9.3
R2595 GND.n3908 GND.n3907 9.3
R2596 GND.n3903 GND.n3902 9.3
R2597 GND.n3900 GND.n3899 9.3
R2598 GND.n3896 GND.n3895 9.3
R2599 GND.n3866 GND.n3865 9.3
R2600 GND.n3806 GND.n3805 9.3
R2601 GND.n3949 GND.n3948 9.3
R2602 GND.n3947 GND.n3946 9.3
R2603 GND.n2172 GND.n2171 9.3
R2604 GND.n2160 GND.n2159 9.3
R2605 GND.n2148 GND.n2147 9.3
R2606 GND.n2136 GND.n2135 9.3
R2607 GND.n2124 GND.n2123 9.3
R2608 GND.n2112 GND.n2111 9.3
R2609 GND.n2094 GND.n2093 9.3
R2610 GND.n2082 GND.n2081 9.3
R2611 GND.n2070 GND.n2069 9.3
R2612 GND.n2058 GND.n2057 9.3
R2613 GND.n2046 GND.n2045 9.3
R2614 GND.n2034 GND.n2033 9.3
R2615 GND.n2022 GND.n2021 9.3
R2616 GND.n2004 GND.n2003 9.3
R2617 GND.n1992 GND.n1991 9.3
R2618 GND.n1980 GND.n1979 9.3
R2619 GND.n1968 GND.n1967 9.3
R2620 GND.n1956 GND.n1955 9.3
R2621 GND.n1944 GND.n1943 9.3
R2622 GND.n1932 GND.n1931 9.3
R2623 GND.n1914 GND.n1913 9.3
R2624 GND.n1902 GND.n1901 9.3
R2625 GND.n1890 GND.n1889 9.3
R2626 GND.n1878 GND.n1877 9.3
R2627 GND.n1866 GND.n1865 9.3
R2628 GND.n1854 GND.n1853 9.3
R2629 GND.n1852 GND.n1851 9.3
R2630 GND.n1864 GND.n1863 9.3
R2631 GND.n1876 GND.n1875 9.3
R2632 GND.n1888 GND.n1887 9.3
R2633 GND.n1900 GND.n1899 9.3
R2634 GND.n1912 GND.n1911 9.3
R2635 GND.n1934 GND.n1933 9.3
R2636 GND.n1946 GND.n1945 9.3
R2637 GND.n1958 GND.n1957 9.3
R2638 GND.n1970 GND.n1969 9.3
R2639 GND.n1982 GND.n1981 9.3
R2640 GND.n1994 GND.n1993 9.3
R2641 GND.n2006 GND.n2005 9.3
R2642 GND.n2020 GND.n2019 9.3
R2643 GND.n2032 GND.n2031 9.3
R2644 GND.n2044 GND.n2043 9.3
R2645 GND.n2056 GND.n2055 9.3
R2646 GND.n2068 GND.n2067 9.3
R2647 GND.n2080 GND.n2079 9.3
R2648 GND.n2092 GND.n2091 9.3
R2649 GND.n2114 GND.n2113 9.3
R2650 GND.n2126 GND.n2125 9.3
R2651 GND.n2138 GND.n2137 9.3
R2652 GND.n2150 GND.n2149 9.3
R2653 GND.n2162 GND.n2161 9.3
R2654 GND.n2174 GND.n2173 9.3
R2655 GND.n2178 GND.n2177 9.3
R2656 GND.n5482 GND.n5481 9.3
R2657 GND.n5470 GND.n5469 9.3
R2658 GND.n5458 GND.n5457 9.3
R2659 GND.n5446 GND.n5445 9.3
R2660 GND.n5434 GND.n5433 9.3
R2661 GND.n5422 GND.n5421 9.3
R2662 GND.n5404 GND.n5403 9.3
R2663 GND.n5392 GND.n5391 9.3
R2664 GND.n5380 GND.n5379 9.3
R2665 GND.n5368 GND.n5367 9.3
R2666 GND.n5356 GND.n5355 9.3
R2667 GND.n5344 GND.n5343 9.3
R2668 GND.n5332 GND.n5331 9.3
R2669 GND.n5314 GND.n5313 9.3
R2670 GND.n5302 GND.n5301 9.3
R2671 GND.n5290 GND.n5289 9.3
R2672 GND.n5278 GND.n5277 9.3
R2673 GND.n5266 GND.n5265 9.3
R2674 GND.n5254 GND.n5253 9.3
R2675 GND.n5242 GND.n5241 9.3
R2676 GND.n5224 GND.n5223 9.3
R2677 GND.n5212 GND.n5211 9.3
R2678 GND.n5200 GND.n5199 9.3
R2679 GND.n5188 GND.n5187 9.3
R2680 GND.n5176 GND.n5175 9.3
R2681 GND.n5164 GND.n5163 9.3
R2682 GND.n5162 GND.n5161 9.3
R2683 GND.n5174 GND.n5173 9.3
R2684 GND.n5186 GND.n5185 9.3
R2685 GND.n5198 GND.n5197 9.3
R2686 GND.n5210 GND.n5209 9.3
R2687 GND.n5222 GND.n5221 9.3
R2688 GND.n5244 GND.n5243 9.3
R2689 GND.n5256 GND.n5255 9.3
R2690 GND.n5268 GND.n5267 9.3
R2691 GND.n5280 GND.n5279 9.3
R2692 GND.n5292 GND.n5291 9.3
R2693 GND.n5304 GND.n5303 9.3
R2694 GND.n5316 GND.n5315 9.3
R2695 GND.n5330 GND.n5329 9.3
R2696 GND.n5342 GND.n5341 9.3
R2697 GND.n5354 GND.n5353 9.3
R2698 GND.n5366 GND.n5365 9.3
R2699 GND.n5378 GND.n5377 9.3
R2700 GND.n5390 GND.n5389 9.3
R2701 GND.n5402 GND.n5401 9.3
R2702 GND.n5424 GND.n5423 9.3
R2703 GND.n5436 GND.n5435 9.3
R2704 GND.n5448 GND.n5447 9.3
R2705 GND.n5460 GND.n5459 9.3
R2706 GND.n5472 GND.n5471 9.3
R2707 GND.n5484 GND.n5483 9.3
R2708 GND.n5488 GND.n5487 9.3
R2709 GND.n5340 GND.n5339 9.3
R2710 GND.n5339 GND.n5338 9.3
R2711 GND.n5352 GND.n5351 9.3
R2712 GND.n5351 GND.n5350 9.3
R2713 GND.n5364 GND.n5363 9.3
R2714 GND.n5363 GND.n5362 9.3
R2715 GND.n5376 GND.n5375 9.3
R2716 GND.n5375 GND.n5374 9.3
R2717 GND.n5388 GND.n5387 9.3
R2718 GND.n5387 GND.n5386 9.3
R2719 GND.n5400 GND.n5399 9.3
R2720 GND.n5399 GND.n5398 9.3
R2721 GND.n5412 GND.n5411 9.3
R2722 GND.n5411 GND.n5410 9.3
R2723 GND.n5420 GND.n5419 9.3
R2724 GND.n5419 GND.n5418 9.3
R2725 GND.n5432 GND.n5431 9.3
R2726 GND.n5431 GND.n5430 9.3
R2727 GND.n5444 GND.n5443 9.3
R2728 GND.n5443 GND.n5442 9.3
R2729 GND.n5456 GND.n5455 9.3
R2730 GND.n5455 GND.n5454 9.3
R2731 GND.n5468 GND.n5467 9.3
R2732 GND.n5467 GND.n5466 9.3
R2733 GND.n5480 GND.n5479 9.3
R2734 GND.n5479 GND.n5478 9.3
R2735 GND.n5156 GND.n5155 9.3
R2736 GND.n5155 GND.n5154 9.3
R2737 GND.n2030 GND.n2029 9.3
R2738 GND.n2029 GND.n2028 9.3
R2739 GND.n2042 GND.n2041 9.3
R2740 GND.n2041 GND.n2040 9.3
R2741 GND.n2054 GND.n2053 9.3
R2742 GND.n2053 GND.n2052 9.3
R2743 GND.n2066 GND.n2065 9.3
R2744 GND.n2065 GND.n2064 9.3
R2745 GND.n2078 GND.n2077 9.3
R2746 GND.n2077 GND.n2076 9.3
R2747 GND.n2090 GND.n2089 9.3
R2748 GND.n2089 GND.n2088 9.3
R2749 GND.n2102 GND.n2101 9.3
R2750 GND.n2101 GND.n2100 9.3
R2751 GND.n2110 GND.n2109 9.3
R2752 GND.n2109 GND.n2108 9.3
R2753 GND.n2122 GND.n2121 9.3
R2754 GND.n2121 GND.n2120 9.3
R2755 GND.n2134 GND.n2133 9.3
R2756 GND.n2133 GND.n2132 9.3
R2757 GND.n2146 GND.n2145 9.3
R2758 GND.n2145 GND.n2144 9.3
R2759 GND.n2158 GND.n2157 9.3
R2760 GND.n2157 GND.n2156 9.3
R2761 GND.n2170 GND.n2169 9.3
R2762 GND.n2169 GND.n2168 9.3
R2763 GND.n1846 GND.n1845 9.3
R2764 GND.n1845 GND.n1844 9.3
R2765 GND.n4738 GND.n4737 9.3
R2766 GND.n4725 GND.n4724 9.3
R2767 GND.n4713 GND.n4712 9.3
R2768 GND.n4700 GND.n4699 9.3
R2769 GND.n4688 GND.n4687 9.3
R2770 GND.n4675 GND.n4674 9.3
R2771 GND.n4656 GND.n4655 9.3
R2772 GND.n4643 GND.n4642 9.3
R2773 GND.n4631 GND.n4630 9.3
R2774 GND.n4618 GND.n4617 9.3
R2775 GND.n4606 GND.n4605 9.3
R2776 GND.n4594 GND.n4593 9.3
R2777 GND.n4582 GND.n4581 9.3
R2778 GND.n4564 GND.n4563 9.3
R2779 GND.n4552 GND.n4551 9.3
R2780 GND.n4540 GND.n4539 9.3
R2781 GND.n4528 GND.n4527 9.3
R2782 GND.n4516 GND.n4515 9.3
R2783 GND.n4504 GND.n4503 9.3
R2784 GND.n4492 GND.n4491 9.3
R2785 GND.n4474 GND.n4473 9.3
R2786 GND.n4462 GND.n4461 9.3
R2787 GND.n4450 GND.n4449 9.3
R2788 GND.n4438 GND.n4437 9.3
R2789 GND.n4426 GND.n4425 9.3
R2790 GND.n4414 GND.n4413 9.3
R2791 GND.n4412 GND.n4411 9.3
R2792 GND.n4424 GND.n4423 9.3
R2793 GND.n4436 GND.n4435 9.3
R2794 GND.n4448 GND.n4447 9.3
R2795 GND.n4460 GND.n4459 9.3
R2796 GND.n4472 GND.n4471 9.3
R2797 GND.n4494 GND.n4493 9.3
R2798 GND.n4506 GND.n4505 9.3
R2799 GND.n4518 GND.n4517 9.3
R2800 GND.n4530 GND.n4529 9.3
R2801 GND.n4542 GND.n4541 9.3
R2802 GND.n4554 GND.n4553 9.3
R2803 GND.n4566 GND.n4565 9.3
R2804 GND.n4580 GND.n4579 9.3
R2805 GND.n4590 GND.n4589 9.3
R2806 GND.n4589 GND.n4588 9.3
R2807 GND.n4592 GND.n4591 9.3
R2808 GND.n4602 GND.n4601 9.3
R2809 GND.n4601 GND.n4600 9.3
R2810 GND.n4604 GND.n4603 9.3
R2811 GND.n4614 GND.n4613 9.3
R2812 GND.n4613 GND.n4612 9.3
R2813 GND.n4616 GND.n4615 9.3
R2814 GND.n4627 GND.n4626 9.3
R2815 GND.n4626 GND.n4625 9.3
R2816 GND.n4629 GND.n4628 9.3
R2817 GND.n4639 GND.n4638 9.3
R2818 GND.n4638 GND.n4637 9.3
R2819 GND.n4641 GND.n4640 9.3
R2820 GND.n4652 GND.n4651 9.3
R2821 GND.n4651 GND.n4650 9.3
R2822 GND.n4654 GND.n4653 9.3
R2823 GND.n4664 GND.n4663 9.3
R2824 GND.n4663 GND.n4662 9.3
R2825 GND.n4673 GND.n4672 9.3
R2826 GND.n4672 GND.n4671 9.3
R2827 GND.n4677 GND.n4676 9.3
R2828 GND.n4686 GND.n4685 9.3
R2829 GND.n4685 GND.n4684 9.3
R2830 GND.n4690 GND.n4689 9.3
R2831 GND.n4698 GND.n4697 9.3
R2832 GND.n4697 GND.n4696 9.3
R2833 GND.n4702 GND.n4701 9.3
R2834 GND.n4711 GND.n4710 9.3
R2835 GND.n4710 GND.n4709 9.3
R2836 GND.n4715 GND.n4714 9.3
R2837 GND.n4723 GND.n4722 9.3
R2838 GND.n4722 GND.n4721 9.3
R2839 GND.n4727 GND.n4726 9.3
R2840 GND.n4736 GND.n4735 9.3
R2841 GND.n4735 GND.n4734 9.3
R2842 GND.n4740 GND.n4739 9.3
R2843 GND.n4744 GND.n4743 9.3
R2844 GND.n4406 GND.n4405 9.3
R2845 GND.n5103 GND.n5102 9.3
R2846 GND.n5091 GND.n5090 9.3
R2847 GND.n5079 GND.n5078 9.3
R2848 GND.n5067 GND.n5066 9.3
R2849 GND.n5055 GND.n5054 9.3
R2850 GND.n5043 GND.n5042 9.3
R2851 GND.n5025 GND.n5024 9.3
R2852 GND.n5013 GND.n5012 9.3
R2853 GND.n5001 GND.n5000 9.3
R2854 GND.n4989 GND.n4988 9.3
R2855 GND.n4977 GND.n4976 9.3
R2856 GND.n4965 GND.n4964 9.3
R2857 GND.n4953 GND.n4952 9.3
R2858 GND.n4935 GND.n4934 9.3
R2859 GND.n4923 GND.n4922 9.3
R2860 GND.n4911 GND.n4910 9.3
R2861 GND.n4899 GND.n4898 9.3
R2862 GND.n4887 GND.n4886 9.3
R2863 GND.n4875 GND.n4874 9.3
R2864 GND.n4863 GND.n4862 9.3
R2865 GND.n4845 GND.n4844 9.3
R2866 GND.n4833 GND.n4832 9.3
R2867 GND.n4821 GND.n4820 9.3
R2868 GND.n4809 GND.n4808 9.3
R2869 GND.n4797 GND.n4796 9.3
R2870 GND.n4785 GND.n4784 9.3
R2871 GND.n4783 GND.n4782 9.3
R2872 GND.n4795 GND.n4794 9.3
R2873 GND.n4807 GND.n4806 9.3
R2874 GND.n4819 GND.n4818 9.3
R2875 GND.n4831 GND.n4830 9.3
R2876 GND.n4843 GND.n4842 9.3
R2877 GND.n4865 GND.n4864 9.3
R2878 GND.n4877 GND.n4876 9.3
R2879 GND.n4889 GND.n4888 9.3
R2880 GND.n4901 GND.n4900 9.3
R2881 GND.n4913 GND.n4912 9.3
R2882 GND.n4925 GND.n4924 9.3
R2883 GND.n4937 GND.n4936 9.3
R2884 GND.n4951 GND.n4950 9.3
R2885 GND.n4961 GND.n4960 9.3
R2886 GND.n4960 GND.n4959 9.3
R2887 GND.n4963 GND.n4962 9.3
R2888 GND.n4973 GND.n4972 9.3
R2889 GND.n4972 GND.n4971 9.3
R2890 GND.n4975 GND.n4974 9.3
R2891 GND.n4985 GND.n4984 9.3
R2892 GND.n4984 GND.n4983 9.3
R2893 GND.n4987 GND.n4986 9.3
R2894 GND.n4997 GND.n4996 9.3
R2895 GND.n4996 GND.n4995 9.3
R2896 GND.n4999 GND.n4998 9.3
R2897 GND.n5009 GND.n5008 9.3
R2898 GND.n5008 GND.n5007 9.3
R2899 GND.n5011 GND.n5010 9.3
R2900 GND.n5021 GND.n5020 9.3
R2901 GND.n5020 GND.n5019 9.3
R2902 GND.n5023 GND.n5022 9.3
R2903 GND.n5033 GND.n5032 9.3
R2904 GND.n5032 GND.n5031 9.3
R2905 GND.n5041 GND.n5040 9.3
R2906 GND.n5040 GND.n5039 9.3
R2907 GND.n5045 GND.n5044 9.3
R2908 GND.n5053 GND.n5052 9.3
R2909 GND.n5052 GND.n5051 9.3
R2910 GND.n5057 GND.n5056 9.3
R2911 GND.n5065 GND.n5064 9.3
R2912 GND.n5064 GND.n5063 9.3
R2913 GND.n5069 GND.n5068 9.3
R2914 GND.n5077 GND.n5076 9.3
R2915 GND.n5076 GND.n5075 9.3
R2916 GND.n5081 GND.n5080 9.3
R2917 GND.n5089 GND.n5088 9.3
R2918 GND.n5088 GND.n5087 9.3
R2919 GND.n5093 GND.n5092 9.3
R2920 GND.n5101 GND.n5100 9.3
R2921 GND.n5100 GND.n5099 9.3
R2922 GND.n5105 GND.n5104 9.3
R2923 GND.n5109 GND.n5108 9.3
R2924 GND.n4777 GND.n4776 9.3
R2925 GND.n4776 GND.n4775 9.3
R2926 GND.n1779 GND.n1778 9.3
R2927 GND.n4793 GND.n4792 9.3
R2928 GND.n4792 GND.n4791 9.3
R2929 GND.n4805 GND.n4804 9.3
R2930 GND.n4804 GND.n4803 9.3
R2931 GND.n4817 GND.n4816 9.3
R2932 GND.n4816 GND.n4815 9.3
R2933 GND.n4829 GND.n4828 9.3
R2934 GND.n4828 GND.n4827 9.3
R2935 GND.n4841 GND.n4840 9.3
R2936 GND.n4840 GND.n4839 9.3
R2937 GND.n4853 GND.n4852 9.3
R2938 GND.n4852 GND.n4851 9.3
R2939 GND.n4861 GND.n4860 9.3
R2940 GND.n4860 GND.n4859 9.3
R2941 GND.n4873 GND.n4872 9.3
R2942 GND.n4872 GND.n4871 9.3
R2943 GND.n4885 GND.n4884 9.3
R2944 GND.n4884 GND.n4883 9.3
R2945 GND.n4897 GND.n4896 9.3
R2946 GND.n4896 GND.n4895 9.3
R2947 GND.n4909 GND.n4908 9.3
R2948 GND.n4908 GND.n4907 9.3
R2949 GND.n4921 GND.n4920 9.3
R2950 GND.n4920 GND.n4919 9.3
R2951 GND.n4933 GND.n4932 9.3
R2952 GND.n4932 GND.n4931 9.3
R2953 GND.n1792 GND.n1791 9.3
R2954 GND.n4422 GND.n4421 9.3
R2955 GND.n4421 GND.n4420 9.3
R2956 GND.n4434 GND.n4433 9.3
R2957 GND.n4433 GND.n4432 9.3
R2958 GND.n4446 GND.n4445 9.3
R2959 GND.n4445 GND.n4444 9.3
R2960 GND.n4458 GND.n4457 9.3
R2961 GND.n4457 GND.n4456 9.3
R2962 GND.n4470 GND.n4469 9.3
R2963 GND.n4469 GND.n4468 9.3
R2964 GND.n4482 GND.n4481 9.3
R2965 GND.n4481 GND.n4480 9.3
R2966 GND.n4490 GND.n4489 9.3
R2967 GND.n4489 GND.n4488 9.3
R2968 GND.n4502 GND.n4501 9.3
R2969 GND.n4501 GND.n4500 9.3
R2970 GND.n4514 GND.n4513 9.3
R2971 GND.n4513 GND.n4512 9.3
R2972 GND.n4526 GND.n4525 9.3
R2973 GND.n4525 GND.n4524 9.3
R2974 GND.n4538 GND.n4537 9.3
R2975 GND.n4537 GND.n4536 9.3
R2976 GND.n4550 GND.n4549 9.3
R2977 GND.n4549 GND.n4548 9.3
R2978 GND.n4562 GND.n4561 9.3
R2979 GND.n4561 GND.n4560 9.3
R2980 GND.n1805 GND.n1804 9.3
R2981 GND.n5172 GND.n5171 9.3
R2982 GND.n5171 GND.n5170 9.3
R2983 GND.n5184 GND.n5183 9.3
R2984 GND.n5183 GND.n5182 9.3
R2985 GND.n5196 GND.n5195 9.3
R2986 GND.n5195 GND.n5194 9.3
R2987 GND.n5208 GND.n5207 9.3
R2988 GND.n5207 GND.n5206 9.3
R2989 GND.n5220 GND.n5219 9.3
R2990 GND.n5219 GND.n5218 9.3
R2991 GND.n5232 GND.n5231 9.3
R2992 GND.n5231 GND.n5230 9.3
R2993 GND.n5240 GND.n5239 9.3
R2994 GND.n5239 GND.n5238 9.3
R2995 GND.n5252 GND.n5251 9.3
R2996 GND.n5251 GND.n5250 9.3
R2997 GND.n5264 GND.n5263 9.3
R2998 GND.n5263 GND.n5262 9.3
R2999 GND.n5276 GND.n5275 9.3
R3000 GND.n5275 GND.n5274 9.3
R3001 GND.n5288 GND.n5287 9.3
R3002 GND.n5287 GND.n5286 9.3
R3003 GND.n5300 GND.n5299 9.3
R3004 GND.n5299 GND.n5298 9.3
R3005 GND.n5312 GND.n5311 9.3
R3006 GND.n5311 GND.n5310 9.3
R3007 GND.n1818 GND.n1817 9.3
R3008 GND.n1862 GND.n1861 9.3
R3009 GND.n1861 GND.n1860 9.3
R3010 GND.n1874 GND.n1873 9.3
R3011 GND.n1873 GND.n1872 9.3
R3012 GND.n1886 GND.n1885 9.3
R3013 GND.n1885 GND.n1884 9.3
R3014 GND.n1898 GND.n1897 9.3
R3015 GND.n1897 GND.n1896 9.3
R3016 GND.n1910 GND.n1909 9.3
R3017 GND.n1909 GND.n1908 9.3
R3018 GND.n1922 GND.n1921 9.3
R3019 GND.n1921 GND.n1920 9.3
R3020 GND.n1930 GND.n1929 9.3
R3021 GND.n1929 GND.n1928 9.3
R3022 GND.n1942 GND.n1941 9.3
R3023 GND.n1941 GND.n1940 9.3
R3024 GND.n1954 GND.n1953 9.3
R3025 GND.n1953 GND.n1952 9.3
R3026 GND.n1966 GND.n1965 9.3
R3027 GND.n1965 GND.n1964 9.3
R3028 GND.n1978 GND.n1977 9.3
R3029 GND.n1977 GND.n1976 9.3
R3030 GND.n1990 GND.n1989 9.3
R3031 GND.n1989 GND.n1988 9.3
R3032 GND.n2002 GND.n2001 9.3
R3033 GND.n2001 GND.n2000 9.3
R3034 GND.n3237 GND.n3236 9.3
R3035 GND.n3250 GND.n3249 9.3
R3036 GND.n3262 GND.n3261 9.3
R3037 GND.n3274 GND.n3273 9.3
R3038 GND.n3286 GND.n3285 9.3
R3039 GND.n3298 GND.n3297 9.3
R3040 GND.n3316 GND.n3315 9.3
R3041 GND.n3328 GND.n3327 9.3
R3042 GND.n3340 GND.n3339 9.3
R3043 GND.n3352 GND.n3351 9.3
R3044 GND.n3364 GND.n3363 9.3
R3045 GND.n3376 GND.n3375 9.3
R3046 GND.n3388 GND.n3387 9.3
R3047 GND.n3406 GND.n3405 9.3
R3048 GND.n3418 GND.n3417 9.3
R3049 GND.n3431 GND.n3430 9.3
R3050 GND.n3443 GND.n3442 9.3
R3051 GND.n3456 GND.n3455 9.3
R3052 GND.n3468 GND.n3467 9.3
R3053 GND.n3481 GND.n3480 9.3
R3054 GND.n3500 GND.n3499 9.3
R3055 GND.n3513 GND.n3512 9.3
R3056 GND.n3525 GND.n3524 9.3
R3057 GND.n3538 GND.n3537 9.3
R3058 GND.n3550 GND.n3549 9.3
R3059 GND.n3563 GND.n3562 9.3
R3060 GND.n3577 GND.n3576 9.3
R3061 GND.n3565 GND.n3564 9.3
R3062 GND.n3561 GND.n3560 9.3
R3063 GND.n3560 GND.n3559 9.3
R3064 GND.n3552 GND.n3551 9.3
R3065 GND.n3548 GND.n3547 9.3
R3066 GND.n3547 GND.n3546 9.3
R3067 GND.n3540 GND.n3539 9.3
R3068 GND.n3536 GND.n3535 9.3
R3069 GND.n3535 GND.n3534 9.3
R3070 GND.n3527 GND.n3526 9.3
R3071 GND.n3523 GND.n3522 9.3
R3072 GND.n3522 GND.n3521 9.3
R3073 GND.n3515 GND.n3514 9.3
R3074 GND.n3511 GND.n3510 9.3
R3075 GND.n3510 GND.n3509 9.3
R3076 GND.n3502 GND.n3501 9.3
R3077 GND.n3498 GND.n3497 9.3
R3078 GND.n3497 GND.n3496 9.3
R3079 GND.n3490 GND.n3489 9.3
R3080 GND.n3489 GND.n3488 9.3
R3081 GND.n3479 GND.n3478 9.3
R3082 GND.n3477 GND.n3476 9.3
R3083 GND.n3476 GND.n3475 9.3
R3084 GND.n3466 GND.n3465 9.3
R3085 GND.n3464 GND.n3463 9.3
R3086 GND.n3463 GND.n3462 9.3
R3087 GND.n3454 GND.n3453 9.3
R3088 GND.n3452 GND.n3451 9.3
R3089 GND.n3451 GND.n3450 9.3
R3090 GND.n3441 GND.n3440 9.3
R3091 GND.n3439 GND.n3438 9.3
R3092 GND.n3438 GND.n3437 9.3
R3093 GND.n3429 GND.n3428 9.3
R3094 GND.n3427 GND.n3426 9.3
R3095 GND.n3426 GND.n3425 9.3
R3096 GND.n3416 GND.n3415 9.3
R3097 GND.n3414 GND.n3413 9.3
R3098 GND.n3413 GND.n3412 9.3
R3099 GND.n3404 GND.n3403 9.3
R3100 GND.n3390 GND.n3389 9.3
R3101 GND.n3386 GND.n3385 9.3
R3102 GND.n3385 GND.n3384 9.3
R3103 GND.n3378 GND.n3377 9.3
R3104 GND.n3374 GND.n3373 9.3
R3105 GND.n3373 GND.n3372 9.3
R3106 GND.n3366 GND.n3365 9.3
R3107 GND.n3362 GND.n3361 9.3
R3108 GND.n3361 GND.n3360 9.3
R3109 GND.n3354 GND.n3353 9.3
R3110 GND.n3350 GND.n3349 9.3
R3111 GND.n3349 GND.n3348 9.3
R3112 GND.n3342 GND.n3341 9.3
R3113 GND.n3338 GND.n3337 9.3
R3114 GND.n3337 GND.n3336 9.3
R3115 GND.n3330 GND.n3329 9.3
R3116 GND.n3326 GND.n3325 9.3
R3117 GND.n3325 GND.n3324 9.3
R3118 GND.n3318 GND.n3317 9.3
R3119 GND.n3314 GND.n3313 9.3
R3120 GND.n3313 GND.n3312 9.3
R3121 GND.n3306 GND.n3305 9.3
R3122 GND.n3305 GND.n3304 9.3
R3123 GND.n3296 GND.n3295 9.3
R3124 GND.n3294 GND.n3293 9.3
R3125 GND.n3293 GND.n3292 9.3
R3126 GND.n3284 GND.n3283 9.3
R3127 GND.n3282 GND.n3281 9.3
R3128 GND.n3281 GND.n3280 9.3
R3129 GND.n3272 GND.n3271 9.3
R3130 GND.n3270 GND.n3269 9.3
R3131 GND.n3269 GND.n3268 9.3
R3132 GND.n3260 GND.n3259 9.3
R3133 GND.n3258 GND.n3257 9.3
R3134 GND.n3257 GND.n3256 9.3
R3135 GND.n3248 GND.n3247 9.3
R3136 GND.n3246 GND.n3245 9.3
R3137 GND.n3245 GND.n3244 9.3
R3138 GND.n3235 GND.n3234 9.3
R3139 GND.n3231 GND.n3230 9.3
R3140 GND.n3207 GND.n3206 9.3
R3141 GND.n5539 GND.n5538 9.3
R3142 GND.n5552 GND.n5551 9.3
R3143 GND.n5564 GND.n5563 9.3
R3144 GND.n5576 GND.n5575 9.3
R3145 GND.n5588 GND.n5587 9.3
R3146 GND.n5600 GND.n5599 9.3
R3147 GND.n5618 GND.n5617 9.3
R3148 GND.n5630 GND.n5629 9.3
R3149 GND.n5642 GND.n5641 9.3
R3150 GND.n5654 GND.n5653 9.3
R3151 GND.n5666 GND.n5665 9.3
R3152 GND.n5678 GND.n5677 9.3
R3153 GND.n5690 GND.n5689 9.3
R3154 GND.n5708 GND.n5707 9.3
R3155 GND.n5720 GND.n5719 9.3
R3156 GND.n5732 GND.n5731 9.3
R3157 GND.n5744 GND.n5743 9.3
R3158 GND.n5756 GND.n5755 9.3
R3159 GND.n5768 GND.n5767 9.3
R3160 GND.n5780 GND.n5779 9.3
R3161 GND.n5798 GND.n5797 9.3
R3162 GND.n5810 GND.n5809 9.3
R3163 GND.n5822 GND.n5821 9.3
R3164 GND.n5834 GND.n5833 9.3
R3165 GND.n5846 GND.n5845 9.3
R3166 GND.n5858 GND.n5857 9.3
R3167 GND.n5872 GND.n5871 9.3
R3168 GND.n5860 GND.n5859 9.3
R3169 GND.n5856 GND.n5855 9.3
R3170 GND.n5855 GND.n5854 9.3
R3171 GND.n5848 GND.n5847 9.3
R3172 GND.n5844 GND.n5843 9.3
R3173 GND.n5843 GND.n5842 9.3
R3174 GND.n5836 GND.n5835 9.3
R3175 GND.n5832 GND.n5831 9.3
R3176 GND.n5831 GND.n5830 9.3
R3177 GND.n5824 GND.n5823 9.3
R3178 GND.n5820 GND.n5819 9.3
R3179 GND.n5819 GND.n5818 9.3
R3180 GND.n5812 GND.n5811 9.3
R3181 GND.n5808 GND.n5807 9.3
R3182 GND.n5807 GND.n5806 9.3
R3183 GND.n5800 GND.n5799 9.3
R3184 GND.n5796 GND.n5795 9.3
R3185 GND.n5795 GND.n5794 9.3
R3186 GND.n5788 GND.n5787 9.3
R3187 GND.n5787 GND.n5786 9.3
R3188 GND.n5778 GND.n5777 9.3
R3189 GND.n5776 GND.n5775 9.3
R3190 GND.n5775 GND.n5774 9.3
R3191 GND.n5766 GND.n5765 9.3
R3192 GND.n5764 GND.n5763 9.3
R3193 GND.n5763 GND.n5762 9.3
R3194 GND.n5754 GND.n5753 9.3
R3195 GND.n5752 GND.n5751 9.3
R3196 GND.n5751 GND.n5750 9.3
R3197 GND.n5742 GND.n5741 9.3
R3198 GND.n5740 GND.n5739 9.3
R3199 GND.n5739 GND.n5738 9.3
R3200 GND.n5730 GND.n5729 9.3
R3201 GND.n5728 GND.n5727 9.3
R3202 GND.n5727 GND.n5726 9.3
R3203 GND.n5718 GND.n5717 9.3
R3204 GND.n5716 GND.n5715 9.3
R3205 GND.n5715 GND.n5714 9.3
R3206 GND.n5706 GND.n5705 9.3
R3207 GND.n5692 GND.n5691 9.3
R3208 GND.n5688 GND.n5687 9.3
R3209 GND.n5687 GND.n5686 9.3
R3210 GND.n5680 GND.n5679 9.3
R3211 GND.n5676 GND.n5675 9.3
R3212 GND.n5675 GND.n5674 9.3
R3213 GND.n5668 GND.n5667 9.3
R3214 GND.n5664 GND.n5663 9.3
R3215 GND.n5663 GND.n5662 9.3
R3216 GND.n5656 GND.n5655 9.3
R3217 GND.n5652 GND.n5651 9.3
R3218 GND.n5651 GND.n5650 9.3
R3219 GND.n5644 GND.n5643 9.3
R3220 GND.n5640 GND.n5639 9.3
R3221 GND.n5639 GND.n5638 9.3
R3222 GND.n5632 GND.n5631 9.3
R3223 GND.n5628 GND.n5627 9.3
R3224 GND.n5627 GND.n5626 9.3
R3225 GND.n5620 GND.n5619 9.3
R3226 GND.n5616 GND.n5615 9.3
R3227 GND.n5615 GND.n5614 9.3
R3228 GND.n5608 GND.n5607 9.3
R3229 GND.n5607 GND.n5606 9.3
R3230 GND.n5598 GND.n5597 9.3
R3231 GND.n5596 GND.n5595 9.3
R3232 GND.n5595 GND.n5594 9.3
R3233 GND.n5586 GND.n5585 9.3
R3234 GND.n5584 GND.n5583 9.3
R3235 GND.n5583 GND.n5582 9.3
R3236 GND.n5574 GND.n5573 9.3
R3237 GND.n5572 GND.n5571 9.3
R3238 GND.n5571 GND.n5570 9.3
R3239 GND.n5562 GND.n5561 9.3
R3240 GND.n5560 GND.n5559 9.3
R3241 GND.n5559 GND.n5558 9.3
R3242 GND.n5550 GND.n5549 9.3
R3243 GND.n5548 GND.n5547 9.3
R3244 GND.n5547 GND.n5546 9.3
R3245 GND.n5537 GND.n5536 9.3
R3246 GND.n5533 GND.n5532 9.3
R3247 GND.n1833 GND.n1832 9.3
R3248 GND.n2415 GND.n2414 9.3
R3249 GND.n2408 GND.n2407 9.3
R3250 GND.n2401 GND.n2400 9.3
R3251 GND.n2394 GND.n2393 9.3
R3252 GND.n2387 GND.n2386 9.3
R3253 GND.n2380 GND.n2379 9.3
R3254 GND.n2373 GND.n2372 9.3
R3255 GND.n2366 GND.n2365 9.3
R3256 GND.n2302 GND.n2301 9.3
R3257 GND.n2313 GND.n2312 9.3
R3258 GND.n2322 GND.n2321 9.3
R3259 GND.n2364 GND.n2363 9.3
R3260 GND.n2324 GND.n2323 9.3
R3261 GND.n2318 GND.n2317 9.3
R3262 GND.n2311 GND.n2310 9.3
R3263 GND.n2307 GND.n2306 9.3
R3264 GND.n2300 GND.n2299 9.3
R3265 GND.n2296 GND.n2295 9.3
R3266 GND.n2290 GND.n2289 9.3
R3267 GND.n2285 GND.n2284 9.3
R3268 GND.n2280 GND.n2279 9.3
R3269 GND.n2275 GND.n2274 9.3
R3270 GND.n2368 GND.n2367 9.3
R3271 GND.n2371 GND.n2370 9.3
R3272 GND.n2376 GND.n2375 9.3
R3273 GND.n2378 GND.n2377 9.3
R3274 GND.n2383 GND.n2382 9.3
R3275 GND.n2385 GND.n2384 9.3
R3276 GND.n2390 GND.n2389 9.3
R3277 GND.n2392 GND.n2391 9.3
R3278 GND.n2397 GND.n2396 9.3
R3279 GND.n2399 GND.n2398 9.3
R3280 GND.n2404 GND.n2403 9.3
R3281 GND.n2406 GND.n2405 9.3
R3282 GND.n2411 GND.n2410 9.3
R3283 GND.n2413 GND.n2412 9.3
R3284 GND.n2417 GND.n2416 9.3
R3285 GND.n2335 GND.n2334 9.3
R3286 GND.n3006 GND.n3005 9.3
R3287 GND.n3001 GND.n3000 9.3
R3288 GND.n2994 GND.n2993 9.3
R3289 GND.n2987 GND.n2986 9.3
R3290 GND.n2980 GND.n2979 9.3
R3291 GND.n2973 GND.n2972 9.3
R3292 GND.n2966 GND.n2965 9.3
R3293 GND.n2959 GND.n2958 9.3
R3294 GND.n2945 GND.n2944 9.3
R3295 GND.n2943 GND.n2942 9.3
R3296 GND.n3004 GND.n3003 9.3
R3297 GND.n2999 GND.n2998 9.3
R3298 GND.n2997 GND.n2996 9.3
R3299 GND.n2992 GND.n2991 9.3
R3300 GND.n2990 GND.n2989 9.3
R3301 GND.n2985 GND.n2984 9.3
R3302 GND.n2983 GND.n2982 9.3
R3303 GND.n2978 GND.n2977 9.3
R3304 GND.n2976 GND.n2975 9.3
R3305 GND.n2971 GND.n2970 9.3
R3306 GND.n2969 GND.n2968 9.3
R3307 GND.n2964 GND.n2963 9.3
R3308 GND.n2962 GND.n2961 9.3
R3309 GND.n2957 GND.n2956 9.3
R3310 GND.n2951 GND.n2950 9.3
R3311 GND.n2939 GND.n2938 9.3
R3312 GND.n2929 GND.n2928 9.3
R3313 GND.n2932 GND.n2931 9.3
R3314 GND.n2934 GND.n2933 9.3
R3315 GND.n3008 GND.n3007 9.3
R3316 GND.n3010 GND.n3009 9.3
R3317 GND.n2913 GND.n2912 9.3
R3318 GND.n2909 GND.n2908 9.3
R3319 GND.n2904 GND.n2903 9.3
R3320 GND.n2900 GND.n2899 9.3
R3321 GND.n2919 GND.n2918 9.3
R3322 GND.n2922 GND.n2921 9.3
R3323 GND.n2924 GND.n2923 9.3
R3324 GND.n2265 GND.n2264 9.3
R3325 GND.n2259 GND.n2258 9.3
R3326 GND.n2263 GND.n2262 9.3
R3327 GND.n2269 GND.n2268 9.3
R3328 GND.n4117 GND.n4116 9.3
R3329 GND.n4112 GND.n4111 9.3
R3330 GND.n4105 GND.n4104 9.3
R3331 GND.n4098 GND.n4097 9.3
R3332 GND.n4091 GND.n4090 9.3
R3333 GND.n4084 GND.n4083 9.3
R3334 GND.n4077 GND.n4076 9.3
R3335 GND.n4070 GND.n4069 9.3
R3336 GND.n4054 GND.n4053 9.3
R3337 GND.n4115 GND.n4114 9.3
R3338 GND.n4110 GND.n4109 9.3
R3339 GND.n4108 GND.n4107 9.3
R3340 GND.n4103 GND.n4102 9.3
R3341 GND.n4101 GND.n4100 9.3
R3342 GND.n4096 GND.n4095 9.3
R3343 GND.n4094 GND.n4093 9.3
R3344 GND.n4089 GND.n4088 9.3
R3345 GND.n4087 GND.n4086 9.3
R3346 GND.n4082 GND.n4081 9.3
R3347 GND.n4080 GND.n4079 9.3
R3348 GND.n4075 GND.n4074 9.3
R3349 GND.n4073 GND.n4072 9.3
R3350 GND.n4068 GND.n4067 9.3
R3351 GND.n4062 GND.n4061 9.3
R3352 GND.n4056 GND.n4055 9.3
R3353 GND.n4050 GND.n4049 9.3
R3354 GND.n4040 GND.n4039 9.3
R3355 GND.n4043 GND.n4042 9.3
R3356 GND.n4045 GND.n4044 9.3
R3357 GND.n4119 GND.n4118 9.3
R3358 GND.n4121 GND.n4120 9.3
R3359 GND.n4024 GND.n4023 9.3
R3360 GND.n4020 GND.n4019 9.3
R3361 GND.n4015 GND.n4014 9.3
R3362 GND.n3988 GND.n3987 9.3
R3363 GND.n4030 GND.n4029 9.3
R3364 GND.n4033 GND.n4032 9.3
R3365 GND.n4035 GND.n4034 9.3
R3366 GND.n2896 GND.n2895 9.3
R3367 GND.n2421 GND.n2420 9.3
R3368 GND.n4304 GND.n4303 9.3
R3369 GND.n4300 GND.n4299 9.3
R3370 GND.n4293 GND.n4292 9.3
R3371 GND.n4281 GND.n4280 9.3
R3372 GND.n4269 GND.n4268 9.3
R3373 GND.n4257 GND.n4256 9.3
R3374 GND.n4245 GND.n4244 9.3
R3375 GND.n4233 GND.n4232 9.3
R3376 GND.n4221 GND.n4220 9.3
R3377 GND.n4203 GND.n4202 9.3
R3378 GND.n4191 GND.n4190 9.3
R3379 GND.n4179 GND.n4178 9.3
R3380 GND.n4167 GND.n4166 9.3
R3381 GND.n4155 GND.n4154 9.3
R3382 GND.n4143 GND.n4142 9.3
R3383 GND.n4130 GND.n4129 9.3
R3384 GND.n3769 GND.n3768 9.3
R3385 GND.n3757 GND.n3756 9.3
R3386 GND.n3745 GND.n3744 9.3
R3387 GND.n3733 GND.n3732 9.3
R3388 GND.n3721 GND.n3720 9.3
R3389 GND.n3709 GND.n3708 9.3
R3390 GND.n3691 GND.n3690 9.3
R3391 GND.n3679 GND.n3678 9.3
R3392 GND.n3667 GND.n3666 9.3
R3393 GND.n3655 GND.n3654 9.3
R3394 GND.n3643 GND.n3642 9.3
R3395 GND.n3631 GND.n3630 9.3
R3396 GND.n3619 GND.n3618 9.3
R3397 GND.n3775 GND.n3774 9.3
R3398 GND.n3771 GND.n3770 9.3
R3399 GND.n3759 GND.n3758 9.3
R3400 GND.n3747 GND.n3746 9.3
R3401 GND.n3735 GND.n3734 9.3
R3402 GND.n3723 GND.n3722 9.3
R3403 GND.n3711 GND.n3710 9.3
R3404 GND.n3689 GND.n3688 9.3
R3405 GND.n3677 GND.n3676 9.3
R3406 GND.n3665 GND.n3664 9.3
R3407 GND.n3653 GND.n3652 9.3
R3408 GND.n3641 GND.n3640 9.3
R3409 GND.n3629 GND.n3628 9.3
R3410 GND.n2443 GND.n2442 9.3
R3411 GND.n4128 GND.n4127 9.3
R3412 GND.n4141 GND.n4140 9.3
R3413 GND.n4153 GND.n4152 9.3
R3414 GND.n4165 GND.n4164 9.3
R3415 GND.n4177 GND.n4176 9.3
R3416 GND.n4189 GND.n4188 9.3
R3417 GND.n4201 GND.n4200 9.3
R3418 GND.n4223 GND.n4222 9.3
R3419 GND.n4235 GND.n4234 9.3
R3420 GND.n4247 GND.n4246 9.3
R3421 GND.n4259 GND.n4258 9.3
R3422 GND.n4271 GND.n4270 9.3
R3423 GND.n4283 GND.n4282 9.3
R3424 GND.n4295 GND.n4294 9.3
R3425 GND.n3616 GND.n3615 9.3
R3426 GND.n3767 GND.n3766 9.3
R3427 GND.n3766 GND.n3765 9.3
R3428 GND.n3755 GND.n3754 9.3
R3429 GND.n3754 GND.n3753 9.3
R3430 GND.n3743 GND.n3742 9.3
R3431 GND.n3742 GND.n3741 9.3
R3432 GND.n3731 GND.n3730 9.3
R3433 GND.n3730 GND.n3729 9.3
R3434 GND.n3719 GND.n3718 9.3
R3435 GND.n3718 GND.n3717 9.3
R3436 GND.n3707 GND.n3706 9.3
R3437 GND.n3706 GND.n3705 9.3
R3438 GND.n3699 GND.n3698 9.3
R3439 GND.n3698 GND.n3697 9.3
R3440 GND.n3687 GND.n3686 9.3
R3441 GND.n3686 GND.n3685 9.3
R3442 GND.n3675 GND.n3674 9.3
R3443 GND.n3674 GND.n3673 9.3
R3444 GND.n3663 GND.n3662 9.3
R3445 GND.n3662 GND.n3661 9.3
R3446 GND.n3651 GND.n3650 9.3
R3447 GND.n3650 GND.n3649 9.3
R3448 GND.n3639 GND.n3638 9.3
R3449 GND.n3638 GND.n3637 9.3
R3450 GND.n3627 GND.n3626 9.3
R3451 GND.n3626 GND.n3625 9.3
R3452 GND.n4139 GND.n4138 9.3
R3453 GND.n4138 GND.n4137 9.3
R3454 GND.n4151 GND.n4150 9.3
R3455 GND.n4150 GND.n4149 9.3
R3456 GND.n4163 GND.n4162 9.3
R3457 GND.n4162 GND.n4161 9.3
R3458 GND.n4175 GND.n4174 9.3
R3459 GND.n4174 GND.n4173 9.3
R3460 GND.n4187 GND.n4186 9.3
R3461 GND.n4186 GND.n4185 9.3
R3462 GND.n4199 GND.n4198 9.3
R3463 GND.n4198 GND.n4197 9.3
R3464 GND.n4211 GND.n4210 9.3
R3465 GND.n4210 GND.n4209 9.3
R3466 GND.n4219 GND.n4218 9.3
R3467 GND.n4218 GND.n4217 9.3
R3468 GND.n4231 GND.n4230 9.3
R3469 GND.n4230 GND.n4229 9.3
R3470 GND.n4243 GND.n4242 9.3
R3471 GND.n4242 GND.n4241 9.3
R3472 GND.n4255 GND.n4254 9.3
R3473 GND.n4254 GND.n4253 9.3
R3474 GND.n4267 GND.n4266 9.3
R3475 GND.n4266 GND.n4265 9.3
R3476 GND.n4279 GND.n4278 9.3
R3477 GND.n4278 GND.n4277 9.3
R3478 GND.n4291 GND.n4290 9.3
R3479 GND.n4290 GND.n4289 9.3
R3480 GND.n3191 GND.n3190 9.3
R3481 GND.n3179 GND.n3178 9.3
R3482 GND.n3167 GND.n3166 9.3
R3483 GND.n3155 GND.n3154 9.3
R3484 GND.n3143 GND.n3142 9.3
R3485 GND.n3131 GND.n3130 9.3
R3486 GND.n3119 GND.n3118 9.3
R3487 GND.n3101 GND.n3100 9.3
R3488 GND.n3089 GND.n3088 9.3
R3489 GND.n3077 GND.n3076 9.3
R3490 GND.n3065 GND.n3064 9.3
R3491 GND.n3053 GND.n3052 9.3
R3492 GND.n3041 GND.n3040 9.3
R3493 GND.n3028 GND.n3027 9.3
R3494 GND.n2725 GND.n2724 9.3
R3495 GND.n2738 GND.n2737 9.3
R3496 GND.n2750 GND.n2749 9.3
R3497 GND.n2762 GND.n2761 9.3
R3498 GND.n2774 GND.n2773 9.3
R3499 GND.n2786 GND.n2785 9.3
R3500 GND.n2798 GND.n2797 9.3
R3501 GND.n2816 GND.n2815 9.3
R3502 GND.n2828 GND.n2827 9.3
R3503 GND.n2840 GND.n2839 9.3
R3504 GND.n2852 GND.n2851 9.3
R3505 GND.n2864 GND.n2863 9.3
R3506 GND.n2876 GND.n2875 9.3
R3507 GND.n2888 GND.n2887 9.3
R3508 GND.n3193 GND.n3192 9.3
R3509 GND.n3189 GND.n3188 9.3
R3510 GND.n3188 GND.n3187 9.3
R3511 GND.n2890 GND.n2889 9.3
R3512 GND.n2886 GND.n2885 9.3
R3513 GND.n2885 GND.n2884 9.3
R3514 GND.n2878 GND.n2877 9.3
R3515 GND.n2874 GND.n2873 9.3
R3516 GND.n2873 GND.n2872 9.3
R3517 GND.n2866 GND.n2865 9.3
R3518 GND.n2862 GND.n2861 9.3
R3519 GND.n2861 GND.n2860 9.3
R3520 GND.n2854 GND.n2853 9.3
R3521 GND.n2850 GND.n2849 9.3
R3522 GND.n2849 GND.n2848 9.3
R3523 GND.n2842 GND.n2841 9.3
R3524 GND.n2838 GND.n2837 9.3
R3525 GND.n2837 GND.n2836 9.3
R3526 GND.n2830 GND.n2829 9.3
R3527 GND.n2826 GND.n2825 9.3
R3528 GND.n2825 GND.n2824 9.3
R3529 GND.n2818 GND.n2817 9.3
R3530 GND.n2814 GND.n2813 9.3
R3531 GND.n2813 GND.n2812 9.3
R3532 GND.n2806 GND.n2805 9.3
R3533 GND.n2805 GND.n2804 9.3
R3534 GND.n2796 GND.n2795 9.3
R3535 GND.n2794 GND.n2793 9.3
R3536 GND.n2793 GND.n2792 9.3
R3537 GND.n2784 GND.n2783 9.3
R3538 GND.n2782 GND.n2781 9.3
R3539 GND.n2781 GND.n2780 9.3
R3540 GND.n2772 GND.n2771 9.3
R3541 GND.n2770 GND.n2769 9.3
R3542 GND.n2769 GND.n2768 9.3
R3543 GND.n2760 GND.n2759 9.3
R3544 GND.n2758 GND.n2757 9.3
R3545 GND.n2757 GND.n2756 9.3
R3546 GND.n2748 GND.n2747 9.3
R3547 GND.n2746 GND.n2745 9.3
R3548 GND.n2745 GND.n2744 9.3
R3549 GND.n2736 GND.n2735 9.3
R3550 GND.n2734 GND.n2733 9.3
R3551 GND.n2733 GND.n2732 9.3
R3552 GND.n2712 GND.n2711 9.3
R3553 GND.n3026 GND.n3025 9.3
R3554 GND.n3037 GND.n3036 9.3
R3555 GND.n3036 GND.n3035 9.3
R3556 GND.n3035 GND.n3034 9.3
R3557 GND.n3039 GND.n3038 9.3
R3558 GND.n3049 GND.n3048 9.3
R3559 GND.n3048 GND.n3047 9.3
R3560 GND.n3051 GND.n3050 9.3
R3561 GND.n3061 GND.n3060 9.3
R3562 GND.n3060 GND.n3059 9.3
R3563 GND.n3063 GND.n3062 9.3
R3564 GND.n3073 GND.n3072 9.3
R3565 GND.n3072 GND.n3071 9.3
R3566 GND.n3075 GND.n3074 9.3
R3567 GND.n3085 GND.n3084 9.3
R3568 GND.n3084 GND.n3083 9.3
R3569 GND.n3087 GND.n3086 9.3
R3570 GND.n3097 GND.n3096 9.3
R3571 GND.n3096 GND.n3095 9.3
R3572 GND.n3099 GND.n3098 9.3
R3573 GND.n3109 GND.n3108 9.3
R3574 GND.n3108 GND.n3107 9.3
R3575 GND.n3117 GND.n3116 9.3
R3576 GND.n3116 GND.n3115 9.3
R3577 GND.n3121 GND.n3120 9.3
R3578 GND.n3129 GND.n3128 9.3
R3579 GND.n3128 GND.n3127 9.3
R3580 GND.n3133 GND.n3132 9.3
R3581 GND.n3141 GND.n3140 9.3
R3582 GND.n3140 GND.n3139 9.3
R3583 GND.n3145 GND.n3144 9.3
R3584 GND.n3153 GND.n3152 9.3
R3585 GND.n3152 GND.n3151 9.3
R3586 GND.n3157 GND.n3156 9.3
R3587 GND.n3165 GND.n3164 9.3
R3588 GND.n3164 GND.n3163 9.3
R3589 GND.n3169 GND.n3168 9.3
R3590 GND.n3177 GND.n3176 9.3
R3591 GND.n3176 GND.n3175 9.3
R3592 GND.n3181 GND.n3180 9.3
R3593 GND.n6158 GND.n6157 9.3
R3594 GND.n676 GND.n675 9.3
R3595 GND.n688 GND.n687 9.3
R3596 GND.n700 GND.n699 9.3
R3597 GND.n712 GND.n711 9.3
R3598 GND.n724 GND.n723 9.3
R3599 GND.n736 GND.n735 9.3
R3600 GND.n754 GND.n753 9.3
R3601 GND.n766 GND.n765 9.3
R3602 GND.n778 GND.n777 9.3
R3603 GND.n790 GND.n789 9.3
R3604 GND.n802 GND.n801 9.3
R3605 GND.n814 GND.n813 9.3
R3606 GND.n1101 GND.n1100 9.3
R3607 GND.n1113 GND.n1112 9.3
R3608 GND.n1125 GND.n1124 9.3
R3609 GND.n1137 GND.n1136 9.3
R3610 GND.n1149 GND.n1148 9.3
R3611 GND.n1161 GND.n1160 9.3
R3612 GND.n1173 GND.n1172 9.3
R3613 GND.n1191 GND.n1190 9.3
R3614 GND.n1203 GND.n1202 9.3
R3615 GND.n1215 GND.n1214 9.3
R3616 GND.n1227 GND.n1226 9.3
R3617 GND.n1239 GND.n1238 9.3
R3618 GND.n1251 GND.n1250 9.3
R3619 GND.n1257 GND.n1256 9.3
R3620 GND.n821 GND.n820 9.3
R3621 GND.n1109 GND.n1108 9.3
R3622 GND.n1108 GND.n1107 9.3
R3623 GND.n1111 GND.n1110 9.3
R3624 GND.n1121 GND.n1120 9.3
R3625 GND.n1120 GND.n1119 9.3
R3626 GND.n1123 GND.n1122 9.3
R3627 GND.n1133 GND.n1132 9.3
R3628 GND.n1132 GND.n1131 9.3
R3629 GND.n1135 GND.n1134 9.3
R3630 GND.n1145 GND.n1144 9.3
R3631 GND.n1144 GND.n1143 9.3
R3632 GND.n1147 GND.n1146 9.3
R3633 GND.n1157 GND.n1156 9.3
R3634 GND.n1156 GND.n1155 9.3
R3635 GND.n1159 GND.n1158 9.3
R3636 GND.n1169 GND.n1168 9.3
R3637 GND.n1168 GND.n1167 9.3
R3638 GND.n1171 GND.n1170 9.3
R3639 GND.n1181 GND.n1180 9.3
R3640 GND.n1180 GND.n1179 9.3
R3641 GND.n1189 GND.n1188 9.3
R3642 GND.n1188 GND.n1187 9.3
R3643 GND.n1193 GND.n1192 9.3
R3644 GND.n1201 GND.n1200 9.3
R3645 GND.n1200 GND.n1199 9.3
R3646 GND.n1205 GND.n1204 9.3
R3647 GND.n1213 GND.n1212 9.3
R3648 GND.n1212 GND.n1211 9.3
R3649 GND.n1217 GND.n1216 9.3
R3650 GND.n1225 GND.n1224 9.3
R3651 GND.n1224 GND.n1223 9.3
R3652 GND.n1229 GND.n1228 9.3
R3653 GND.n1237 GND.n1236 9.3
R3654 GND.n1236 GND.n1235 9.3
R3655 GND.n1241 GND.n1240 9.3
R3656 GND.n1249 GND.n1248 9.3
R3657 GND.n1248 GND.n1247 9.3
R3658 GND.n1253 GND.n1252 9.3
R3659 GND.n1098 GND.n1097 9.3
R3660 GND.n6160 GND.n6159 9.3
R3661 GND.n6156 GND.n6155 9.3
R3662 GND.n6155 GND.n6154 9.3
R3663 GND.n674 GND.n673 9.3
R3664 GND.n684 GND.n683 9.3
R3665 GND.n683 GND.n682 9.3
R3666 GND.n686 GND.n685 9.3
R3667 GND.n696 GND.n695 9.3
R3668 GND.n695 GND.n694 9.3
R3669 GND.n698 GND.n697 9.3
R3670 GND.n708 GND.n707 9.3
R3671 GND.n707 GND.n706 9.3
R3672 GND.n710 GND.n709 9.3
R3673 GND.n720 GND.n719 9.3
R3674 GND.n719 GND.n718 9.3
R3675 GND.n722 GND.n721 9.3
R3676 GND.n732 GND.n731 9.3
R3677 GND.n731 GND.n730 9.3
R3678 GND.n734 GND.n733 9.3
R3679 GND.n744 GND.n743 9.3
R3680 GND.n743 GND.n742 9.3
R3681 GND.n752 GND.n751 9.3
R3682 GND.n751 GND.n750 9.3
R3683 GND.n756 GND.n755 9.3
R3684 GND.n764 GND.n763 9.3
R3685 GND.n763 GND.n762 9.3
R3686 GND.n768 GND.n767 9.3
R3687 GND.n776 GND.n775 9.3
R3688 GND.n775 GND.n774 9.3
R3689 GND.n780 GND.n779 9.3
R3690 GND.n788 GND.n787 9.3
R3691 GND.n787 GND.n786 9.3
R3692 GND.n792 GND.n791 9.3
R3693 GND.n800 GND.n799 9.3
R3694 GND.n799 GND.n798 9.3
R3695 GND.n804 GND.n803 9.3
R3696 GND.n812 GND.n811 9.3
R3697 GND.n811 GND.n810 9.3
R3698 GND.n816 GND.n815 9.3
R3699 GND.n669 GND.n668 9.3
R3700 GND.n668 GND.n667 9.3
R3701 GND.n819 GND.n671 9.3
R3702 GND.n1463 GND.n1462 9.3
R3703 GND.n1449 GND.n1448 9.3
R3704 GND.n1436 GND.n1435 9.3
R3705 GND.n1424 GND.n1423 9.3
R3706 GND.n1412 GND.n1411 9.3
R3707 GND.n1400 GND.n1399 9.3
R3708 GND.n1388 GND.n1387 9.3
R3709 GND.n1370 GND.n1369 9.3
R3710 GND.n1358 GND.n1357 9.3
R3711 GND.n1346 GND.n1345 9.3
R3712 GND.n1334 GND.n1333 9.3
R3713 GND.n1322 GND.n1321 9.3
R3714 GND.n1310 GND.n1309 9.3
R3715 GND.n1297 GND.n1296 9.3
R3716 GND.n1614 GND.n1613 9.3
R3717 GND.n1613 GND.n1612 9.3
R3718 GND.n1612 GND.n1611 9.3
R3719 GND.n1618 GND.n1617 9.3
R3720 GND.n1630 GND.n1629 9.3
R3721 GND.n1642 GND.n1641 9.3
R3722 GND.n1654 GND.n1653 9.3
R3723 GND.n1666 GND.n1665 9.3
R3724 GND.n1678 GND.n1677 9.3
R3725 GND.n1696 GND.n1695 9.3
R3726 GND.n1708 GND.n1707 9.3
R3727 GND.n1720 GND.n1719 9.3
R3728 GND.n1732 GND.n1731 9.3
R3729 GND.n1744 GND.n1743 9.3
R3730 GND.n1756 GND.n1755 9.3
R3731 GND.n1770 GND.n1769 9.3
R3732 GND.n1616 GND.n1615 9.3
R3733 GND.n1626 GND.n1625 9.3
R3734 GND.n1625 GND.n1624 9.3
R3735 GND.n1628 GND.n1627 9.3
R3736 GND.n1638 GND.n1637 9.3
R3737 GND.n1637 GND.n1636 9.3
R3738 GND.n1640 GND.n1639 9.3
R3739 GND.n1650 GND.n1649 9.3
R3740 GND.n1649 GND.n1648 9.3
R3741 GND.n1652 GND.n1651 9.3
R3742 GND.n1662 GND.n1661 9.3
R3743 GND.n1661 GND.n1660 9.3
R3744 GND.n1664 GND.n1663 9.3
R3745 GND.n1674 GND.n1673 9.3
R3746 GND.n1673 GND.n1672 9.3
R3747 GND.n1676 GND.n1675 9.3
R3748 GND.n1686 GND.n1685 9.3
R3749 GND.n1685 GND.n1684 9.3
R3750 GND.n1694 GND.n1693 9.3
R3751 GND.n1693 GND.n1692 9.3
R3752 GND.n1698 GND.n1697 9.3
R3753 GND.n1706 GND.n1705 9.3
R3754 GND.n1705 GND.n1704 9.3
R3755 GND.n1710 GND.n1709 9.3
R3756 GND.n1718 GND.n1717 9.3
R3757 GND.n1717 GND.n1716 9.3
R3758 GND.n1722 GND.n1721 9.3
R3759 GND.n1730 GND.n1729 9.3
R3760 GND.n1729 GND.n1728 9.3
R3761 GND.n1734 GND.n1733 9.3
R3762 GND.n1742 GND.n1741 9.3
R3763 GND.n1741 GND.n1740 9.3
R3764 GND.n1746 GND.n1745 9.3
R3765 GND.n1754 GND.n1753 9.3
R3766 GND.n1753 GND.n1752 9.3
R3767 GND.n1758 GND.n1757 9.3
R3768 GND.n1766 GND.n1765 9.3
R3769 GND.n1765 GND.n1764 9.3
R3770 GND.n1768 GND.n1767 9.3
R3771 GND.n1605 GND.n1604 9.3
R3772 GND.n1603 GND.n1602 9.3
R3773 GND.n1451 GND.n1450 9.3
R3774 GND.n1447 GND.n1446 9.3
R3775 GND.n1446 GND.n1445 9.3
R3776 GND.n1438 GND.n1437 9.3
R3777 GND.n1434 GND.n1433 9.3
R3778 GND.n1433 GND.n1432 9.3
R3779 GND.n1426 GND.n1425 9.3
R3780 GND.n1422 GND.n1421 9.3
R3781 GND.n1421 GND.n1420 9.3
R3782 GND.n1414 GND.n1413 9.3
R3783 GND.n1410 GND.n1409 9.3
R3784 GND.n1409 GND.n1408 9.3
R3785 GND.n1402 GND.n1401 9.3
R3786 GND.n1398 GND.n1397 9.3
R3787 GND.n1397 GND.n1396 9.3
R3788 GND.n1390 GND.n1389 9.3
R3789 GND.n1386 GND.n1385 9.3
R3790 GND.n1385 GND.n1384 9.3
R3791 GND.n1378 GND.n1377 9.3
R3792 GND.n1377 GND.n1376 9.3
R3793 GND.n1368 GND.n1367 9.3
R3794 GND.n1366 GND.n1365 9.3
R3795 GND.n1365 GND.n1364 9.3
R3796 GND.n1356 GND.n1355 9.3
R3797 GND.n1354 GND.n1353 9.3
R3798 GND.n1353 GND.n1352 9.3
R3799 GND.n1344 GND.n1343 9.3
R3800 GND.n1342 GND.n1341 9.3
R3801 GND.n1341 GND.n1340 9.3
R3802 GND.n1332 GND.n1331 9.3
R3803 GND.n1330 GND.n1329 9.3
R3804 GND.n1329 GND.n1328 9.3
R3805 GND.n1320 GND.n1319 9.3
R3806 GND.n1318 GND.n1317 9.3
R3807 GND.n1317 GND.n1316 9.3
R3808 GND.n1308 GND.n1307 9.3
R3809 GND.n1306 GND.n1305 9.3
R3810 GND.n1305 GND.n1304 9.3
R3811 GND.n1288 GND.n1287 9.3
R3812 GND.n1461 GND.n1460 9.3
R3813 GND.n1459 GND.n1458 9.3
R3814 GND.n1458 GND.n1457 9.3
R3815 GND.n1587 GND.n1586 9.3
R3816 GND.n1580 GND.n1579 9.3
R3817 GND.n1573 GND.n1572 9.3
R3818 GND.n1566 GND.n1565 9.3
R3819 GND.n1559 GND.n1558 9.3
R3820 GND.n1552 GND.n1551 9.3
R3821 GND.n1545 GND.n1544 9.3
R3822 GND.n1538 GND.n1537 9.3
R3823 GND.n1517 GND.n1516 9.3
R3824 GND.n1508 GND.n1507 9.3
R3825 GND.n1519 GND.n1518 9.3
R3826 GND.n1513 GND.n1512 9.3
R3827 GND.n1506 GND.n1505 9.3
R3828 GND.n1502 GND.n1501 9.3
R3829 GND.n1530 GND.n1529 9.3
R3830 GND.n1536 GND.n1535 9.3
R3831 GND.n1541 GND.n1540 9.3
R3832 GND.n1543 GND.n1542 9.3
R3833 GND.n1548 GND.n1547 9.3
R3834 GND.n1550 GND.n1549 9.3
R3835 GND.n1555 GND.n1554 9.3
R3836 GND.n1557 GND.n1556 9.3
R3837 GND.n1562 GND.n1561 9.3
R3838 GND.n1564 GND.n1563 9.3
R3839 GND.n1569 GND.n1568 9.3
R3840 GND.n1571 GND.n1570 9.3
R3841 GND.n1576 GND.n1575 9.3
R3842 GND.n1578 GND.n1577 9.3
R3843 GND.n1583 GND.n1582 9.3
R3844 GND.n1585 GND.n1584 9.3
R3845 GND.n1589 GND.n1588 9.3
R3846 GND.n1486 GND.n1485 9.3
R3847 GND.n1482 GND.n1481 9.3
R3848 GND.n1477 GND.n1476 9.3
R3849 GND.n1473 GND.n1472 9.3
R3850 GND.n1492 GND.n1491 9.3
R3851 GND.n1495 GND.n1494 9.3
R3852 GND.n1497 GND.n1496 9.3
R3853 GND.n493 GND.n492 9.3
R3854 GND.n499 GND.n498 9.3
R3855 GND.n497 GND.n496 9.3
R3856 GND.n503 GND.n502 9.3
R3857 GND.n6171 GND.n6170 9.3
R3858 GND.n6176 GND.n6175 9.3
R3859 GND.n6183 GND.n6182 9.3
R3860 GND.n6190 GND.n6189 9.3
R3861 GND.n6197 GND.n6196 9.3
R3862 GND.n6204 GND.n6203 9.3
R3863 GND.n6211 GND.n6210 9.3
R3864 GND.n6218 GND.n6217 9.3
R3865 GND.n6240 GND.n6239 9.3
R3866 GND.n6249 GND.n6248 9.3
R3867 GND.n6174 GND.n6173 9.3
R3868 GND.n6178 GND.n6177 9.3
R3869 GND.n6181 GND.n6180 9.3
R3870 GND.n6185 GND.n6184 9.3
R3871 GND.n6188 GND.n6187 9.3
R3872 GND.n6192 GND.n6191 9.3
R3873 GND.n6195 GND.n6194 9.3
R3874 GND.n6199 GND.n6198 9.3
R3875 GND.n6202 GND.n6201 9.3
R3876 GND.n6206 GND.n6205 9.3
R3877 GND.n6209 GND.n6208 9.3
R3878 GND.n6213 GND.n6212 9.3
R3879 GND.n6216 GND.n6215 9.3
R3880 GND.n6221 GND.n6220 9.3
R3881 GND.n6227 GND.n6226 9.3
R3882 GND.n6238 GND.n6237 9.3
R3883 GND.n6245 GND.n6244 9.3
R3884 GND.n6251 GND.n6250 9.3
R3885 GND.n6256 GND.n6255 9.3
R3886 GND.n6169 GND.n6168 9.3
R3887 GND.n6167 GND.n6166 9.3
R3888 GND.n6272 GND.n6271 9.3
R3889 GND.n6278 GND.n6277 9.3
R3890 GND.n6282 GND.n6281 9.3
R3891 GND.n6310 GND.n6309 9.3
R3892 GND.n6267 GND.n6266 9.3
R3893 GND.n6262 GND.n6261 9.3
R3894 GND.n6260 GND.n6259 9.3
R3895 GND.n6313 GND.n6312 9.3
R3896 GND.n661 GND.n660 9.3
R3897 GND.n655 GND.n654 9.3
R3898 GND.n1469 GND.n1468 9.3
R3899 GND.n8223 GND.n8222 9.3
R3900 GND.n8257 GND.n8256 9.3
R3901 GND.n8287 GND.n8286 9.3
R3902 GND.n8246 GND.n8245 9.3
R3903 GND.n8229 GND.n8228 9.3
R3904 GND.n8233 GND.n8232 9.3
R3905 GND.n8240 GND.n8239 9.3
R3906 GND.n8244 GND.n8243 9.3
R3907 GND.n8251 GND.n8250 9.3
R3908 GND.n8255 GND.n8254 9.3
R3909 GND.n8263 GND.n8262 9.3
R3910 GND.n8285 GND.n8284 9.3
R3911 GND.n8277 GND.n8276 9.3
R3912 GND.n8218 GND.n8217 9.3
R3913 GND.n8174 GND.n8173 9.3
R3914 GND.n8185 GND.n8184 9.3
R3915 GND.n8191 GND.n8190 9.3
R3916 GND.n8183 GND.n8182 9.3
R3917 GND.n8179 GND.n8178 9.3
R3918 GND.n8172 GND.n8171 9.3
R3919 GND.n8168 GND.n8167 9.3
R3920 GND.n8161 GND.n8160 9.3
R3921 GND.n8157 GND.n8156 9.3
R3922 GND.n8151 GND.n8150 9.3
R3923 GND.n8146 GND.n8145 9.3
R3924 GND.n8204 GND.n8203 9.3
R3925 GND.n8212 GND.n8211 9.3
R3926 GND.n8214 GND.n8213 9.3
R3927 GND.n8330 GND.n8329 9.3
R3928 GND.n8353 GND.n8352 9.3
R3929 GND.n8336 GND.n8335 9.3
R3930 GND.n8340 GND.n8339 9.3
R3931 GND.n8347 GND.n8346 9.3
R3932 GND.n8351 GND.n8350 9.3
R3933 GND.n8358 GND.n8357 9.3
R3934 GND.n8362 GND.n8361 9.3
R3935 GND.n8364 GND.n8363 9.3
R3936 GND.n8394 GND.n8393 9.3
R3937 GND.n8370 GND.n8369 9.3
R3938 GND.n8392 GND.n8391 9.3
R3939 GND.n8384 GND.n8383 9.3
R3940 GND.n8325 GND.n8324 9.3
R3941 GND.n8425 GND.n8424 9.3
R3942 GND.n8419 GND.n8418 9.3
R3943 GND.n8430 GND.n8429 9.3
R3944 GND.n8408 GND.n8407 9.3
R3945 GND.n8402 GND.n8401 9.3
R3946 GND.n8397 GND.n8396 9.3
R3947 GND.n8412 GND.n8411 9.3
R3948 GND.n8436 GND.n8435 9.3
R3949 GND.n8465 GND.n8464 9.3
R3950 GND.n8434 GND.n8433 9.3
R3951 GND.n8442 GND.n8441 9.3
R3952 GND.n8463 GND.n8462 9.3
R3953 GND.n8455 GND.n8454 9.3
R3954 GND.n8423 GND.n8422 9.3
R3955 GND.n8515 GND.n8514 9.3
R3956 GND.n8538 GND.n8537 9.3
R3957 GND.n8521 GND.n8520 9.3
R3958 GND.n8525 GND.n8524 9.3
R3959 GND.n8532 GND.n8531 9.3
R3960 GND.n8536 GND.n8535 9.3
R3961 GND.n8543 GND.n8542 9.3
R3962 GND.n8547 GND.n8546 9.3
R3963 GND.n8549 GND.n8548 9.3
R3964 GND.n8579 GND.n8578 9.3
R3965 GND.n8555 GND.n8554 9.3
R3966 GND.n8577 GND.n8576 9.3
R3967 GND.n8569 GND.n8568 9.3
R3968 GND.n8510 GND.n8509 9.3
R3969 GND.n8610 GND.n8609 9.3
R3970 GND.n8604 GND.n8603 9.3
R3971 GND.n8615 GND.n8614 9.3
R3972 GND.n8593 GND.n8592 9.3
R3973 GND.n8587 GND.n8586 9.3
R3974 GND.n8582 GND.n8581 9.3
R3975 GND.n8597 GND.n8596 9.3
R3976 GND.n8621 GND.n8620 9.3
R3977 GND.n8650 GND.n8649 9.3
R3978 GND.n8619 GND.n8618 9.3
R3979 GND.n8627 GND.n8626 9.3
R3980 GND.n8648 GND.n8647 9.3
R3981 GND.n8640 GND.n8639 9.3
R3982 GND.n8608 GND.n8607 9.3
R3983 GND.n8700 GND.n8699 9.3
R3984 GND.n8723 GND.n8722 9.3
R3985 GND.n8706 GND.n8705 9.3
R3986 GND.n8710 GND.n8709 9.3
R3987 GND.n8717 GND.n8716 9.3
R3988 GND.n8721 GND.n8720 9.3
R3989 GND.n8728 GND.n8727 9.3
R3990 GND.n8732 GND.n8731 9.3
R3991 GND.n8734 GND.n8733 9.3
R3992 GND.n8764 GND.n8763 9.3
R3993 GND.n8740 GND.n8739 9.3
R3994 GND.n8762 GND.n8761 9.3
R3995 GND.n8754 GND.n8753 9.3
R3996 GND.n8695 GND.n8694 9.3
R3997 GND.n8795 GND.n8794 9.3
R3998 GND.n8789 GND.n8788 9.3
R3999 GND.n8800 GND.n8799 9.3
R4000 GND.n8778 GND.n8777 9.3
R4001 GND.n8772 GND.n8771 9.3
R4002 GND.n8767 GND.n8766 9.3
R4003 GND.n8782 GND.n8781 9.3
R4004 GND.n8806 GND.n8805 9.3
R4005 GND.n8835 GND.n8834 9.3
R4006 GND.n8804 GND.n8803 9.3
R4007 GND.n8812 GND.n8811 9.3
R4008 GND.n8833 GND.n8832 9.3
R4009 GND.n8825 GND.n8824 9.3
R4010 GND.n8793 GND.n8792 9.3
R4011 GND.n8885 GND.n8884 9.3
R4012 GND.n8908 GND.n8907 9.3
R4013 GND.n8891 GND.n8890 9.3
R4014 GND.n8895 GND.n8894 9.3
R4015 GND.n8902 GND.n8901 9.3
R4016 GND.n8906 GND.n8905 9.3
R4017 GND.n8913 GND.n8912 9.3
R4018 GND.n8917 GND.n8916 9.3
R4019 GND.n8919 GND.n8918 9.3
R4020 GND.n8949 GND.n8948 9.3
R4021 GND.n8925 GND.n8924 9.3
R4022 GND.n8947 GND.n8946 9.3
R4023 GND.n8939 GND.n8938 9.3
R4024 GND.n8880 GND.n8879 9.3
R4025 GND.n8980 GND.n8979 9.3
R4026 GND.n8974 GND.n8973 9.3
R4027 GND.n8985 GND.n8984 9.3
R4028 GND.n8963 GND.n8962 9.3
R4029 GND.n8957 GND.n8956 9.3
R4030 GND.n8952 GND.n8951 9.3
R4031 GND.n8967 GND.n8966 9.3
R4032 GND.n8991 GND.n8990 9.3
R4033 GND.n9020 GND.n9019 9.3
R4034 GND.n8989 GND.n8988 9.3
R4035 GND.n8997 GND.n8996 9.3
R4036 GND.n9018 GND.n9017 9.3
R4037 GND.n9010 GND.n9009 9.3
R4038 GND.n8978 GND.n8977 9.3
R4039 GND.n9070 GND.n9069 9.3
R4040 GND.n9093 GND.n9092 9.3
R4041 GND.n9076 GND.n9075 9.3
R4042 GND.n9080 GND.n9079 9.3
R4043 GND.n9087 GND.n9086 9.3
R4044 GND.n9091 GND.n9090 9.3
R4045 GND.n9098 GND.n9097 9.3
R4046 GND.n9102 GND.n9101 9.3
R4047 GND.n9104 GND.n9103 9.3
R4048 GND.n9134 GND.n9133 9.3
R4049 GND.n9110 GND.n9109 9.3
R4050 GND.n9132 GND.n9131 9.3
R4051 GND.n9124 GND.n9123 9.3
R4052 GND.n9065 GND.n9064 9.3
R4053 GND.n9165 GND.n9164 9.3
R4054 GND.n9159 GND.n9158 9.3
R4055 GND.n9170 GND.n9169 9.3
R4056 GND.n9148 GND.n9147 9.3
R4057 GND.n9142 GND.n9141 9.3
R4058 GND.n9137 GND.n9136 9.3
R4059 GND.n9152 GND.n9151 9.3
R4060 GND.n9176 GND.n9175 9.3
R4061 GND.n9205 GND.n9204 9.3
R4062 GND.n9174 GND.n9173 9.3
R4063 GND.n9182 GND.n9181 9.3
R4064 GND.n9203 GND.n9202 9.3
R4065 GND.n9195 GND.n9194 9.3
R4066 GND.n9163 GND.n9162 9.3
R4067 GND.n31 GND.n30 9.3
R4068 GND.n54 GND.n53 9.3
R4069 GND.n37 GND.n36 9.3
R4070 GND.n41 GND.n40 9.3
R4071 GND.n48 GND.n47 9.3
R4072 GND.n52 GND.n51 9.3
R4073 GND.n59 GND.n58 9.3
R4074 GND.n63 GND.n62 9.3
R4075 GND.n65 GND.n64 9.3
R4076 GND.n95 GND.n94 9.3
R4077 GND.n71 GND.n70 9.3
R4078 GND.n93 GND.n92 9.3
R4079 GND.n85 GND.n84 9.3
R4080 GND.n26 GND.n25 9.3
R4081 GND.n126 GND.n125 9.3
R4082 GND.n120 GND.n119 9.3
R4083 GND.n131 GND.n130 9.3
R4084 GND.n109 GND.n108 9.3
R4085 GND.n103 GND.n102 9.3
R4086 GND.n98 GND.n97 9.3
R4087 GND.n113 GND.n112 9.3
R4088 GND.n137 GND.n136 9.3
R4089 GND.n166 GND.n165 9.3
R4090 GND.n135 GND.n134 9.3
R4091 GND.n143 GND.n142 9.3
R4092 GND.n164 GND.n163 9.3
R4093 GND.n156 GND.n155 9.3
R4094 GND.n124 GND.n123 9.3
R4095 GND.n5531 GND.n1835 9.154
R4096 GND.n2180 GND.n2179 9.154
R4097 GND.n2008 GND.n2007 9.154
R4098 GND.n2011 GND.n2010 9.154
R4099 GND.n2014 GND.n2013 9.154
R4100 GND.n2017 GND.n2016 9.154
R4101 GND.n1821 GND.n1810 9.154
R4102 GND.n5490 GND.n5489 9.154
R4103 GND.n5318 GND.n5317 9.154
R4104 GND.n5321 GND.n5320 9.154
R4105 GND.n5324 GND.n5323 9.154
R4106 GND.n5327 GND.n5326 9.154
R4107 GND.n1808 GND.n1797 9.154
R4108 GND.n4746 GND.n4745 9.154
R4109 GND.n4568 GND.n4567 9.154
R4110 GND.n4571 GND.n4570 9.154
R4111 GND.n4574 GND.n4573 9.154
R4112 GND.n4577 GND.n4576 9.154
R4113 GND.n1795 GND.n1784 9.154
R4114 GND.n5111 GND.n5110 9.154
R4115 GND.n4939 GND.n4938 9.154
R4116 GND.n4942 GND.n4941 9.154
R4117 GND.n4945 GND.n4944 9.154
R4118 GND.n4948 GND.n4947 9.154
R4119 GND.n1782 GND.n1771 9.154
R4120 GND.n3229 GND.n3209 9.154
R4121 GND.n3401 GND.n3400 9.154
R4122 GND.n3398 GND.n3397 9.154
R4123 GND.n3395 GND.n3394 9.154
R4124 GND.n3392 GND.n3391 9.154
R4125 GND.n3580 GND.n3569 9.154
R4126 GND.n5703 GND.n5702 9.154
R4127 GND.n5700 GND.n5699 9.154
R4128 GND.n5697 GND.n5696 9.154
R4129 GND.n5694 GND.n5693 9.154
R4130 GND.n5875 GND.n5864 9.154
R4131 GND.n2441 GND.n2440 9.154
R4132 GND.n3975 GND.n3974 9.154
R4133 GND.n3972 GND.n3971 9.154
R4134 GND.n3969 GND.n3968 9.154
R4135 GND.n3777 GND.n3776 9.154
R4136 GND.n4125 GND.n4124 9.154
R4137 GND.n3195 GND.n3194 9.154
R4138 GND.n2892 GND.n2891 9.154
R4139 GND.n3014 GND.n3013 9.154
R4140 GND.n3017 GND.n3016 9.154
R4141 GND.n3020 GND.n3019 9.154
R4142 GND.n3023 GND.n3022 9.154
R4143 GND.n3198 GND.n3197 9.154
R4144 GND.n3798 GND.n3797 9.154
R4145 GND.n3792 GND.n3791 9.154
R4146 GND.n3785 GND.n3784 9.154
R4147 GND.n3782 GND.n3780 9.154
R4148 GND.n3607 GND.n3606 9.154
R4149 GND.n3604 GND.n3603 9.154
R4150 GND.n3601 GND.n3600 9.154
R4151 GND.n3598 GND.n3597 9.154
R4152 GND.n3594 GND.n3593 9.154
R4153 GND.n3589 GND.n3588 9.154
R4154 GND.n3586 GND.n3585 9.154
R4155 GND.n3583 GND.n3582 9.154
R4156 GND.n1824 GND.n1823 9.154
R4157 GND.n5881 GND.n5880 9.154
R4158 GND.n5884 GND.n5883 9.154
R4159 GND.n5887 GND.n5886 9.154
R4160 GND.n5890 GND.n5889 9.154
R4161 GND.n5893 GND.n5892 9.154
R4162 GND.n5899 GND.n5898 9.154
R4163 GND.n5902 GND.n5901 9.154
R4164 GND.n5905 GND.n5904 9.154
R4165 GND.n5908 GND.n5907 9.154
R4166 GND.n5911 GND.n5910 9.154
R4167 GND.n5917 GND.n5916 9.154
R4168 GND.n5920 GND.n5919 9.154
R4169 GND.n5923 GND.n5922 9.154
R4170 GND.n5926 GND.n5925 9.154
R4171 GND.n5929 GND.n5928 9.154
R4172 GND.n5935 GND.n5934 9.154
R4173 GND.n5938 GND.n5937 9.154
R4174 GND.n5941 GND.n5940 9.154
R4175 GND.n5944 GND.n5943 9.154
R4176 GND.n5947 GND.n5946 9.154
R4177 GND.n5953 GND.n5952 9.154
R4178 GND.n5956 GND.n5955 9.154
R4179 GND.n5959 GND.n5958 9.154
R4180 GND.n5962 GND.n5961 9.154
R4181 GND.n5965 GND.n5964 9.154
R4182 GND.n5973 GND.n5972 9.154
R4183 GND.n1285 GND.n1284 9.154
R4184 GND.n1273 GND.n1272 9.154
R4185 GND.n1264 GND.n1090 9.154
R4186 GND.n1263 GND.n1262 9.154
R4187 GND.n6141 GND.n6140 9.154
R4188 GND.n6144 GND.n6143 9.154
R4189 GND.n6147 GND.n6146 9.154
R4190 GND.n1259 GND.n1258 9.154
R4191 GND.n2256 GND.n2255 9.154
R4192 GND.n2251 GND.n2250 9.154
R4193 GND.n2424 GND.n2423 9.154
R4194 GND.n2438 GND.n2437 9.154
R4195 GND.n2433 GND.n2432 9.154
R4196 GND.n2430 GND.n2429 9.154
R4197 GND.n2427 GND.n2426 9.154
R4198 GND.n3211 GND.n3210 9.154
R4199 GND.n3225 GND.n3224 9.154
R4200 GND.n3220 GND.n3219 9.154
R4201 GND.n3217 GND.n3216 9.154
R4202 GND.n3214 GND.n3213 9.154
R4203 GND.n1837 GND.n1836 9.154
R4204 GND.n5527 GND.n5526 9.154
R4205 GND.n5522 GND.n5521 9.154
R4206 GND.n5519 GND.n5518 9.154
R4207 GND.n5516 GND.n5515 9.154
R4208 GND.n5513 GND.n5512 9.154
R4209 GND.n5509 GND.n5508 9.154
R4210 GND.n5504 GND.n5503 9.154
R4211 GND.n5501 GND.n5500 9.154
R4212 GND.n5497 GND.n5496 9.154
R4213 GND.n5494 GND.n5493 9.154
R4214 GND.n5147 GND.n5146 9.154
R4215 GND.n5142 GND.n5141 9.154
R4216 GND.n5139 GND.n5138 9.154
R4217 GND.n5136 GND.n5135 9.154
R4218 GND.n5133 GND.n5132 9.154
R4219 GND.n5129 GND.n5128 9.154
R4220 GND.n5124 GND.n5123 9.154
R4221 GND.n5121 GND.n5120 9.154
R4222 GND.n5118 GND.n5117 9.154
R4223 GND.n5115 GND.n5114 9.154
R4224 GND.n4768 GND.n4767 9.154
R4225 GND.n4763 GND.n4762 9.154
R4226 GND.n4760 GND.n4759 9.154
R4227 GND.n4757 GND.n4756 9.154
R4228 GND.n4754 GND.n4753 9.154
R4229 GND.n2254 GND.n2253 9.154
R4230 GND.n1290 GND.n1289 9.154
R4231 GND.n1594 GND.n1593 9.154
R4232 GND.n1597 GND.n1596 9.154
R4233 GND.n1600 GND.n1599 9.154
R4234 GND.n5968 GND.n5967 9.154
R4235 GND.n6162 GND.n6161 9.154
R4236 GND.n6317 GND.n672 9.154
R4237 GND.n1465 GND.n1464 9.154
R4238 GND.n4751 GND.n4750 9.154
R4239 GND.n490 GND.n489 9.154
R4240 GND.n6324 GND.n6323 9.154
R4241 GND.n6321 GND.n6320 9.154
R4242 GND.n6319 GND.n6318 9.154
R4243 GND.n8003 GND.n7997 9
R4244 GND.n8029 GND.n8028 9
R4245 GND.n7944 GND.n7941 9
R4246 GND.n7982 GND.n7977 9
R4247 GND.n8006 GND.n8005 9
R4248 GND.n7845 GND.n7844 9
R4249 GND.n7955 GND.n7952 9
R4250 GND.n7991 GND.n7988 9
R4251 GND.n7901 GND.n7895 9
R4252 GND.n7911 GND.n7910 9
R4253 GND.n7858 GND.n7857 9
R4254 GND.n7875 GND.n7874 9
R4255 GND.n7929 GND.n7923 9
R4256 GND.n7881 GND.n7878 9
R4257 GND.n7776 GND.n7770 9
R4258 GND.n7802 GND.n7801 9
R4259 GND.n7717 GND.n7714 9
R4260 GND.n7755 GND.n7750 9
R4261 GND.n7779 GND.n7778 9
R4262 GND.n7618 GND.n7617 9
R4263 GND.n7728 GND.n7725 9
R4264 GND.n7764 GND.n7761 9
R4265 GND.n7674 GND.n7668 9
R4266 GND.n7684 GND.n7683 9
R4267 GND.n7631 GND.n7630 9
R4268 GND.n7648 GND.n7647 9
R4269 GND.n7702 GND.n7696 9
R4270 GND.n7654 GND.n7651 9
R4271 GND.n7549 GND.n7543 9
R4272 GND.n7575 GND.n7574 9
R4273 GND.n7490 GND.n7487 9
R4274 GND.n7528 GND.n7523 9
R4275 GND.n7552 GND.n7551 9
R4276 GND.n7391 GND.n7390 9
R4277 GND.n7501 GND.n7498 9
R4278 GND.n7537 GND.n7534 9
R4279 GND.n7447 GND.n7441 9
R4280 GND.n7457 GND.n7456 9
R4281 GND.n7404 GND.n7403 9
R4282 GND.n7421 GND.n7420 9
R4283 GND.n7475 GND.n7469 9
R4284 GND.n7427 GND.n7424 9
R4285 GND.n7322 GND.n7316 9
R4286 GND.n7348 GND.n7347 9
R4287 GND.n7263 GND.n7260 9
R4288 GND.n7301 GND.n7296 9
R4289 GND.n7325 GND.n7324 9
R4290 GND.n7164 GND.n7163 9
R4291 GND.n7274 GND.n7271 9
R4292 GND.n7310 GND.n7307 9
R4293 GND.n7220 GND.n7214 9
R4294 GND.n7230 GND.n7229 9
R4295 GND.n7177 GND.n7176 9
R4296 GND.n7194 GND.n7193 9
R4297 GND.n7248 GND.n7242 9
R4298 GND.n7200 GND.n7197 9
R4299 GND.n7095 GND.n7089 9
R4300 GND.n7121 GND.n7120 9
R4301 GND.n7036 GND.n7033 9
R4302 GND.n7074 GND.n7069 9
R4303 GND.n7098 GND.n7097 9
R4304 GND.n6937 GND.n6936 9
R4305 GND.n7047 GND.n7044 9
R4306 GND.n7083 GND.n7080 9
R4307 GND.n6993 GND.n6987 9
R4308 GND.n7003 GND.n7002 9
R4309 GND.n6950 GND.n6949 9
R4310 GND.n6967 GND.n6966 9
R4311 GND.n7021 GND.n7015 9
R4312 GND.n6973 GND.n6970 9
R4313 GND.n6868 GND.n6862 9
R4314 GND.n6894 GND.n6893 9
R4315 GND.n6809 GND.n6806 9
R4316 GND.n6847 GND.n6842 9
R4317 GND.n6871 GND.n6870 9
R4318 GND.n6710 GND.n6709 9
R4319 GND.n6820 GND.n6817 9
R4320 GND.n6856 GND.n6853 9
R4321 GND.n6766 GND.n6760 9
R4322 GND.n6776 GND.n6775 9
R4323 GND.n6723 GND.n6722 9
R4324 GND.n6740 GND.n6739 9
R4325 GND.n6794 GND.n6788 9
R4326 GND.n6746 GND.n6743 9
R4327 GND.n6536 GND.n6530 9
R4328 GND.n6562 GND.n6561 9
R4329 GND.n6477 GND.n6474 9
R4330 GND.n6515 GND.n6510 9
R4331 GND.n6539 GND.n6538 9
R4332 GND.n6378 GND.n6377 9
R4333 GND.n6397 GND.n6391 9
R4334 GND.n6408 GND.n6402 9
R4335 GND.n6488 GND.n6485 9
R4336 GND.n6524 GND.n6521 9
R4337 GND.n6420 GND.n6416 9
R4338 GND.n6455 GND.n6454 9
R4339 GND.n6439 GND.n6438 9
R4340 GND.n6426 GND.n6423 9
R4341 GND.n511 GND.n510 9
R4342 GND.n522 GND.n521 9
R4343 GND.n532 GND.n531 9
R4344 GND.n593 GND.n570 9
R4345 GND.n543 GND.n542 9
R4346 GND.n554 GND.n553 9
R4347 GND.n560 GND.n559 9
R4348 GND.n1084 GND.n1083 9
R4349 GND.n1035 GND.n1034 9
R4350 GND.n1041 GND.n1040 9
R4351 GND.n1052 GND.n1051 9
R4352 GND.n1063 GND.n1062 9
R4353 GND.n1073 GND.n1072 9
R4354 GND.n1023 GND.n1022 9
R4355 GND.n886 GND.n885 9
R4356 GND.n837 GND.n836 9
R4357 GND.n847 GND.n846 9
R4358 GND.n858 GND.n857 9
R4359 GND.n869 GND.n868 9
R4360 GND.n875 GND.n874 9
R4361 GND.n826 GND.n825 9
R4362 GND.n6063 GND.n6039 9
R4363 GND.n6001 GND.n6000 9
R4364 GND.n5991 GND.n5990 9
R4365 GND.n6012 GND.n6011 9
R4366 GND.n6023 GND.n6022 9
R4367 GND.n6029 GND.n6028 9
R4368 GND.n5980 GND.n5979 9
R4369 GND.n2706 GND.n2705 9
R4370 GND.n2657 GND.n2656 9
R4371 GND.n2663 GND.n2662 9
R4372 GND.n2674 GND.n2673 9
R4373 GND.n2685 GND.n2684 9
R4374 GND.n2695 GND.n2694 9
R4375 GND.n2645 GND.n2644 9
R4376 GND.n2508 GND.n2507 9
R4377 GND.n2459 GND.n2458 9
R4378 GND.n2469 GND.n2468 9
R4379 GND.n2480 GND.n2479 9
R4380 GND.n2491 GND.n2490 9
R4381 GND.n2497 GND.n2496 9
R4382 GND.n2448 GND.n2447 9
R4383 GND.n3891 GND.n3867 9
R4384 GND.n3829 GND.n3828 9
R4385 GND.n3819 GND.n3818 9
R4386 GND.n3840 GND.n3839 9
R4387 GND.n3851 GND.n3850 9
R4388 GND.n3857 GND.n3856 9
R4389 GND.n3808 GND.n3807 9
R4390 GND.n2359 GND.n2336 9
R4391 GND.n2277 GND.n2276 9
R4392 GND.n2288 GND.n2287 9
R4393 GND.n2298 GND.n2297 9
R4394 GND.n2309 GND.n2308 9
R4395 GND.n2320 GND.n2319 9
R4396 GND.n2326 GND.n2325 9
R4397 GND.n2901 GND.n2723 9
R4398 GND.n2911 GND.n2722 9
R4399 GND.n2920 GND.n2721 9
R4400 GND.n2952 GND.n2713 9
R4401 GND.n2930 GND.n2720 9
R4402 GND.n2946 GND.n2719 9
R4403 GND.n2941 GND.n2940 9
R4404 GND.n4012 GND.n3986 9
R4405 GND.n4022 GND.n3985 9
R4406 GND.n4031 GND.n3984 9
R4407 GND.n4041 GND.n3983 9
R4408 GND.n4063 GND.n3977 9
R4409 GND.n4057 GND.n3982 9
R4410 GND.n4052 GND.n4051 9
R4411 GND.n1531 GND.n1291 9
R4412 GND.n1474 GND.n1295 9
R4413 GND.n1484 GND.n1294 9
R4414 GND.n1493 GND.n1293 9
R4415 GND.n1520 GND.n1292 9
R4416 GND.n1515 GND.n1514 9
R4417 GND.n1504 GND.n1503 9
R4418 GND.n6308 GND.n6284 9
R4419 GND.n6274 GND.n6273 9
R4420 GND.n6264 GND.n6263 9
R4421 GND.n6225 GND.n6224 9
R4422 GND.n6236 GND.n6235 9
R4423 GND.n6242 GND.n6241 9
R4424 GND.n6253 GND.n6252 9
R4425 GND.n8210 GND.n8192 9
R4426 GND.n8202 GND.n8201 9
R4427 GND.n8275 GND.n8269 9
R4428 GND.n8148 GND.n8147 9
R4429 GND.n8159 GND.n8158 9
R4430 GND.n8170 GND.n8169 9
R4431 GND.n8181 GND.n8180 9
R4432 GND.n8288 GND.n8264 9
R4433 GND.n8216 GND.n8215 9
R4434 GND.n8283 GND.n8265 9
R4435 GND.n8231 GND.n8230 9
R4436 GND.n8242 GND.n8241 9
R4437 GND.n8253 GND.n8252 9
R4438 GND.n8220 GND.n8219 9
R4439 GND.n8453 GND.n8447 9
R4440 GND.n8382 GND.n8376 9
R4441 GND.n8399 GND.n8398 9
R4442 GND.n8410 GND.n8409 9
R4443 GND.n8349 GND.n8348 9
R4444 GND.n8360 GND.n8359 9
R4445 GND.n8432 GND.n8431 9
R4446 GND.n8467 GND.n8466 9
R4447 GND.n8390 GND.n8372 9
R4448 GND.n8338 GND.n8337 9
R4449 GND.n8395 GND.n8371 9
R4450 GND.n8461 GND.n8443 9
R4451 GND.n8327 GND.n8326 9
R4452 GND.n8421 GND.n8420 9
R4453 GND.n8638 GND.n8632 9
R4454 GND.n8567 GND.n8561 9
R4455 GND.n8584 GND.n8583 9
R4456 GND.n8595 GND.n8594 9
R4457 GND.n8534 GND.n8533 9
R4458 GND.n8545 GND.n8544 9
R4459 GND.n8617 GND.n8616 9
R4460 GND.n8652 GND.n8651 9
R4461 GND.n8575 GND.n8557 9
R4462 GND.n8523 GND.n8522 9
R4463 GND.n8580 GND.n8556 9
R4464 GND.n8646 GND.n8628 9
R4465 GND.n8512 GND.n8511 9
R4466 GND.n8606 GND.n8605 9
R4467 GND.n8823 GND.n8817 9
R4468 GND.n8752 GND.n8746 9
R4469 GND.n8769 GND.n8768 9
R4470 GND.n8780 GND.n8779 9
R4471 GND.n8719 GND.n8718 9
R4472 GND.n8730 GND.n8729 9
R4473 GND.n8802 GND.n8801 9
R4474 GND.n8837 GND.n8836 9
R4475 GND.n8760 GND.n8742 9
R4476 GND.n8708 GND.n8707 9
R4477 GND.n8765 GND.n8741 9
R4478 GND.n8831 GND.n8813 9
R4479 GND.n8697 GND.n8696 9
R4480 GND.n8791 GND.n8790 9
R4481 GND.n9008 GND.n9002 9
R4482 GND.n8937 GND.n8931 9
R4483 GND.n8954 GND.n8953 9
R4484 GND.n8965 GND.n8964 9
R4485 GND.n8904 GND.n8903 9
R4486 GND.n8915 GND.n8914 9
R4487 GND.n8987 GND.n8986 9
R4488 GND.n9022 GND.n9021 9
R4489 GND.n8945 GND.n8927 9
R4490 GND.n8893 GND.n8892 9
R4491 GND.n8950 GND.n8926 9
R4492 GND.n9016 GND.n8998 9
R4493 GND.n8882 GND.n8881 9
R4494 GND.n8976 GND.n8975 9
R4495 GND.n9193 GND.n9187 9
R4496 GND.n9122 GND.n9116 9
R4497 GND.n9139 GND.n9138 9
R4498 GND.n9150 GND.n9149 9
R4499 GND.n9089 GND.n9088 9
R4500 GND.n9100 GND.n9099 9
R4501 GND.n9172 GND.n9171 9
R4502 GND.n9207 GND.n9206 9
R4503 GND.n9130 GND.n9112 9
R4504 GND.n9078 GND.n9077 9
R4505 GND.n9135 GND.n9111 9
R4506 GND.n9201 GND.n9183 9
R4507 GND.n9067 GND.n9066 9
R4508 GND.n9161 GND.n9160 9
R4509 GND.n154 GND.n148 9
R4510 GND.n83 GND.n77 9
R4511 GND.n100 GND.n99 9
R4512 GND.n111 GND.n110 9
R4513 GND.n50 GND.n49 9
R4514 GND.n61 GND.n60 9
R4515 GND.n133 GND.n132 9
R4516 GND.n168 GND.n167 9
R4517 GND.n91 GND.n73 9
R4518 GND.n39 GND.n38 9
R4519 GND.n96 GND.n72 9
R4520 GND.n162 GND.n144 9
R4521 GND.n28 GND.n27 9
R4522 GND.n122 GND.n121 9
R4523 GND.n6130 GND.n6129 8.764
R4524 GND.n1276 GND.n1275 8.764
R4525 GND.n3958 GND.n3957 8.764
R4526 GND.n3795 GND.n3794 8.764
R4527 GND.n2271 GND.n2270 8.764
R4528 GND.n4306 GND.n4305 8.764
R4529 GND.n505 GND.n504 8.764
R4530 GND.n657 GND.n656 8.764
R4531 GND.n1831 GND.n1828 8.522
R4532 GND.n4404 GND.n4403 8.522
R4533 GND.n1777 GND.n1774 8.522
R4534 GND.n1790 GND.n1787 8.522
R4535 GND.n1803 GND.n1800 8.522
R4536 GND.n1816 GND.n1813 8.522
R4537 GND.n5870 GND.n5867 8.522
R4538 GND.n3205 GND.n3202 8.522
R4539 GND.n3575 GND.n3574 8.522
R4540 GND.n3614 GND.n3611 8.522
R4541 GND.n4136 GND.n4133 8.522
R4542 GND.n2731 GND.n2728 8.522
R4543 GND.n1096 GND.n1093 8.522
R4544 GND.n1303 GND.n1300 8.522
R4545 GND.n5917 GND.n5914 8.282
R4546 GND.n5147 GND.n5144 8.282
R4547 GND.n563 GND.n562 7.99
R4548 GND.n1030 GND.n1029 7.99
R4549 GND.n878 GND.n877 7.99
R4550 GND.n2652 GND.n2651 7.99
R4551 GND.n2500 GND.n2499 7.99
R4552 GND.n2329 GND.n2328 7.99
R4553 GND.n2717 GND.n2716 7.99
R4554 GND.n3980 GND.n3979 7.99
R4555 GND.n1525 GND.n1524 7.99
R4556 GND.n6231 GND.n6230 7.99
R4557 GND.n6032 GND.n6031 7.99
R4558 GND.n3860 GND.n3859 7.99
R4559 GND.n4403 GND.n4402 7.027
R4560 GND.n3780 GND.n3779 6.793
R4561 GND.n2437 GND.n2436 6.793
R4562 GND.n1610 GND.n1609 6.716
R4563 GND.n5713 GND.n5712 6.716
R4564 GND.n1999 GND.n1998 6.716
R4565 GND.n1842 GND.n1841 6.716
R4566 GND.n5309 GND.n5308 6.716
R4567 GND.n5152 GND.n5151 6.716
R4568 GND.n5153 GND.n5152 6.716
R4569 GND.n1843 GND.n1842 6.716
R4570 GND.n4559 GND.n4558 6.716
R4571 GND.n4930 GND.n4929 6.716
R4572 GND.n4773 GND.n4772 6.716
R4573 GND.n4774 GND.n4773 6.716
R4574 GND.n4929 GND.n4928 6.716
R4575 GND.n4558 GND.n4557 6.716
R4576 GND.n5308 GND.n5307 6.716
R4577 GND.n1998 GND.n1997 6.716
R4578 GND.n5712 GND.n5711 6.716
R4579 GND.n3624 GND.n3623 6.716
R4580 GND.n4287 GND.n4286 6.716
R4581 GND.n3623 GND.n3622 6.716
R4582 GND.n4288 GND.n4287 6.716
R4583 GND.n1106 GND.n1105 6.716
R4584 GND.n666 GND.n665 6.716
R4585 GND.n3033 GND.n3032 6.716
R4586 GND.n2883 GND.n2882 6.716
R4587 GND.n2882 GND.n2881 6.716
R4588 GND.n3032 GND.n3031 6.716
R4589 GND.n1105 GND.n1104 6.716
R4590 GND.n665 GND.n664 6.716
R4591 GND.n1609 GND.n1608 6.716
R4592 GND.n5790 GND.n5789 6.023
R4593 GND.n5782 GND.n5781 6.023
R4594 GND.n5610 GND.n5609 6.023
R4595 GND.n5602 GND.n5601 6.023
R4596 GND.n1916 GND.n1915 6.023
R4597 GND.n1924 GND.n1923 6.023
R4598 GND.n2096 GND.n2095 6.023
R4599 GND.n2104 GND.n2103 6.023
R4600 GND.n5226 GND.n5225 6.023
R4601 GND.n5234 GND.n5233 6.023
R4602 GND.n5406 GND.n5405 6.023
R4603 GND.n5414 GND.n5413 6.023
R4604 GND.n4476 GND.n4475 6.023
R4605 GND.n4484 GND.n4483 6.023
R4606 GND.n4658 GND.n4657 6.023
R4607 GND.n4666 GND.n4665 6.023
R4608 GND.n4847 GND.n4846 6.023
R4609 GND.n4855 GND.n4854 6.023
R4610 GND.n5027 GND.n5026 6.023
R4611 GND.n5035 GND.n5034 6.023
R4612 GND.n3492 GND.n3491 6.023
R4613 GND.n3483 GND.n3482 6.023
R4614 GND.n3308 GND.n3307 6.023
R4615 GND.n3300 GND.n3299 6.023
R4616 GND.n3701 GND.n3700 6.023
R4617 GND.n3693 GND.n3692 6.023
R4618 GND.n4205 GND.n4204 6.023
R4619 GND.n4213 GND.n4212 6.023
R4620 GND.n3111 GND.n3110 6.023
R4621 GND.n3103 GND.n3102 6.023
R4622 GND.n2800 GND.n2799 6.023
R4623 GND.n2808 GND.n2807 6.023
R4624 GND.n5899 GND.n5896 6.023
R4625 GND.n1183 GND.n1182 6.023
R4626 GND.n1175 GND.n1174 6.023
R4627 GND.n738 GND.n737 6.023
R4628 GND.n746 GND.n745 6.023
R4629 GND.n5509 GND.n5506 6.023
R4630 GND.n1688 GND.n1687 6.023
R4631 GND.n1680 GND.n1679 6.023
R4632 GND.n1372 GND.n1371 6.023
R4633 GND.n1380 GND.n1379 6.023
R4634 GND.n5802 GND.n5801 5.27
R4635 GND.n5770 GND.n5769 5.27
R4636 GND.n5622 GND.n5621 5.27
R4637 GND.n5590 GND.n5589 5.27
R4638 GND.n1904 GND.n1903 5.27
R4639 GND.n1936 GND.n1935 5.27
R4640 GND.n2084 GND.n2083 5.27
R4641 GND.n2116 GND.n2115 5.27
R4642 GND.n5214 GND.n5213 5.27
R4643 GND.n5246 GND.n5245 5.27
R4644 GND.n5394 GND.n5393 5.27
R4645 GND.n5426 GND.n5425 5.27
R4646 GND.n4464 GND.n4463 5.27
R4647 GND.n4496 GND.n4495 5.27
R4648 GND.n4645 GND.n4644 5.27
R4649 GND.n4679 GND.n4678 5.27
R4650 GND.n4835 GND.n4834 5.27
R4651 GND.n4867 GND.n4866 5.27
R4652 GND.n5015 GND.n5014 5.27
R4653 GND.n5047 GND.n5046 5.27
R4654 GND.n3504 GND.n3503 5.27
R4655 GND.n3470 GND.n3469 5.27
R4656 GND.n3320 GND.n3319 5.27
R4657 GND.n3288 GND.n3287 5.27
R4658 GND.n3713 GND.n3712 5.27
R4659 GND.n3681 GND.n3680 5.27
R4660 GND.n4193 GND.n4192 5.27
R4661 GND.n4225 GND.n4224 5.27
R4662 GND.n3123 GND.n3122 5.27
R4663 GND.n3091 GND.n3090 5.27
R4664 GND.n2788 GND.n2787 5.27
R4665 GND.n2820 GND.n2819 5.27
R4666 GND.n1195 GND.n1194 5.27
R4667 GND.n1163 GND.n1162 5.27
R4668 GND.n726 GND.n725 5.27
R4669 GND.n758 GND.n757 5.27
R4670 GND.n1700 GND.n1699 5.27
R4671 GND.n1668 GND.n1667 5.27
R4672 GND.n1360 GND.n1359 5.27
R4673 GND.n1392 GND.n1391 5.27
R4674 GND.n5873 GND.n5872 4.894
R4675 GND.n5872 GND.n5866 4.894
R4676 GND.n5715 GND.n5710 4.894
R4677 GND.n5687 GND.n5682 4.894
R4678 GND.n1833 GND.n1827 4.894
R4679 GND.n1834 GND.n1833 4.894
R4680 GND.n1819 GND.n1818 4.894
R4681 GND.n1818 GND.n1812 4.894
R4682 GND.n2001 GND.n1996 4.894
R4683 GND.n2029 GND.n2024 4.894
R4684 GND.n1846 GND.n1840 4.894
R4685 GND.n1847 GND.n1846 4.894
R4686 GND.n1806 GND.n1805 4.894
R4687 GND.n1805 GND.n1799 4.894
R4688 GND.n5311 GND.n5306 4.894
R4689 GND.n5339 GND.n5334 4.894
R4690 GND.n5156 GND.n5150 4.894
R4691 GND.n5157 GND.n5156 4.894
R4692 GND.n1793 GND.n1792 4.894
R4693 GND.n1792 GND.n1786 4.894
R4694 GND.n4561 GND.n4556 4.894
R4695 GND.n4589 GND.n4584 4.894
R4696 GND.n4406 GND.n4399 4.894
R4697 GND.n4407 GND.n4406 4.894
R4698 GND.n1780 GND.n1779 4.894
R4699 GND.n1779 GND.n1773 4.894
R4700 GND.n4932 GND.n4927 4.894
R4701 GND.n4960 GND.n4955 4.894
R4702 GND.n4777 GND.n4771 4.894
R4703 GND.n4778 GND.n4777 4.894
R4704 GND.n3578 GND.n3577 4.894
R4705 GND.n3577 GND.n3571 4.894
R4706 GND.n3413 GND.n3408 4.894
R4707 GND.n3385 GND.n3380 4.894
R4708 GND.n3207 GND.n3201 4.894
R4709 GND.n3208 GND.n3207 4.894
R4710 GND.n3617 GND.n3616 4.894
R4711 GND.n3616 GND.n3610 4.894
R4712 GND.n3626 GND.n3621 4.894
R4713 GND.n4138 GND.n4132 4.894
R4714 GND.n4290 GND.n4285 4.894
R4715 GND.n3188 GND.n3183 4.894
R4716 GND.n3036 GND.n3030 4.894
R4717 GND.n2733 GND.n2727 4.894
R4718 GND.n2885 GND.n2880 4.894
R4719 GND.n1099 GND.n1098 4.894
R4720 GND.n1098 GND.n1092 4.894
R4721 GND.n1108 GND.n1103 4.894
R4722 GND.n6155 GND.n6150 4.894
R4723 GND.n669 GND.n663 4.894
R4724 GND.n670 GND.n669 4.894
R4725 GND.n1765 GND.n1760 4.894
R4726 GND.n1613 GND.n1607 4.894
R4727 GND.n1305 GND.n1299 4.894
R4728 GND.n1458 GND.n1453 4.894
R4729 GND.n6131 GND.n6130 4.65
R4730 GND.n1277 GND.n1276 4.65
R4731 GND.n3959 GND.n3958 4.65
R4732 GND.n3796 GND.n3795 4.65
R4733 GND.n2009 GND.n2008 4.65
R4734 GND.n2012 GND.n2011 4.65
R4735 GND.n2015 GND.n2014 4.65
R4736 GND.n2018 GND.n2017 4.65
R4737 GND.n1822 GND.n1821 4.65
R4738 GND.n2181 GND.n2180 4.65
R4739 GND.n5319 GND.n5318 4.65
R4740 GND.n5322 GND.n5321 4.65
R4741 GND.n5325 GND.n5324 4.65
R4742 GND.n5328 GND.n5327 4.65
R4743 GND.n1809 GND.n1808 4.65
R4744 GND.n5491 GND.n5490 4.65
R4745 GND.n4569 GND.n4568 4.65
R4746 GND.n4572 GND.n4571 4.65
R4747 GND.n4575 GND.n4574 4.65
R4748 GND.n4578 GND.n4577 4.65
R4749 GND.n1796 GND.n1795 4.65
R4750 GND.n4747 GND.n4746 4.65
R4751 GND.n4940 GND.n4939 4.65
R4752 GND.n4943 GND.n4942 4.65
R4753 GND.n4946 GND.n4945 4.65
R4754 GND.n4949 GND.n4948 4.65
R4755 GND.n1783 GND.n1782 4.65
R4756 GND.n5112 GND.n5111 4.65
R4757 GND.n3402 GND.n3401 4.65
R4758 GND.n3399 GND.n3398 4.65
R4759 GND.n3396 GND.n3395 4.65
R4760 GND.n3393 GND.n3392 4.65
R4761 GND.n3581 GND.n3580 4.65
R4762 GND.n3229 GND.n3228 4.65
R4763 GND.n5704 GND.n5703 4.65
R4764 GND.n5701 GND.n5700 4.65
R4765 GND.n5698 GND.n5697 4.65
R4766 GND.n5695 GND.n5694 4.65
R4767 GND.n5876 GND.n5875 4.65
R4768 GND.n5531 GND.n5530 4.65
R4769 GND.n2272 GND.n2271 4.65
R4770 GND.n4307 GND.n4306 4.65
R4771 GND.n3976 GND.n3975 4.65
R4772 GND.n4296 GND.n2441 4.65
R4773 GND.n3973 GND.n3972 4.65
R4774 GND.n3970 GND.n3969 4.65
R4775 GND.n3778 GND.n3777 4.65
R4776 GND.n4126 GND.n4125 4.65
R4777 GND.n3021 GND.n3020 4.65
R4778 GND.n2893 GND.n2892 4.65
R4779 GND.n3015 GND.n3014 4.65
R4780 GND.n3018 GND.n3017 4.65
R4781 GND.n3024 GND.n3023 4.65
R4782 GND.n3196 GND.n3195 4.65
R4783 GND.n3199 GND.n3198 4.65
R4784 GND.n3799 GND.n3798 4.65
R4785 GND.n3793 GND.n3792 4.65
R4786 GND.n3786 GND.n3785 4.65
R4787 GND.n3783 GND.n3782 4.65
R4788 GND.n3608 GND.n3607 4.65
R4789 GND.n3605 GND.n3604 4.65
R4790 GND.n3602 GND.n3601 4.65
R4791 GND.n3599 GND.n3598 4.65
R4792 GND.n3595 GND.n3594 4.65
R4793 GND.n3590 GND.n3589 4.65
R4794 GND.n3587 GND.n3586 4.65
R4795 GND.n3584 GND.n3583 4.65
R4796 GND.n1825 GND.n1824 4.65
R4797 GND.n5882 GND.n5881 4.65
R4798 GND.n5885 GND.n5884 4.65
R4799 GND.n5888 GND.n5887 4.65
R4800 GND.n5891 GND.n5890 4.65
R4801 GND.n5894 GND.n5893 4.65
R4802 GND.n5900 GND.n5899 4.65
R4803 GND.n5903 GND.n5902 4.65
R4804 GND.n5906 GND.n5905 4.65
R4805 GND.n5909 GND.n5908 4.65
R4806 GND.n5912 GND.n5911 4.65
R4807 GND.n5918 GND.n5917 4.65
R4808 GND.n5921 GND.n5920 4.65
R4809 GND.n5924 GND.n5923 4.65
R4810 GND.n5927 GND.n5926 4.65
R4811 GND.n5930 GND.n5929 4.65
R4812 GND.n5936 GND.n5935 4.65
R4813 GND.n5939 GND.n5938 4.65
R4814 GND.n5942 GND.n5941 4.65
R4815 GND.n5945 GND.n5944 4.65
R4816 GND.n5948 GND.n5947 4.65
R4817 GND.n5954 GND.n5953 4.65
R4818 GND.n5957 GND.n5956 4.65
R4819 GND.n5960 GND.n5959 4.65
R4820 GND.n5963 GND.n5962 4.65
R4821 GND.n5966 GND.n5965 4.65
R4822 GND.n5974 GND.n5973 4.65
R4823 GND.n1286 GND.n1285 4.65
R4824 GND.n1274 GND.n1273 4.65
R4825 GND.n1265 GND.n1264 4.65
R4826 GND.n1263 GND.n1261 4.65
R4827 GND.n6142 GND.n6141 4.65
R4828 GND.n6145 GND.n6144 4.65
R4829 GND.n6148 GND.n6147 4.65
R4830 GND.n1260 GND.n1259 4.65
R4831 GND.n2252 GND.n2251 4.65
R4832 GND.n2425 GND.n2424 4.65
R4833 GND.n2438 GND.n2435 4.65
R4834 GND.n2434 GND.n2433 4.65
R4835 GND.n2431 GND.n2430 4.65
R4836 GND.n2428 GND.n2427 4.65
R4837 GND.n3212 GND.n3211 4.65
R4838 GND.n3226 GND.n3225 4.65
R4839 GND.n3221 GND.n3220 4.65
R4840 GND.n3218 GND.n3217 4.65
R4841 GND.n3215 GND.n3214 4.65
R4842 GND.n1838 GND.n1837 4.65
R4843 GND.n5528 GND.n5527 4.65
R4844 GND.n5523 GND.n5522 4.65
R4845 GND.n5520 GND.n5519 4.65
R4846 GND.n5517 GND.n5516 4.65
R4847 GND.n5514 GND.n5513 4.65
R4848 GND.n5510 GND.n5509 4.65
R4849 GND.n5505 GND.n5504 4.65
R4850 GND.n5502 GND.n5501 4.65
R4851 GND.n5498 GND.n5497 4.65
R4852 GND.n5495 GND.n5494 4.65
R4853 GND.n5148 GND.n5147 4.65
R4854 GND.n5143 GND.n5142 4.65
R4855 GND.n5140 GND.n5139 4.65
R4856 GND.n5137 GND.n5136 4.65
R4857 GND.n5134 GND.n5133 4.65
R4858 GND.n5130 GND.n5129 4.65
R4859 GND.n5125 GND.n5124 4.65
R4860 GND.n5122 GND.n5121 4.65
R4861 GND.n5119 GND.n5118 4.65
R4862 GND.n5116 GND.n5115 4.65
R4863 GND.n4769 GND.n4768 4.65
R4864 GND.n4764 GND.n4763 4.65
R4865 GND.n4761 GND.n4760 4.65
R4866 GND.n4758 GND.n4757 4.65
R4867 GND.n4755 GND.n4754 4.65
R4868 GND.n1595 GND.n1594 4.65
R4869 GND.n1598 GND.n1597 4.65
R4870 GND.n1601 GND.n1600 4.65
R4871 GND.n5969 GND.n5968 4.65
R4872 GND.n1592 GND.n1290 4.65
R4873 GND.n6163 GND.n6162 4.65
R4874 GND.n506 GND.n505 4.65
R4875 GND.n6317 GND.n6316 4.65
R4876 GND.n6326 GND.n657 4.65
R4877 GND.n1466 GND.n1465 4.65
R4878 GND.n4752 GND.n4751 4.65
R4879 GND.n491 GND.n490 4.65
R4880 GND.n6325 GND.n6324 4.65
R4881 GND.n3802 GND.n3801 4.589
R4882 GND.n3790 GND.n3789 4.589
R4883 GND.n7970 GND.n7969 4.574
R4884 GND.n7964 GND.n7962 4.574
R4885 GND.n7743 GND.n7742 4.574
R4886 GND.n7737 GND.n7735 4.574
R4887 GND.n7516 GND.n7515 4.574
R4888 GND.n7510 GND.n7508 4.574
R4889 GND.n7289 GND.n7288 4.574
R4890 GND.n7283 GND.n7281 4.574
R4891 GND.n7062 GND.n7061 4.574
R4892 GND.n7056 GND.n7054 4.574
R4893 GND.n6835 GND.n6834 4.574
R4894 GND.n6829 GND.n6827 4.574
R4895 GND.n6503 GND.n6502 4.574
R4896 GND.n6497 GND.n6495 4.574
R4897 GND.n566 GND.n565 4.574
R4898 GND.n1032 GND.n1031 4.574
R4899 GND.n881 GND.n880 4.574
R4900 GND.n6035 GND.n6034 4.574
R4901 GND.n2654 GND.n2653 4.574
R4902 GND.n2503 GND.n2502 4.574
R4903 GND.n3863 GND.n3862 4.574
R4904 GND.n2332 GND.n2331 4.574
R4905 GND.n2948 GND.n2718 4.574
R4906 GND.n4059 GND.n3981 4.574
R4907 GND.n1527 GND.n1526 4.574
R4908 GND.n6233 GND.n6232 4.574
R4909 GND.n8206 GND.n8195 4.574
R4910 GND.n8279 GND.n8268 4.574
R4911 GND.n8386 GND.n8375 4.574
R4912 GND.n8457 GND.n8446 4.574
R4913 GND.n8571 GND.n8560 4.574
R4914 GND.n8642 GND.n8631 4.574
R4915 GND.n8756 GND.n8745 4.574
R4916 GND.n8827 GND.n8816 4.574
R4917 GND.n8941 GND.n8930 4.574
R4918 GND.n9012 GND.n9001 4.574
R4919 GND.n9126 GND.n9115 4.574
R4920 GND.n9197 GND.n9186 4.574
R4921 GND.n87 GND.n76 4.574
R4922 GND.n158 GND.n147 4.574
R4923 GND.n5814 GND.n5813 4.517
R4924 GND.n5758 GND.n5757 4.517
R4925 GND.n5634 GND.n5633 4.517
R4926 GND.n5578 GND.n5577 4.517
R4927 GND.n1892 GND.n1891 4.517
R4928 GND.n1948 GND.n1947 4.517
R4929 GND.n2072 GND.n2071 4.517
R4930 GND.n2128 GND.n2127 4.517
R4931 GND.n5202 GND.n5201 4.517
R4932 GND.n5258 GND.n5257 4.517
R4933 GND.n5382 GND.n5381 4.517
R4934 GND.n5438 GND.n5437 4.517
R4935 GND.n4452 GND.n4451 4.517
R4936 GND.n4508 GND.n4507 4.517
R4937 GND.n4633 GND.n4632 4.517
R4938 GND.n4692 GND.n4691 4.517
R4939 GND.n4823 GND.n4822 4.517
R4940 GND.n4879 GND.n4878 4.517
R4941 GND.n5003 GND.n5002 4.517
R4942 GND.n5059 GND.n5058 4.517
R4943 GND.n3517 GND.n3516 4.517
R4944 GND.n3458 GND.n3457 4.517
R4945 GND.n3332 GND.n3331 4.517
R4946 GND.n3276 GND.n3275 4.517
R4947 GND.n3725 GND.n3724 4.517
R4948 GND.n3669 GND.n3668 4.517
R4949 GND.n4181 GND.n4180 4.517
R4950 GND.n4237 GND.n4236 4.517
R4951 GND.n3135 GND.n3134 4.517
R4952 GND.n3079 GND.n3078 4.517
R4953 GND.n2776 GND.n2775 4.517
R4954 GND.n2832 GND.n2831 4.517
R4955 GND.n1207 GND.n1206 4.517
R4956 GND.n1151 GND.n1150 4.517
R4957 GND.n714 GND.n713 4.517
R4958 GND.n770 GND.n769 4.517
R4959 GND.n1712 GND.n1711 4.517
R4960 GND.n1656 GND.n1655 4.517
R4961 GND.n1348 GND.n1347 4.517
R4962 GND.n1404 GND.n1403 4.517
R4963 GND.n5855 GND.n5850 4.141
R4964 GND.n5727 GND.n5722 4.141
R4965 GND.n5675 GND.n5670 4.141
R4966 GND.n5547 GND.n5541 4.141
R4967 GND.n1861 GND.n1856 4.141
R4968 GND.n1989 GND.n1984 4.141
R4969 GND.n2041 GND.n2036 4.141
R4970 GND.n2169 GND.n2164 4.141
R4971 GND.n5171 GND.n5166 4.141
R4972 GND.n5299 GND.n5294 4.141
R4973 GND.n5351 GND.n5346 4.141
R4974 GND.n5479 GND.n5474 4.141
R4975 GND.n4421 GND.n4416 4.141
R4976 GND.n4549 GND.n4544 4.141
R4977 GND.n4601 GND.n4596 4.141
R4978 GND.n4735 GND.n4729 4.141
R4979 GND.n4792 GND.n4787 4.141
R4980 GND.n4920 GND.n4915 4.141
R4981 GND.n4972 GND.n4967 4.141
R4982 GND.n5100 GND.n5095 4.141
R4983 GND.n3560 GND.n3554 4.141
R4984 GND.n3426 GND.n3420 4.141
R4985 GND.n3373 GND.n3368 4.141
R4986 GND.n3245 GND.n3239 4.141
R4987 GND.n3766 GND.n3761 4.141
R4988 GND.n3638 GND.n3633 4.141
R4989 GND.n4150 GND.n4145 4.141
R4990 GND.n4278 GND.n4273 4.141
R4991 GND.n3176 GND.n3171 4.141
R4992 GND.n3048 GND.n3043 4.141
R4993 GND.n2745 GND.n2740 4.141
R4994 GND.n2873 GND.n2868 4.141
R4995 GND.n1248 GND.n1243 4.141
R4996 GND.n1120 GND.n1115 4.141
R4997 GND.n683 GND.n678 4.141
R4998 GND.n811 GND.n806 4.141
R4999 GND.n1753 GND.n1748 4.141
R5000 GND.n1625 GND.n1620 4.141
R5001 GND.n1317 GND.n1312 4.141
R5002 GND.n1446 GND.n1440 4.141
R5003 GND.n5826 GND.n5825 3.764
R5004 GND.n5746 GND.n5745 3.764
R5005 GND.n5646 GND.n5645 3.764
R5006 GND.n5566 GND.n5565 3.764
R5007 GND.n1880 GND.n1879 3.764
R5008 GND.n1960 GND.n1959 3.764
R5009 GND.n2060 GND.n2059 3.764
R5010 GND.n2140 GND.n2139 3.764
R5011 GND.n5190 GND.n5189 3.764
R5012 GND.n5270 GND.n5269 3.764
R5013 GND.n5370 GND.n5369 3.764
R5014 GND.n5450 GND.n5449 3.764
R5015 GND.n4440 GND.n4439 3.764
R5016 GND.n4520 GND.n4519 3.764
R5017 GND.n4620 GND.n4619 3.764
R5018 GND.n4704 GND.n4703 3.764
R5019 GND.n4811 GND.n4810 3.764
R5020 GND.n4891 GND.n4890 3.764
R5021 GND.n4991 GND.n4990 3.764
R5022 GND.n5071 GND.n5070 3.764
R5023 GND.n3529 GND.n3528 3.764
R5024 GND.n3445 GND.n3444 3.764
R5025 GND.n3344 GND.n3343 3.764
R5026 GND.n3264 GND.n3263 3.764
R5027 GND.n3737 GND.n3736 3.764
R5028 GND.n3657 GND.n3656 3.764
R5029 GND.n4169 GND.n4168 3.764
R5030 GND.n4249 GND.n4248 3.764
R5031 GND.n3147 GND.n3146 3.764
R5032 GND.n3067 GND.n3066 3.764
R5033 GND.n2764 GND.n2763 3.764
R5034 GND.n2844 GND.n2843 3.764
R5035 GND.n5881 GND.n5878 3.764
R5036 GND.n1219 GND.n1218 3.764
R5037 GND.n1139 GND.n1138 3.764
R5038 GND.n702 GND.n701 3.764
R5039 GND.n782 GND.n781 3.764
R5040 GND.n5527 GND.n5524 3.764
R5041 GND.n1724 GND.n1723 3.764
R5042 GND.n1644 GND.n1643 3.764
R5043 GND.n1336 GND.n1335 3.764
R5044 GND.n1416 GND.n1415 3.764
R5045 GND.n6322 GND.n6319 3.669
R5046 GND.n2257 GND.n2254 3.588
R5047 GND.n2257 GND.n2256 3.549
R5048 GND.n6322 GND.n6321 3.538
R5049 GND.n1684 GND.n1683 3.396
R5050 GND.n1384 GND.n1383 3.396
R5051 GND.n5786 GND.n5785 3.396
R5052 GND.n5606 GND.n5605 3.396
R5053 GND.n1928 GND.n1927 3.396
R5054 GND.n2108 GND.n2107 3.396
R5055 GND.n5238 GND.n5237 3.396
R5056 GND.n5418 GND.n5417 3.396
R5057 GND.n4488 GND.n4487 3.396
R5058 GND.n4859 GND.n4858 3.396
R5059 GND.n5039 GND.n5038 3.396
R5060 GND.n3304 GND.n3303 3.396
R5061 GND.n3697 GND.n3696 3.396
R5062 GND.n4217 GND.n4216 3.396
R5063 GND.n1179 GND.n1178 3.396
R5064 GND.n750 GND.n749 3.396
R5065 GND.n3107 GND.n3106 3.396
R5066 GND.n2812 GND.n2811 3.396
R5067 GND.n7969 GND.n7967 3.388
R5068 GND.n7962 GND.n7960 3.388
R5069 GND.n7742 GND.n7740 3.388
R5070 GND.n7735 GND.n7733 3.388
R5071 GND.n7515 GND.n7513 3.388
R5072 GND.n7508 GND.n7506 3.388
R5073 GND.n7288 GND.n7286 3.388
R5074 GND.n7281 GND.n7279 3.388
R5075 GND.n7061 GND.n7059 3.388
R5076 GND.n7054 GND.n7052 3.388
R5077 GND.n6834 GND.n6832 3.388
R5078 GND.n6827 GND.n6825 3.388
R5079 GND.n6502 GND.n6500 3.388
R5080 GND.n6495 GND.n6493 3.388
R5081 GND.n6232 GND.n6229 3.388
R5082 GND.n565 GND.n564 3.388
R5083 GND.n6034 GND.n6033 3.388
R5084 GND.n1031 GND.n1027 3.388
R5085 GND.n880 GND.n879 3.388
R5086 GND.n3862 GND.n3861 3.388
R5087 GND.n2653 GND.n2649 3.388
R5088 GND.n2502 GND.n2501 3.388
R5089 GND.n5843 GND.n5838 3.388
R5090 GND.n5739 GND.n5734 3.388
R5091 GND.n5663 GND.n5658 3.388
R5092 GND.n5559 GND.n5554 3.388
R5093 GND.n1873 GND.n1868 3.388
R5094 GND.n1977 GND.n1972 3.388
R5095 GND.n2053 GND.n2048 3.388
R5096 GND.n2157 GND.n2152 3.388
R5097 GND.n5183 GND.n5178 3.388
R5098 GND.n5287 GND.n5282 3.388
R5099 GND.n5363 GND.n5358 3.388
R5100 GND.n5467 GND.n5462 3.388
R5101 GND.n4433 GND.n4428 3.388
R5102 GND.n4537 GND.n4532 3.388
R5103 GND.n4613 GND.n4608 3.388
R5104 GND.n4722 GND.n4717 3.388
R5105 GND.n4804 GND.n4799 3.388
R5106 GND.n4908 GND.n4903 3.388
R5107 GND.n4984 GND.n4979 3.388
R5108 GND.n5088 GND.n5083 3.388
R5109 GND.n3547 GND.n3542 3.388
R5110 GND.n3438 GND.n3433 3.388
R5111 GND.n3361 GND.n3356 3.388
R5112 GND.n3257 GND.n3252 3.388
R5113 GND.n3981 GND.n3978 3.388
R5114 GND.n2331 GND.n2330 3.388
R5115 GND.n2718 GND.n2714 3.388
R5116 GND.n3754 GND.n3749 3.388
R5117 GND.n3650 GND.n3645 3.388
R5118 GND.n4162 GND.n4157 3.388
R5119 GND.n4266 GND.n4261 3.388
R5120 GND.n3164 GND.n3159 3.388
R5121 GND.n3060 GND.n3055 3.388
R5122 GND.n2757 GND.n2752 3.388
R5123 GND.n2861 GND.n2856 3.388
R5124 GND.n1236 GND.n1231 3.388
R5125 GND.n1132 GND.n1127 3.388
R5126 GND.n695 GND.n690 3.388
R5127 GND.n799 GND.n794 3.388
R5128 GND.n1741 GND.n1736 3.388
R5129 GND.n1637 GND.n1632 3.388
R5130 GND.n1329 GND.n1324 3.388
R5131 GND.n1433 GND.n1428 3.388
R5132 GND.n1526 GND.n1522 3.388
R5133 GND.n8268 GND.n8267 3.388
R5134 GND.n8195 GND.n8194 3.388
R5135 GND.n8375 GND.n8374 3.388
R5136 GND.n8446 GND.n8445 3.388
R5137 GND.n8560 GND.n8559 3.388
R5138 GND.n8631 GND.n8630 3.388
R5139 GND.n8745 GND.n8744 3.388
R5140 GND.n8816 GND.n8815 3.388
R5141 GND.n8930 GND.n8929 3.388
R5142 GND.n9001 GND.n9000 3.388
R5143 GND.n9115 GND.n9114 3.388
R5144 GND.n9186 GND.n9185 3.388
R5145 GND.n76 GND.n75 3.388
R5146 GND.n147 GND.n146 3.388
R5147 GND.n7937 GND.t1 3.326
R5148 GND.n7947 GND.t47 3.326
R5149 GND.n7710 GND.t75 3.326
R5150 GND.n7720 GND.t69 3.326
R5151 GND.n7483 GND.t45 3.326
R5152 GND.n7493 GND.t83 3.326
R5153 GND.n7256 GND.t65 3.326
R5154 GND.n7266 GND.t53 3.326
R5155 GND.n7029 GND.t5 3.326
R5156 GND.n7039 GND.t89 3.326
R5157 GND.n6802 GND.t61 3.326
R5158 GND.n6812 GND.t71 3.326
R5159 GND.n6470 GND.t67 3.326
R5160 GND.n6480 GND.t63 3.326
R5161 GND.n6230 GND.t20 3.326
R5162 GND.n562 GND.t19 3.326
R5163 GND.n1029 GND.n1028 3.326
R5164 GND.n1029 GND.t27 3.326
R5165 GND.n877 GND.t28 3.326
R5166 GND.n2651 GND.n2650 3.326
R5167 GND.n2651 GND.t15 3.326
R5168 GND.n2499 GND.t16 3.326
R5169 GND.n3979 GND.t24 3.326
R5170 GND.n2328 GND.t23 3.326
R5171 GND.n2716 GND.n2715 3.326
R5172 GND.n1524 GND.n1523 3.326
R5173 GND.n8270 GND.t3 3.326
R5174 GND.n8196 GND.t7 3.326
R5175 GND.n8377 GND.t51 3.326
R5176 GND.n8448 GND.t73 3.326
R5177 GND.n8562 GND.t85 3.326
R5178 GND.n8633 GND.t81 3.326
R5179 GND.n8747 GND.t59 3.326
R5180 GND.n8818 GND.t55 3.326
R5181 GND.n8932 GND.t49 3.326
R5182 GND.n9003 GND.t91 3.326
R5183 GND.n9117 GND.t77 3.326
R5184 GND.n9188 GND.t57 3.326
R5185 GND.n78 GND.t79 3.326
R5186 GND.n149 GND.t87 3.326
R5187 GND.n1691 GND.n1690 3.324
R5188 GND.n1375 GND.n1374 3.324
R5189 GND.n5793 GND.n5792 3.324
R5190 GND.n5613 GND.n5612 3.324
R5191 GND.n1919 GND.n1918 3.324
R5192 GND.n2099 GND.n2098 3.324
R5193 GND.n5229 GND.n5228 3.324
R5194 GND.n5409 GND.n5408 3.324
R5195 GND.n4479 GND.n4478 3.324
R5196 GND.n4670 GND.n4669 3.324
R5197 GND.n4661 GND.n4660 3.324
R5198 GND.n4850 GND.n4849 3.324
R5199 GND.n5030 GND.n5029 3.324
R5200 GND.n3487 GND.n3486 3.324
R5201 GND.n3311 GND.n3310 3.324
R5202 GND.n3495 GND.n3494 3.324
R5203 GND.n3704 GND.n3703 3.324
R5204 GND.n4208 GND.n4207 3.324
R5205 GND.n1186 GND.n1185 3.324
R5206 GND.n741 GND.n740 3.324
R5207 GND.n3114 GND.n3113 3.324
R5208 GND.n2803 GND.n2802 3.324
R5209 GND.n5838 GND.n5837 3.011
R5210 GND.n5734 GND.n5733 3.011
R5211 GND.n5658 GND.n5657 3.011
R5212 GND.n5554 GND.n5553 3.011
R5213 GND.n1868 GND.n1867 3.011
R5214 GND.n1972 GND.n1971 3.011
R5215 GND.n2048 GND.n2047 3.011
R5216 GND.n2152 GND.n2151 3.011
R5217 GND.n5178 GND.n5177 3.011
R5218 GND.n5282 GND.n5281 3.011
R5219 GND.n5358 GND.n5357 3.011
R5220 GND.n5462 GND.n5461 3.011
R5221 GND.n4428 GND.n4427 3.011
R5222 GND.n4532 GND.n4531 3.011
R5223 GND.n4608 GND.n4607 3.011
R5224 GND.n4717 GND.n4716 3.011
R5225 GND.n4799 GND.n4798 3.011
R5226 GND.n4903 GND.n4902 3.011
R5227 GND.n4979 GND.n4978 3.011
R5228 GND.n5083 GND.n5082 3.011
R5229 GND.n3542 GND.n3541 3.011
R5230 GND.n3433 GND.n3432 3.011
R5231 GND.n3356 GND.n3355 3.011
R5232 GND.n3252 GND.n3251 3.011
R5233 GND.n3749 GND.n3748 3.011
R5234 GND.n3645 GND.n3644 3.011
R5235 GND.n4157 GND.n4156 3.011
R5236 GND.n4261 GND.n4260 3.011
R5237 GND.n3159 GND.n3158 3.011
R5238 GND.n3055 GND.n3054 3.011
R5239 GND.n2752 GND.n2751 3.011
R5240 GND.n2856 GND.n2855 3.011
R5241 GND.n1231 GND.n1230 3.011
R5242 GND.n1127 GND.n1126 3.011
R5243 GND.n690 GND.n689 3.011
R5244 GND.n794 GND.n793 3.011
R5245 GND.n1736 GND.n1735 3.011
R5246 GND.n1632 GND.n1631 3.011
R5247 GND.n1324 GND.n1323 3.011
R5248 GND.n1428 GND.n1427 3.011
R5249 GND.n8004 GND.n8003 3
R5250 GND.n7956 GND.n7955 3
R5251 GND.n7965 GND.n7964 3
R5252 GND.n7992 GND.n7991 3
R5253 GND.n7902 GND.n7901 3
R5254 GND.n7876 GND.n7875 3
R5255 GND.n7930 GND.n7929 3
R5256 GND.n8030 GND.n8029 3
R5257 GND.n7777 GND.n7776 3
R5258 GND.n7729 GND.n7728 3
R5259 GND.n7738 GND.n7737 3
R5260 GND.n7765 GND.n7764 3
R5261 GND.n7675 GND.n7674 3
R5262 GND.n7649 GND.n7648 3
R5263 GND.n7703 GND.n7702 3
R5264 GND.n7803 GND.n7802 3
R5265 GND.n7550 GND.n7549 3
R5266 GND.n7502 GND.n7501 3
R5267 GND.n7511 GND.n7510 3
R5268 GND.n7538 GND.n7537 3
R5269 GND.n7448 GND.n7447 3
R5270 GND.n7422 GND.n7421 3
R5271 GND.n7476 GND.n7475 3
R5272 GND.n7576 GND.n7575 3
R5273 GND.n7323 GND.n7322 3
R5274 GND.n7275 GND.n7274 3
R5275 GND.n7284 GND.n7283 3
R5276 GND.n7311 GND.n7310 3
R5277 GND.n7221 GND.n7220 3
R5278 GND.n7195 GND.n7194 3
R5279 GND.n7249 GND.n7248 3
R5280 GND.n7349 GND.n7348 3
R5281 GND.n7096 GND.n7095 3
R5282 GND.n7048 GND.n7047 3
R5283 GND.n7057 GND.n7056 3
R5284 GND.n7084 GND.n7083 3
R5285 GND.n6994 GND.n6993 3
R5286 GND.n6968 GND.n6967 3
R5287 GND.n7022 GND.n7021 3
R5288 GND.n7122 GND.n7121 3
R5289 GND.n6869 GND.n6868 3
R5290 GND.n6821 GND.n6820 3
R5291 GND.n6830 GND.n6829 3
R5292 GND.n6857 GND.n6856 3
R5293 GND.n6767 GND.n6766 3
R5294 GND.n6741 GND.n6740 3
R5295 GND.n6795 GND.n6794 3
R5296 GND.n6895 GND.n6894 3
R5297 GND.n6537 GND.n6536 3
R5298 GND.n6463 GND.n6397 3
R5299 GND.n6489 GND.n6488 3
R5300 GND.n6498 GND.n6497 3
R5301 GND.n6525 GND.n6524 3
R5302 GND.n6421 GND.n6420 3
R5303 GND.n6446 GND.n6408 3
R5304 GND.n6563 GND.n6562 3
R5305 GND.n593 GND.n592 3
R5306 GND.n6063 GND.n6062 3
R5307 GND.n3891 GND.n3890 3
R5308 GND.n2359 GND.n2358 3
R5309 GND.n4012 GND.n4011 3
R5310 GND.n6308 GND.n6307 3
R5311 GND.n5831 GND.n5826 2.635
R5312 GND.n5751 GND.n5746 2.635
R5313 GND.n5651 GND.n5646 2.635
R5314 GND.n5571 GND.n5566 2.635
R5315 GND.n1885 GND.n1880 2.635
R5316 GND.n1965 GND.n1960 2.635
R5317 GND.n2065 GND.n2060 2.635
R5318 GND.n2145 GND.n2140 2.635
R5319 GND.n5195 GND.n5190 2.635
R5320 GND.n5275 GND.n5270 2.635
R5321 GND.n5375 GND.n5370 2.635
R5322 GND.n5455 GND.n5450 2.635
R5323 GND.n4445 GND.n4440 2.635
R5324 GND.n4525 GND.n4520 2.635
R5325 GND.n4626 GND.n4620 2.635
R5326 GND.n4710 GND.n4704 2.635
R5327 GND.n4816 GND.n4811 2.635
R5328 GND.n4896 GND.n4891 2.635
R5329 GND.n4996 GND.n4991 2.635
R5330 GND.n5076 GND.n5071 2.635
R5331 GND.n3535 GND.n3529 2.635
R5332 GND.n3451 GND.n3445 2.635
R5333 GND.n3349 GND.n3344 2.635
R5334 GND.n3269 GND.n3264 2.635
R5335 GND.n3742 GND.n3737 2.635
R5336 GND.n3662 GND.n3657 2.635
R5337 GND.n4174 GND.n4169 2.635
R5338 GND.n4254 GND.n4249 2.635
R5339 GND.n3152 GND.n3147 2.635
R5340 GND.n3072 GND.n3067 2.635
R5341 GND.n2769 GND.n2764 2.635
R5342 GND.n2849 GND.n2844 2.635
R5343 GND.n1224 GND.n1219 2.635
R5344 GND.n1144 GND.n1139 2.635
R5345 GND.n707 GND.n702 2.635
R5346 GND.n787 GND.n782 2.635
R5347 GND.n1729 GND.n1724 2.635
R5348 GND.n1649 GND.n1644 2.635
R5349 GND.n1341 GND.n1336 2.635
R5350 GND.n1421 GND.n1416 2.635
R5351 GND.n7885 GND.n7884 2.473
R5352 GND.n7984 GND.n7983 2.473
R5353 GND.n7890 GND.n7863 2.473
R5354 GND.n7918 GND.n7917 2.473
R5355 GND.n7934 GND.n7853 2.473
R5356 GND.n8013 GND.n8012 2.473
R5357 GND.n7972 GND.n7971 2.473
R5358 GND.n7946 GND.n7945 2.473
R5359 GND.n7658 GND.n7657 2.473
R5360 GND.n7757 GND.n7756 2.473
R5361 GND.n7663 GND.n7636 2.473
R5362 GND.n7691 GND.n7690 2.473
R5363 GND.n7707 GND.n7626 2.473
R5364 GND.n7786 GND.n7785 2.473
R5365 GND.n7745 GND.n7744 2.473
R5366 GND.n7719 GND.n7718 2.473
R5367 GND.n7431 GND.n7430 2.473
R5368 GND.n7530 GND.n7529 2.473
R5369 GND.n7436 GND.n7409 2.473
R5370 GND.n7464 GND.n7463 2.473
R5371 GND.n7480 GND.n7399 2.473
R5372 GND.n7559 GND.n7558 2.473
R5373 GND.n7518 GND.n7517 2.473
R5374 GND.n7492 GND.n7491 2.473
R5375 GND.n7204 GND.n7203 2.473
R5376 GND.n7303 GND.n7302 2.473
R5377 GND.n7209 GND.n7182 2.473
R5378 GND.n7237 GND.n7236 2.473
R5379 GND.n7253 GND.n7172 2.473
R5380 GND.n7332 GND.n7331 2.473
R5381 GND.n7291 GND.n7290 2.473
R5382 GND.n7265 GND.n7264 2.473
R5383 GND.n6977 GND.n6976 2.473
R5384 GND.n7076 GND.n7075 2.473
R5385 GND.n6982 GND.n6955 2.473
R5386 GND.n7010 GND.n7009 2.473
R5387 GND.n7026 GND.n6945 2.473
R5388 GND.n7105 GND.n7104 2.473
R5389 GND.n7064 GND.n7063 2.473
R5390 GND.n7038 GND.n7037 2.473
R5391 GND.n6750 GND.n6749 2.473
R5392 GND.n6849 GND.n6848 2.473
R5393 GND.n6755 GND.n6728 2.473
R5394 GND.n6783 GND.n6782 2.473
R5395 GND.n6799 GND.n6718 2.473
R5396 GND.n6878 GND.n6877 2.473
R5397 GND.n6837 GND.n6836 2.473
R5398 GND.n6811 GND.n6810 2.473
R5399 GND.n6430 GND.n6429 2.473
R5400 GND.n6517 GND.n6516 2.473
R5401 GND.n6445 GND.n6444 2.473
R5402 GND.n6462 GND.n6461 2.473
R5403 GND.n6467 GND.n6386 2.473
R5404 GND.n6546 GND.n6545 2.473
R5405 GND.n6505 GND.n6504 2.473
R5406 GND.n6479 GND.n6478 2.473
R5407 GND.n5850 GND.n5849 2.258
R5408 GND.n5722 GND.n5721 2.258
R5409 GND.n5670 GND.n5669 2.258
R5410 GND.n5541 GND.n5540 2.258
R5411 GND.n1856 GND.n1855 2.258
R5412 GND.n1984 GND.n1983 2.258
R5413 GND.n2036 GND.n2035 2.258
R5414 GND.n2164 GND.n2163 2.258
R5415 GND.n5166 GND.n5165 2.258
R5416 GND.n5294 GND.n5293 2.258
R5417 GND.n5346 GND.n5345 2.258
R5418 GND.n5474 GND.n5473 2.258
R5419 GND.n4416 GND.n4415 2.258
R5420 GND.n4544 GND.n4543 2.258
R5421 GND.n4596 GND.n4595 2.258
R5422 GND.n4729 GND.n4728 2.258
R5423 GND.n4787 GND.n4786 2.258
R5424 GND.n4915 GND.n4914 2.258
R5425 GND.n4967 GND.n4966 2.258
R5426 GND.n5095 GND.n5094 2.258
R5427 GND.n3554 GND.n3553 2.258
R5428 GND.n3420 GND.n3419 2.258
R5429 GND.n3368 GND.n3367 2.258
R5430 GND.n3239 GND.n3238 2.258
R5431 GND.n3761 GND.n3760 2.258
R5432 GND.n3633 GND.n3632 2.258
R5433 GND.n4145 GND.n4144 2.258
R5434 GND.n4273 GND.n4272 2.258
R5435 GND.n3171 GND.n3170 2.258
R5436 GND.n3043 GND.n3042 2.258
R5437 GND.n2740 GND.n2739 2.258
R5438 GND.n2868 GND.n2867 2.258
R5439 GND.n1243 GND.n1242 2.258
R5440 GND.n1115 GND.n1114 2.258
R5441 GND.n678 GND.n677 2.258
R5442 GND.n806 GND.n805 2.258
R5443 GND.n1748 GND.n1747 2.258
R5444 GND.n1620 GND.n1619 2.258
R5445 GND.n1312 GND.n1311 2.258
R5446 GND.n1440 GND.n1439 2.258
R5447 GND.n4684 GND.n4683 2.163
R5448 GND.n4709 GND.n4708 2.163
R5449 GND.n4734 GND.n4733 2.163
R5450 GND.n4625 GND.n4624 2.163
R5451 GND.n4650 GND.n4649 2.163
R5452 GND.n3475 GND.n3474 2.163
R5453 GND.n3450 GND.n3449 2.163
R5454 GND.n3425 GND.n3424 2.163
R5455 GND.n3559 GND.n3558 2.163
R5456 GND.n3534 GND.n3533 2.163
R5457 GND.n3509 GND.n3508 2.163
R5458 GND.n3244 GND.n3243 2.163
R5459 GND.n5546 GND.n5545 2.163
R5460 GND.n1445 GND.n1444 2.163
R5461 GND.n5819 GND.n5814 1.882
R5462 GND.n5763 GND.n5758 1.882
R5463 GND.n5639 GND.n5634 1.882
R5464 GND.n5583 GND.n5578 1.882
R5465 GND.n1897 GND.n1892 1.882
R5466 GND.n1953 GND.n1948 1.882
R5467 GND.n2077 GND.n2072 1.882
R5468 GND.n2133 GND.n2128 1.882
R5469 GND.n5207 GND.n5202 1.882
R5470 GND.n5263 GND.n5258 1.882
R5471 GND.n5387 GND.n5382 1.882
R5472 GND.n5443 GND.n5438 1.882
R5473 GND.n4457 GND.n4452 1.882
R5474 GND.n4513 GND.n4508 1.882
R5475 GND.n4638 GND.n4633 1.882
R5476 GND.n4697 GND.n4692 1.882
R5477 GND.n4828 GND.n4823 1.882
R5478 GND.n4884 GND.n4879 1.882
R5479 GND.n5008 GND.n5003 1.882
R5480 GND.n5064 GND.n5059 1.882
R5481 GND.n3522 GND.n3517 1.882
R5482 GND.n3463 GND.n3458 1.882
R5483 GND.n3337 GND.n3332 1.882
R5484 GND.n3281 GND.n3276 1.882
R5485 GND.n3730 GND.n3725 1.882
R5486 GND.n3674 GND.n3669 1.882
R5487 GND.n4186 GND.n4181 1.882
R5488 GND.n4242 GND.n4237 1.882
R5489 GND.n3140 GND.n3135 1.882
R5490 GND.n3084 GND.n3079 1.882
R5491 GND.n2781 GND.n2776 1.882
R5492 GND.n2837 GND.n2832 1.882
R5493 GND.n1212 GND.n1207 1.882
R5494 GND.n1156 GND.n1151 1.882
R5495 GND.n719 GND.n714 1.882
R5496 GND.n775 GND.n770 1.882
R5497 GND.n1717 GND.n1712 1.882
R5498 GND.n1661 GND.n1656 1.882
R5499 GND.n1353 GND.n1348 1.882
R5500 GND.n1409 GND.n1404 1.882
R5501 GND.n1021 GND.n1020 1.801
R5502 GND.n2643 GND.n2642 1.801
R5503 GND.n8289 GND.n8216 1.596
R5504 GND.n8468 GND.n8467 1.596
R5505 GND.n8653 GND.n8652 1.596
R5506 GND.n8838 GND.n8837 1.596
R5507 GND.n9023 GND.n9022 1.596
R5508 GND.n9208 GND.n9207 1.596
R5509 GND.n169 GND.n168 1.596
R5510 GND.n5874 GND.n5873 1.505
R5511 GND.n5866 GND.n5865 1.505
R5512 GND.n5710 GND.n5709 1.505
R5513 GND.n5682 GND.n5681 1.505
R5514 GND.n1827 GND.n1826 1.505
R5515 GND.n5532 GND.n1834 1.505
R5516 GND.n1820 GND.n1819 1.505
R5517 GND.n1812 GND.n1811 1.505
R5518 GND.n1996 GND.n1995 1.505
R5519 GND.n2024 GND.n2023 1.505
R5520 GND.n1840 GND.n1839 1.505
R5521 GND.n2178 GND.n1847 1.505
R5522 GND.n1807 GND.n1806 1.505
R5523 GND.n1799 GND.n1798 1.505
R5524 GND.n5306 GND.n5305 1.505
R5525 GND.n5334 GND.n5333 1.505
R5526 GND.n5150 GND.n5149 1.505
R5527 GND.n5488 GND.n5157 1.505
R5528 GND.n1794 GND.n1793 1.505
R5529 GND.n1786 GND.n1785 1.505
R5530 GND.n4556 GND.n4555 1.505
R5531 GND.n4584 GND.n4583 1.505
R5532 GND.n4399 GND.n4398 1.505
R5533 GND.n4744 GND.n4407 1.505
R5534 GND.n1781 GND.n1780 1.505
R5535 GND.n1773 GND.n1772 1.505
R5536 GND.n4927 GND.n4926 1.505
R5537 GND.n4955 GND.n4954 1.505
R5538 GND.n4771 GND.n4770 1.505
R5539 GND.n5109 GND.n4778 1.505
R5540 GND.n3579 GND.n3578 1.505
R5541 GND.n3571 GND.n3570 1.505
R5542 GND.n3408 GND.n3407 1.505
R5543 GND.n3380 GND.n3379 1.505
R5544 GND.n3201 GND.n3200 1.505
R5545 GND.n3230 GND.n3208 1.505
R5546 GND.n3775 GND.n3617 1.505
R5547 GND.n3610 GND.n3609 1.505
R5548 GND.n3621 GND.n3620 1.505
R5549 GND.n4132 GND.n4131 1.505
R5550 GND.n4285 GND.n4284 1.505
R5551 GND.n3183 GND.n3182 1.505
R5552 GND.n3030 GND.n3029 1.505
R5553 GND.n2727 GND.n2726 1.505
R5554 GND.n2880 GND.n2879 1.505
R5555 GND.n3594 GND.n3591 1.505
R5556 GND.n1257 GND.n1099 1.505
R5557 GND.n1092 GND.n1091 1.505
R5558 GND.n1103 GND.n1102 1.505
R5559 GND.n6150 GND.n6149 1.505
R5560 GND.n663 GND.n662 1.505
R5561 GND.n671 GND.n670 1.505
R5562 GND.n3225 GND.n3222 1.505
R5563 GND.n1760 GND.n1759 1.505
R5564 GND.n1607 GND.n1606 1.505
R5565 GND.n1299 GND.n1298 1.505
R5566 GND.n1453 GND.n1452 1.505
R5567 GND.n8289 GND.n8288 1.356
R5568 GND.n8468 GND.n8395 1.356
R5569 GND.n8653 GND.n8580 1.356
R5570 GND.n8838 GND.n8765 1.356
R5571 GND.n9023 GND.n8950 1.356
R5572 GND.n9208 GND.n9135 1.356
R5573 GND.n169 GND.n96 1.356
R5574 GND.n8271 GND.n8270 1.155
R5575 GND.n8378 GND.n8377 1.155
R5576 GND.n8563 GND.n8562 1.155
R5577 GND.n8748 GND.n8747 1.155
R5578 GND.n8933 GND.n8932 1.155
R5579 GND.n9118 GND.n9117 1.155
R5580 GND.n79 GND.n78 1.155
R5581 GND.n8197 GND.n8196 1.155
R5582 GND.n8449 GND.n8448 1.155
R5583 GND.n8634 GND.n8633 1.155
R5584 GND.n8819 GND.n8818 1.155
R5585 GND.n9004 GND.n9003 1.155
R5586 GND.n9189 GND.n9188 1.155
R5587 GND.n150 GND.n149 1.155
R5588 GND.n7938 GND.n7937 1.155
R5589 GND.n7948 GND.n7947 1.155
R5590 GND.n7711 GND.n7710 1.155
R5591 GND.n7721 GND.n7720 1.155
R5592 GND.n7484 GND.n7483 1.155
R5593 GND.n7494 GND.n7493 1.155
R5594 GND.n7257 GND.n7256 1.155
R5595 GND.n7267 GND.n7266 1.155
R5596 GND.n7030 GND.n7029 1.155
R5597 GND.n7040 GND.n7039 1.155
R5598 GND.n6803 GND.n6802 1.155
R5599 GND.n6813 GND.n6812 1.155
R5600 GND.n6471 GND.n6470 1.155
R5601 GND.n6481 GND.n6480 1.155
R5602 GND.n5807 GND.n5802 1.129
R5603 GND.n5775 GND.n5770 1.129
R5604 GND.n5627 GND.n5622 1.129
R5605 GND.n5595 GND.n5590 1.129
R5606 GND.n1909 GND.n1904 1.129
R5607 GND.n1941 GND.n1936 1.129
R5608 GND.n2089 GND.n2084 1.129
R5609 GND.n2121 GND.n2116 1.129
R5610 GND.n5219 GND.n5214 1.129
R5611 GND.n5251 GND.n5246 1.129
R5612 GND.n5399 GND.n5394 1.129
R5613 GND.n5431 GND.n5426 1.129
R5614 GND.n4469 GND.n4464 1.129
R5615 GND.n4501 GND.n4496 1.129
R5616 GND.n4651 GND.n4645 1.129
R5617 GND.n4685 GND.n4679 1.129
R5618 GND.n4840 GND.n4835 1.129
R5619 GND.n4872 GND.n4867 1.129
R5620 GND.n5020 GND.n5015 1.129
R5621 GND.n5052 GND.n5047 1.129
R5622 GND.n3510 GND.n3504 1.129
R5623 GND.n3476 GND.n3470 1.129
R5624 GND.n3325 GND.n3320 1.129
R5625 GND.n3293 GND.n3288 1.129
R5626 GND.n3718 GND.n3713 1.129
R5627 GND.n3686 GND.n3681 1.129
R5628 GND.n4198 GND.n4193 1.129
R5629 GND.n4230 GND.n4225 1.129
R5630 GND.n3128 GND.n3123 1.129
R5631 GND.n3096 GND.n3091 1.129
R5632 GND.n2793 GND.n2788 1.129
R5633 GND.n2825 GND.n2820 1.129
R5634 GND.n1200 GND.n1195 1.129
R5635 GND.n1168 GND.n1163 1.129
R5636 GND.n731 GND.n726 1.129
R5637 GND.n763 GND.n758 1.129
R5638 GND.n1705 GND.n1700 1.129
R5639 GND.n1673 GND.n1668 1.129
R5640 GND.n1365 GND.n1360 1.129
R5641 GND.n1397 GND.n1392 1.129
R5642 GND.n7939 GND.n7938 0.879
R5643 GND.n7949 GND.n7948 0.879
R5644 GND.n7712 GND.n7711 0.879
R5645 GND.n7722 GND.n7721 0.879
R5646 GND.n7485 GND.n7484 0.879
R5647 GND.n7495 GND.n7494 0.879
R5648 GND.n7258 GND.n7257 0.879
R5649 GND.n7268 GND.n7267 0.879
R5650 GND.n7031 GND.n7030 0.879
R5651 GND.n7041 GND.n7040 0.879
R5652 GND.n6804 GND.n6803 0.879
R5653 GND.n6814 GND.n6813 0.879
R5654 GND.n6472 GND.n6471 0.879
R5655 GND.n6482 GND.n6481 0.879
R5656 GND.n8272 GND.n8271 0.857
R5657 GND.n8379 GND.n8378 0.857
R5658 GND.n8564 GND.n8563 0.857
R5659 GND.n8749 GND.n8748 0.857
R5660 GND.n8934 GND.n8933 0.857
R5661 GND.n9119 GND.n9118 0.857
R5662 GND.n80 GND.n79 0.857
R5663 GND.n8198 GND.n8197 0.857
R5664 GND.n8450 GND.n8449 0.857
R5665 GND.n8635 GND.n8634 0.857
R5666 GND.n8820 GND.n8819 0.857
R5667 GND.n9005 GND.n9004 0.857
R5668 GND.n9190 GND.n9189 0.857
R5669 GND.n151 GND.n150 0.857
R5670 GND.n8109 GND.n8108 0.853
R5671 GND.n8142 GND.n8123 0.853
R5672 GND.n8290 GND.n8289 0.853
R5673 GND.n8297 GND.n8296 0.853
R5674 GND.n8121 GND.n8120 0.853
R5675 GND.n8101 GND.n8100 0.853
R5676 GND.n8128 GND.n8127 0.853
R5677 GND.n8141 GND.n8140 0.853
R5678 GND.n445 GND.n444 0.853
R5679 GND.n8489 GND.n8488 0.853
R5680 GND.n8469 GND.n8468 0.853
R5681 GND.n419 GND.n418 0.853
R5682 GND.n411 GND.n410 0.853
R5683 GND.n438 GND.n437 0.853
R5684 GND.n450 GND.n448 0.853
R5685 GND.n8480 GND.n8479 0.853
R5686 GND.n8490 GND.n8473 0.853
R5687 GND.n421 GND.n414 0.853
R5688 GND.n435 GND.n434 0.853
R5689 GND.n396 GND.n395 0.853
R5690 GND.n8674 GND.n8673 0.853
R5691 GND.n8654 GND.n8653 0.853
R5692 GND.n370 GND.n369 0.853
R5693 GND.n362 GND.n361 0.853
R5694 GND.n389 GND.n388 0.853
R5695 GND.n401 GND.n399 0.853
R5696 GND.n8665 GND.n8664 0.853
R5697 GND.n8675 GND.n8658 0.853
R5698 GND.n372 GND.n365 0.853
R5699 GND.n386 GND.n385 0.853
R5700 GND.n347 GND.n346 0.853
R5701 GND.n8859 GND.n8858 0.853
R5702 GND.n8839 GND.n8838 0.853
R5703 GND.n321 GND.n320 0.853
R5704 GND.n313 GND.n312 0.853
R5705 GND.n340 GND.n339 0.853
R5706 GND.n352 GND.n350 0.853
R5707 GND.n8850 GND.n8849 0.853
R5708 GND.n8860 GND.n8843 0.853
R5709 GND.n323 GND.n316 0.853
R5710 GND.n337 GND.n336 0.853
R5711 GND.n298 GND.n297 0.853
R5712 GND.n9044 GND.n9043 0.853
R5713 GND.n9024 GND.n9023 0.853
R5714 GND.n272 GND.n271 0.853
R5715 GND.n264 GND.n263 0.853
R5716 GND.n291 GND.n290 0.853
R5717 GND.n303 GND.n301 0.853
R5718 GND.n9035 GND.n9034 0.853
R5719 GND.n9045 GND.n9028 0.853
R5720 GND.n274 GND.n267 0.853
R5721 GND.n288 GND.n287 0.853
R5722 GND.n249 GND.n248 0.853
R5723 GND.n9229 GND.n9228 0.853
R5724 GND.n9209 GND.n9208 0.853
R5725 GND.n223 GND.n222 0.853
R5726 GND.n215 GND.n214 0.853
R5727 GND.n242 GND.n241 0.853
R5728 GND.n254 GND.n252 0.853
R5729 GND.n9220 GND.n9219 0.853
R5730 GND.n9230 GND.n9213 0.853
R5731 GND.n225 GND.n218 0.853
R5732 GND.n239 GND.n238 0.853
R5733 GND.n9259 GND.n9258 0.853
R5734 GND.n8302 GND.n8301 0.853
R5735 GND.n8112 GND.n8111 0.853
R5736 GND.n8098 GND.n8097 0.853
R5737 GND.n8131 GND.n8130 0.853
R5738 GND.n654 GND.n653 0.77
R5739 GND.n660 GND.n659 0.77
R5740 GND.n496 GND.n495 0.77
R5741 GND.n502 GND.n501 0.77
R5742 GND.n1280 GND.n1279 0.77
R5743 GND.n1270 GND.n1269 0.77
R5744 GND.n6127 GND.n6126 0.77
R5745 GND.n6134 GND.n6133 0.77
R5746 GND.n3955 GND.n3954 0.77
R5747 GND.n3962 GND.n3961 0.77
R5748 GND.n2420 GND.n2419 0.77
R5749 GND.n4303 GND.n4302 0.77
R5750 GND.n2262 GND.n2261 0.77
R5751 GND.n2268 GND.n2267 0.77
R5752 GND.n3782 GND.n3781 0.752
R5753 GND.n2439 GND.n2438 0.752
R5754 GND.n6325 GND.n6322 0.739
R5755 GND.n1457 GND.n1456 0.644
R5756 GND.n5338 GND.n5337 0.644
R5757 GND.n2028 GND.n2027 0.644
R5758 GND.n4588 GND.n4587 0.644
R5759 GND.n4405 GND.n4404 0.644
R5760 GND.n4959 GND.n4958 0.644
R5761 GND.n1778 GND.n1777 0.644
R5762 GND.n1791 GND.n1790 0.644
R5763 GND.n1804 GND.n1803 0.644
R5764 GND.n1817 GND.n1816 0.644
R5765 GND.n3576 GND.n3575 0.644
R5766 GND.n3412 GND.n3411 0.644
R5767 GND.n3384 GND.n3383 0.644
R5768 GND.n3206 GND.n3205 0.644
R5769 GND.n5871 GND.n5870 0.644
R5770 GND.n5686 GND.n5685 0.644
R5771 GND.n1832 GND.n1831 0.644
R5772 GND.n3615 GND.n3614 0.644
R5773 GND.n4137 GND.n4136 0.644
R5774 GND.n3187 GND.n3186 0.644
R5775 GND.n2732 GND.n2731 0.644
R5776 GND.n1097 GND.n1096 0.644
R5777 GND.n6154 GND.n6153 0.644
R5778 GND.n1764 GND.n1763 0.644
R5779 GND.n1304 GND.n1303 0.644
R5780 GND.n4307 GND.n2257 0.582
R5781 GND.n5350 GND.n5349 0.551
R5782 GND.n2040 GND.n2039 0.551
R5783 GND.n4971 GND.n4970 0.551
R5784 GND.n4791 GND.n4790 0.551
R5785 GND.n4420 GND.n4419 0.551
R5786 GND.n5170 GND.n5169 0.551
R5787 GND.n1860 GND.n1859 0.551
R5788 GND.n3372 GND.n3371 0.551
R5789 GND.n5854 GND.n5853 0.551
R5790 GND.n5674 GND.n5673 0.551
R5791 GND.n3765 GND.n3764 0.551
R5792 GND.n4149 GND.n4148 0.551
R5793 GND.n2744 GND.n2743 0.551
R5794 GND.n3175 GND.n3174 0.551
R5795 GND.n1247 GND.n1246 0.551
R5796 GND.n682 GND.n681 0.551
R5797 GND.n1752 GND.n1751 0.551
R5798 GND.n1316 GND.n1315 0.551
R5799 GND.n6220 GND.n6219 0.536
R5800 GND.n597 GND.n596 0.536
R5801 GND.n609 GND.n608 0.536
R5802 GND.n6079 GND.n6078 0.536
R5803 GND.n987 GND.n986 0.536
R5804 GND.n999 GND.n998 0.536
R5805 GND.n3907 GND.n3906 0.536
R5806 GND.n2609 GND.n2608 0.536
R5807 GND.n2621 GND.n2620 0.536
R5808 GND.n4067 GND.n4066 0.536
R5809 GND.n2363 GND.n2362 0.536
R5810 GND.n2375 GND.n2374 0.536
R5811 GND.n2956 GND.n2955 0.536
R5812 GND.n1535 GND.n1534 0.536
R5813 GND.n890 GND.n889 0.536
R5814 GND.n902 GND.n901 0.536
R5815 GND.n6067 GND.n6066 0.536
R5816 GND.n2512 GND.n2511 0.536
R5817 GND.n2524 GND.n2523 0.536
R5818 GND.n3895 GND.n3894 0.536
R5819 GND.n2968 GND.n2967 0.536
R5820 GND.n4079 GND.n4078 0.536
R5821 GND.n1547 GND.n1546 0.536
R5822 GND.n6208 GND.n6207 0.536
R5823 GND.n7969 GND.n7968 0.506
R5824 GND.n7962 GND.n7961 0.506
R5825 GND.n7742 GND.n7741 0.506
R5826 GND.n7735 GND.n7734 0.506
R5827 GND.n7515 GND.n7514 0.506
R5828 GND.n7508 GND.n7507 0.506
R5829 GND.n7288 GND.n7287 0.506
R5830 GND.n7281 GND.n7280 0.506
R5831 GND.n7061 GND.n7060 0.506
R5832 GND.n7054 GND.n7053 0.506
R5833 GND.n6834 GND.n6833 0.506
R5834 GND.n6827 GND.n6826 0.506
R5835 GND.n6502 GND.n6501 0.506
R5836 GND.n6495 GND.n6494 0.506
R5837 GND.n6232 GND.n6231 0.506
R5838 GND.n565 GND.n563 0.506
R5839 GND.n616 GND.n615 0.506
R5840 GND.n6086 GND.n6085 0.506
R5841 GND.n980 GND.n979 0.506
R5842 GND.n1031 GND.n1030 0.506
R5843 GND.n909 GND.n908 0.506
R5844 GND.n880 GND.n878 0.506
R5845 GND.n3914 GND.n3913 0.506
R5846 GND.n2602 GND.n2601 0.506
R5847 GND.n2653 GND.n2652 0.506
R5848 GND.n2531 GND.n2530 0.506
R5849 GND.n2502 GND.n2500 0.506
R5850 GND.n3981 GND.n3980 0.506
R5851 GND.n2331 GND.n2329 0.506
R5852 GND.n2382 GND.n2381 0.506
R5853 GND.n2718 GND.n2717 0.506
R5854 GND.n1526 GND.n1525 0.506
R5855 GND.n8195 GND.n8193 0.506
R5856 GND.n8446 GND.n8444 0.506
R5857 GND.n8631 GND.n8629 0.506
R5858 GND.n8816 GND.n8814 0.506
R5859 GND.n9001 GND.n8999 0.506
R5860 GND.n9186 GND.n9184 0.506
R5861 GND.n147 GND.n145 0.506
R5862 GND.n6034 GND.n6032 0.506
R5863 GND.n3862 GND.n3860 0.506
R5864 GND.n2975 GND.n2974 0.506
R5865 GND.n4086 GND.n4085 0.506
R5866 GND.n1554 GND.n1553 0.506
R5867 GND.n6201 GND.n6200 0.506
R5868 GND.n8268 GND.n8266 0.506
R5869 GND.n8375 GND.n8373 0.506
R5870 GND.n8560 GND.n8558 0.506
R5871 GND.n8745 GND.n8743 0.506
R5872 GND.n8930 GND.n8928 0.506
R5873 GND.n9115 GND.n9113 0.506
R5874 GND.n76 GND.n74 0.506
R5875 GND.n8008 GND.n8007 0.476
R5876 GND.n8001 GND.n8000 0.476
R5877 GND.n7781 GND.n7780 0.476
R5878 GND.n7774 GND.n7773 0.476
R5879 GND.n7554 GND.n7553 0.476
R5880 GND.n7547 GND.n7546 0.476
R5881 GND.n7327 GND.n7326 0.476
R5882 GND.n7320 GND.n7319 0.476
R5883 GND.n7100 GND.n7099 0.476
R5884 GND.n7093 GND.n7092 0.476
R5885 GND.n6873 GND.n6872 0.476
R5886 GND.n6866 GND.n6865 0.476
R5887 GND.n6541 GND.n6540 0.476
R5888 GND.n6534 GND.n6533 0.476
R5889 GND.n6244 GND.n6243 0.476
R5890 GND.n551 GND.n550 0.476
R5891 GND.n623 GND.n622 0.476
R5892 GND.n6093 GND.n6092 0.476
R5893 GND.n973 GND.n972 0.476
R5894 GND.n1043 GND.n1042 0.476
R5895 GND.n3921 GND.n3920 0.476
R5896 GND.n2595 GND.n2594 0.476
R5897 GND.n2665 GND.n2664 0.476
R5898 GND.n4049 GND.n4048 0.476
R5899 GND.n2317 GND.n2316 0.476
R5900 GND.n2389 GND.n2388 0.476
R5901 GND.n2938 GND.n2937 0.476
R5902 GND.n1512 GND.n1511 0.476
R5903 GND.n866 GND.n865 0.475
R5904 GND.n916 GND.n915 0.475
R5905 GND.n6020 GND.n6019 0.475
R5906 GND.n2488 GND.n2487 0.475
R5907 GND.n2538 GND.n2537 0.475
R5908 GND.n3848 GND.n3847 0.475
R5909 GND.n2982 GND.n2981 0.475
R5910 GND.n4093 GND.n4092 0.475
R5911 GND.n1561 GND.n1560 0.475
R5912 GND.n6194 GND.n6193 0.475
R5913 GND.n8262 GND.n8261 0.475
R5914 GND.n8190 GND.n8189 0.475
R5915 GND.n8369 GND.n8368 0.475
R5916 GND.n8441 GND.n8440 0.475
R5917 GND.n8554 GND.n8553 0.475
R5918 GND.n8626 GND.n8625 0.475
R5919 GND.n8739 GND.n8738 0.475
R5920 GND.n8811 GND.n8810 0.475
R5921 GND.n8924 GND.n8923 0.475
R5922 GND.n8996 GND.n8995 0.475
R5923 GND.n9109 GND.n9108 0.475
R5924 GND.n9181 GND.n9180 0.475
R5925 GND.n70 GND.n69 0.475
R5926 GND.n142 GND.n141 0.475
R5927 GND.n5362 GND.n5361 0.455
R5928 GND.n2052 GND.n2051 0.455
R5929 GND.n4612 GND.n4611 0.455
R5930 GND.n4721 GND.n4720 0.455
R5931 GND.n4983 GND.n4982 0.455
R5932 GND.n4803 GND.n4802 0.455
R5933 GND.n4432 GND.n4431 0.455
R5934 GND.n5182 GND.n5181 0.455
R5935 GND.n1872 GND.n1871 0.455
R5936 GND.n3546 GND.n3545 0.455
R5937 GND.n3437 GND.n3436 0.455
R5938 GND.n3360 GND.n3359 0.455
R5939 GND.n5842 GND.n5841 0.455
R5940 GND.n5662 GND.n5661 0.455
R5941 GND.n3753 GND.n3752 0.455
R5942 GND.n4161 GND.n4160 0.455
R5943 GND.n2756 GND.n2755 0.455
R5944 GND.n3163 GND.n3162 0.455
R5945 GND.n1235 GND.n1234 0.455
R5946 GND.n694 GND.n693 0.455
R5947 GND.n1740 GND.n1739 0.455
R5948 GND.n1328 GND.n1327 0.455
R5949 GND.n6339 GND.n6338 0.453
R5950 GND.n7847 GND.n7846 0.445
R5951 GND.n8026 GND.n8025 0.445
R5952 GND.n7620 GND.n7619 0.445
R5953 GND.n7799 GND.n7798 0.445
R5954 GND.n7393 GND.n7392 0.445
R5955 GND.n7572 GND.n7571 0.445
R5956 GND.n7166 GND.n7165 0.445
R5957 GND.n7345 GND.n7344 0.445
R5958 GND.n6939 GND.n6938 0.445
R5959 GND.n7118 GND.n7117 0.445
R5960 GND.n6712 GND.n6711 0.445
R5961 GND.n6891 GND.n6890 0.445
R5962 GND.n6380 GND.n6379 0.445
R5963 GND.n6559 GND.n6558 0.445
R5964 GND.n6255 GND.n6254 0.445
R5965 GND.n540 GND.n539 0.445
R5966 GND.n630 GND.n629 0.445
R5967 GND.n6100 GND.n6099 0.445
R5968 GND.n966 GND.n965 0.445
R5969 GND.n1054 GND.n1053 0.445
R5970 GND.n923 GND.n922 0.445
R5971 GND.n3928 GND.n3927 0.445
R5972 GND.n2588 GND.n2587 0.445
R5973 GND.n2676 GND.n2675 0.445
R5974 GND.n2545 GND.n2544 0.445
R5975 GND.n4039 GND.n4038 0.445
R5976 GND.n2306 GND.n2305 0.445
R5977 GND.n2396 GND.n2395 0.445
R5978 GND.n2928 GND.n2927 0.445
R5979 GND.n1501 GND.n1500 0.445
R5980 GND.n855 GND.n854 0.445
R5981 GND.n6009 GND.n6008 0.445
R5982 GND.n2477 GND.n2476 0.445
R5983 GND.n3837 GND.n3836 0.445
R5984 GND.n2989 GND.n2988 0.445
R5985 GND.n4100 GND.n4099 0.445
R5986 GND.n1568 GND.n1567 0.445
R5987 GND.n6187 GND.n6186 0.445
R5988 GND.n8250 GND.n8249 0.445
R5989 GND.n8178 GND.n8177 0.445
R5990 GND.n8357 GND.n8356 0.445
R5991 GND.n8429 GND.n8428 0.445
R5992 GND.n8542 GND.n8541 0.445
R5993 GND.n8614 GND.n8613 0.445
R5994 GND.n8727 GND.n8726 0.445
R5995 GND.n8799 GND.n8798 0.445
R5996 GND.n8912 GND.n8911 0.445
R5997 GND.n8984 GND.n8983 0.445
R5998 GND.n9097 GND.n9096 0.445
R5999 GND.n9169 GND.n9168 0.445
R6000 GND.n58 GND.n57 0.445
R6001 GND.n130 GND.n129 0.445
R6002 GND.n8032 GND.n8031 0.426
R6003 GND.n7805 GND.n7804 0.426
R6004 GND.n7578 GND.n7577 0.426
R6005 GND.n7351 GND.n7350 0.426
R6006 GND.n7124 GND.n7123 0.426
R6007 GND.n6897 GND.n6896 0.426
R6008 GND.n6580 GND.n6564 0.426
R6009 GND.n7913 GND.n7912 0.414
R6010 GND.n7927 GND.n7926 0.414
R6011 GND.n7686 GND.n7685 0.414
R6012 GND.n7700 GND.n7699 0.414
R6013 GND.n7459 GND.n7458 0.414
R6014 GND.n7473 GND.n7472 0.414
R6015 GND.n7232 GND.n7231 0.414
R6016 GND.n7246 GND.n7245 0.414
R6017 GND.n7005 GND.n7004 0.414
R6018 GND.n7019 GND.n7018 0.414
R6019 GND.n6778 GND.n6777 0.414
R6020 GND.n6792 GND.n6791 0.414
R6021 GND.n6457 GND.n6456 0.414
R6022 GND.n6395 GND.n6394 0.414
R6023 GND.n6266 GND.n6265 0.414
R6024 GND.n529 GND.n528 0.414
R6025 GND.n637 GND.n636 0.414
R6026 GND.n6107 GND.n6106 0.414
R6027 GND.n959 GND.n958 0.414
R6028 GND.n1065 GND.n1064 0.414
R6029 GND.n3935 GND.n3934 0.414
R6030 GND.n2581 GND.n2580 0.414
R6031 GND.n2687 GND.n2686 0.414
R6032 GND.n4029 GND.n4028 0.414
R6033 GND.n2295 GND.n2294 0.414
R6034 GND.n2403 GND.n2402 0.414
R6035 GND.n2918 GND.n2917 0.414
R6036 GND.n1491 GND.n1490 0.414
R6037 GND.n844 GND.n843 0.413
R6038 GND.n930 GND.n929 0.413
R6039 GND.n5998 GND.n5997 0.413
R6040 GND.n2466 GND.n2465 0.413
R6041 GND.n2552 GND.n2551 0.413
R6042 GND.n3826 GND.n3825 0.413
R6043 GND.n2996 GND.n2995 0.413
R6044 GND.n4107 GND.n4106 0.413
R6045 GND.n1575 GND.n1574 0.413
R6046 GND.n6180 GND.n6179 0.413
R6047 GND.n8239 GND.n8238 0.413
R6048 GND.n8167 GND.n8166 0.413
R6049 GND.n8346 GND.n8345 0.413
R6050 GND.n8418 GND.n8417 0.413
R6051 GND.n8531 GND.n8530 0.413
R6052 GND.n8603 GND.n8602 0.413
R6053 GND.n8716 GND.n8715 0.413
R6054 GND.n8788 GND.n8787 0.413
R6055 GND.n8901 GND.n8900 0.413
R6056 GND.n8973 GND.n8972 0.413
R6057 GND.n9086 GND.n9085 0.413
R6058 GND.n9158 GND.n9157 0.413
R6059 GND.n47 GND.n46 0.413
R6060 GND.n119 GND.n118 0.413
R6061 GND.n4397 GND.n4396 0.412
R6062 GND.n2211 GND.n2210 0.412
R6063 GND.n2190 GND.n2189 0.412
R6064 GND.n5499 GND.n4388 0.412
R6065 GND.n4330 GND.n4329 0.412
R6066 GND.n4315 GND.n4314 0.412
R6067 GND.n4309 GND.n4308 0.412
R6068 GND.n2238 GND.n2237 0.412
R6069 GND.n7860 GND.n7859 0.382
R6070 GND.n7899 GND.n7898 0.382
R6071 GND.n7633 GND.n7632 0.382
R6072 GND.n7672 GND.n7671 0.382
R6073 GND.n7406 GND.n7405 0.382
R6074 GND.n7445 GND.n7444 0.382
R6075 GND.n7179 GND.n7178 0.382
R6076 GND.n7218 GND.n7217 0.382
R6077 GND.n6952 GND.n6951 0.382
R6078 GND.n6991 GND.n6990 0.382
R6079 GND.n6725 GND.n6724 0.382
R6080 GND.n6764 GND.n6763 0.382
R6081 GND.n6441 GND.n6440 0.382
R6082 GND.n6406 GND.n6405 0.382
R6083 GND.n6277 GND.n6276 0.382
R6084 GND.n518 GND.n517 0.382
R6085 GND.n644 GND.n643 0.382
R6086 GND.n6114 GND.n6113 0.382
R6087 GND.n952 GND.n951 0.382
R6088 GND.n1076 GND.n1075 0.382
R6089 GND.n937 GND.n936 0.382
R6090 GND.n3942 GND.n3941 0.382
R6091 GND.n2574 GND.n2573 0.382
R6092 GND.n2698 GND.n2697 0.382
R6093 GND.n2559 GND.n2558 0.382
R6094 GND.n4019 GND.n4018 0.382
R6095 GND.n2284 GND.n2283 0.382
R6096 GND.n2410 GND.n2409 0.382
R6097 GND.n2908 GND.n2907 0.382
R6098 GND.n1481 GND.n1480 0.382
R6099 GND.n833 GND.n832 0.382
R6100 GND.n5987 GND.n5986 0.382
R6101 GND.n2455 GND.n2454 0.382
R6102 GND.n3815 GND.n3814 0.382
R6103 GND.n3003 GND.n3002 0.382
R6104 GND.n4114 GND.n4113 0.382
R6105 GND.n1582 GND.n1581 0.382
R6106 GND.n6173 GND.n6172 0.382
R6107 GND.n8228 GND.n8227 0.382
R6108 GND.n8156 GND.n8155 0.382
R6109 GND.n8335 GND.n8334 0.382
R6110 GND.n8407 GND.n8406 0.382
R6111 GND.n8520 GND.n8519 0.382
R6112 GND.n8592 GND.n8591 0.382
R6113 GND.n8705 GND.n8704 0.382
R6114 GND.n8777 GND.n8776 0.382
R6115 GND.n8890 GND.n8889 0.382
R6116 GND.n8962 GND.n8961 0.382
R6117 GND.n9075 GND.n9074 0.382
R6118 GND.n9147 GND.n9146 0.382
R6119 GND.n36 GND.n35 0.382
R6120 GND.n108 GND.n107 0.382
R6121 GND.n5795 GND.n5790 0.376
R6122 GND.n5787 GND.n5782 0.376
R6123 GND.n5615 GND.n5610 0.376
R6124 GND.n5607 GND.n5602 0.376
R6125 GND.n1921 GND.n1916 0.376
R6126 GND.n1929 GND.n1924 0.376
R6127 GND.n2101 GND.n2096 0.376
R6128 GND.n2109 GND.n2104 0.376
R6129 GND.n5231 GND.n5226 0.376
R6130 GND.n5239 GND.n5234 0.376
R6131 GND.n5411 GND.n5406 0.376
R6132 GND.n5419 GND.n5414 0.376
R6133 GND.n4481 GND.n4476 0.376
R6134 GND.n4489 GND.n4484 0.376
R6135 GND.n4663 GND.n4658 0.376
R6136 GND.n4672 GND.n4666 0.376
R6137 GND.n4852 GND.n4847 0.376
R6138 GND.n4860 GND.n4855 0.376
R6139 GND.n5032 GND.n5027 0.376
R6140 GND.n5040 GND.n5035 0.376
R6141 GND.n3497 GND.n3492 0.376
R6142 GND.n3489 GND.n3483 0.376
R6143 GND.n3313 GND.n3308 0.376
R6144 GND.n3305 GND.n3300 0.376
R6145 GND.n3706 GND.n3701 0.376
R6146 GND.n3698 GND.n3693 0.376
R6147 GND.n4210 GND.n4205 0.376
R6148 GND.n4218 GND.n4213 0.376
R6149 GND.n3116 GND.n3111 0.376
R6150 GND.n3108 GND.n3103 0.376
R6151 GND.n2805 GND.n2800 0.376
R6152 GND.n2813 GND.n2808 0.376
R6153 GND.n1188 GND.n1183 0.376
R6154 GND.n1180 GND.n1175 0.376
R6155 GND.n743 GND.n738 0.376
R6156 GND.n751 GND.n746 0.376
R6157 GND.n1693 GND.n1688 0.376
R6158 GND.n1685 GND.n1680 0.376
R6159 GND.n1377 GND.n1372 0.376
R6160 GND.n1385 GND.n1380 0.376
R6161 GND.n5374 GND.n5373 0.358
R6162 GND.n2064 GND.n2063 0.358
R6163 GND.n4995 GND.n4994 0.358
R6164 GND.n4815 GND.n4814 0.358
R6165 GND.n4444 GND.n4443 0.358
R6166 GND.n5194 GND.n5193 0.358
R6167 GND.n1884 GND.n1883 0.358
R6168 GND.n3348 GND.n3347 0.358
R6169 GND.n5830 GND.n5829 0.358
R6170 GND.n5650 GND.n5649 0.358
R6171 GND.n3741 GND.n3740 0.358
R6172 GND.n4173 GND.n4172 0.358
R6173 GND.n2768 GND.n2767 0.358
R6174 GND.n3151 GND.n3150 0.358
R6175 GND.n1223 GND.n1222 0.358
R6176 GND.n706 GND.n705 0.358
R6177 GND.n1728 GND.n1727 0.358
R6178 GND.n1340 GND.n1339 0.358
R6179 GND.n8069 GND.n6586 0.285
R6180 GND.n8303 GND.n8302 0.285
R6181 GND.n5386 GND.n5385 0.259
R6182 GND.n2076 GND.n2075 0.259
R6183 GND.n4637 GND.n4636 0.259
R6184 GND.n4696 GND.n4695 0.259
R6185 GND.n5007 GND.n5006 0.259
R6186 GND.n4827 GND.n4826 0.259
R6187 GND.n4456 GND.n4455 0.259
R6188 GND.n5206 GND.n5205 0.259
R6189 GND.n1896 GND.n1895 0.259
R6190 GND.n3521 GND.n3520 0.259
R6191 GND.n3462 GND.n3461 0.259
R6192 GND.n3336 GND.n3335 0.259
R6193 GND.n5818 GND.n5817 0.259
R6194 GND.n5638 GND.n5637 0.259
R6195 GND.n3729 GND.n3728 0.259
R6196 GND.n4185 GND.n4184 0.259
R6197 GND.n2780 GND.n2779 0.259
R6198 GND.n3139 GND.n3138 0.259
R6199 GND.n1211 GND.n1210 0.259
R6200 GND.n718 GND.n717 0.259
R6201 GND.n1716 GND.n1715 0.259
R6202 GND.n1352 GND.n1351 0.259
R6203 GND.n1601 GND.n1088 0.208
R6204 GND.n3024 GND.n2710 0.208
R6205 GND.n3015 GND.n3012 0.208
R6206 GND.n1592 GND.n1591 0.208
R6207 GND.n9251 GND.n9248 0.19
R6208 GND.n9251 GND.n9242 0.19
R6209 GND.n9251 GND.n9238 0.19
R6210 GND.n9232 GND.n9231 0.19
R6211 GND.n9058 GND.n255 0.19
R6212 GND.n9234 GND.n228 0.19
R6213 GND.n9047 GND.n9046 0.19
R6214 GND.n8873 GND.n304 0.19
R6215 GND.n9049 GND.n277 0.19
R6216 GND.n8862 GND.n8861 0.19
R6217 GND.n8688 GND.n353 0.19
R6218 GND.n8864 GND.n326 0.19
R6219 GND.n8677 GND.n8676 0.19
R6220 GND.n8503 GND.n402 0.19
R6221 GND.n8679 GND.n375 0.19
R6222 GND.n8492 GND.n8491 0.19
R6223 GND.n8318 GND.n451 0.19
R6224 GND.n8494 GND.n424 0.19
R6225 GND.n6922 GND.n6921 0.19
R6226 GND.n6902 GND.n6696 0.19
R6227 GND.n7149 GND.n7148 0.19
R6228 GND.n7129 GND.n6679 0.19
R6229 GND.n7376 GND.n7375 0.19
R6230 GND.n7356 GND.n6662 0.19
R6231 GND.n7603 GND.n7602 0.19
R6232 GND.n7583 GND.n6645 0.19
R6233 GND.n7830 GND.n7829 0.19
R6234 GND.n7810 GND.n6628 0.19
R6235 GND.n8057 GND.n8056 0.19
R6236 GND.n8037 GND.n6611 0.19
R6237 GND.n6899 GND.n6898 0.19
R6238 GND.n7126 GND.n7125 0.19
R6239 GND.n7353 GND.n7352 0.19
R6240 GND.n7580 GND.n7579 0.19
R6241 GND.n7807 GND.n7806 0.19
R6242 GND.n8034 GND.n8033 0.19
R6243 GND.n6142 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/GATE 0.181
R6244 GND.n3970 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/GATE 0.181
R6245 GND.n4126 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/GATE 0.181
R6246 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/GATE GND.n6163 0.181
R6247 GND.n1598 GND.n1595 0.172
R6248 GND.n6148 GND.n6145 0.172
R6249 GND.n3021 GND.n3018 0.172
R6250 GND.n3976 GND.n3973 0.172
R6251 GND.n2012 GND.n2009 0.172
R6252 GND.n2015 GND.n2012 0.172
R6253 GND.n2018 GND.n2015 0.172
R6254 GND.n5322 GND.n5319 0.172
R6255 GND.n5325 GND.n5322 0.172
R6256 GND.n5328 GND.n5325 0.172
R6257 GND.n4572 GND.n4569 0.172
R6258 GND.n4575 GND.n4572 0.172
R6259 GND.n4578 GND.n4575 0.172
R6260 GND.n5143 GND.n5140 0.172
R6261 GND.n5140 GND.n5137 0.172
R6262 GND.n5137 GND.n5134 0.172
R6263 GND.n5130 GND.n5125 0.172
R6264 GND.n5125 GND.n5122 0.172
R6265 GND.n5122 GND.n5119 0.172
R6266 GND.n5119 GND.n5116 0.172
R6267 GND.n4769 GND.n4764 0.172
R6268 GND.n4764 GND.n4761 0.172
R6269 GND.n4761 GND.n4758 0.172
R6270 GND.n4758 GND.n4755 0.172
R6271 GND.n4755 GND.n4752 0.172
R6272 GND.n4943 GND.n4940 0.172
R6273 GND.n4946 GND.n4943 0.172
R6274 GND.n4949 GND.n4946 0.172
R6275 GND.n3402 GND.n3399 0.172
R6276 GND.n3399 GND.n3396 0.172
R6277 GND.n3396 GND.n3393 0.172
R6278 GND.n3608 GND.n3605 0.172
R6279 GND.n3605 GND.n3602 0.172
R6280 GND.n3602 GND.n3599 0.172
R6281 GND.n3595 GND.n3590 0.172
R6282 GND.n3590 GND.n3587 0.172
R6283 GND.n3587 GND.n3584 0.172
R6284 GND.n3584 GND.n1825 0.172
R6285 GND.n5885 GND.n5882 0.172
R6286 GND.n5888 GND.n5885 0.172
R6287 GND.n5891 GND.n5888 0.172
R6288 GND.n5894 GND.n5891 0.172
R6289 GND.n5903 GND.n5900 0.172
R6290 GND.n5906 GND.n5903 0.172
R6291 GND.n5909 GND.n5906 0.172
R6292 GND.n5912 GND.n5909 0.172
R6293 GND.n5921 GND.n5918 0.172
R6294 GND.n5924 GND.n5921 0.172
R6295 GND.n5927 GND.n5924 0.172
R6296 GND.n5930 GND.n5927 0.172
R6297 GND.n5939 GND.n5936 0.172
R6298 GND.n5942 GND.n5939 0.172
R6299 GND.n5945 GND.n5942 0.172
R6300 GND.n5948 GND.n5945 0.172
R6301 GND.n5957 GND.n5954 0.172
R6302 GND.n5960 GND.n5957 0.172
R6303 GND.n5963 GND.n5960 0.172
R6304 GND.n5966 GND.n5963 0.172
R6305 GND.n5704 GND.n5701 0.172
R6306 GND.n5701 GND.n5698 0.172
R6307 GND.n5698 GND.n5695 0.172
R6308 GND.n2434 GND.n2431 0.172
R6309 GND.n2431 GND.n2428 0.172
R6310 GND.n3226 GND.n3221 0.172
R6311 GND.n3221 GND.n3218 0.172
R6312 GND.n3218 GND.n3215 0.172
R6313 GND.n3215 GND.n1838 0.172
R6314 GND.n5528 GND.n5523 0.172
R6315 GND.n5523 GND.n5520 0.172
R6316 GND.n5520 GND.n5517 0.172
R6317 GND.n5517 GND.n5514 0.172
R6318 GND.n4752 GND.n491 0.172
R6319 GND.n605 GND.n602 0.168
R6320 GND.n995 GND.n992 0.168
R6321 GND.n898 GND.n895 0.168
R6322 GND.n6075 GND.n6072 0.168
R6323 GND.n2617 GND.n2614 0.168
R6324 GND.n2520 GND.n2517 0.168
R6325 GND.n3903 GND.n3900 0.168
R6326 GND.n2371 GND.n2368 0.168
R6327 GND.n2964 GND.n2962 0.168
R6328 GND.n4075 GND.n4073 0.168
R6329 GND.n1543 GND.n1541 0.168
R6330 GND.n6216 GND.n6213 0.168
R6331 GND.n5895 GND.n1822 0.165
R6332 GND.n5511 GND.n2181 0.165
R6333 GND.n5913 GND.n1809 0.165
R6334 GND.n5492 GND.n5491 0.165
R6335 GND.n5931 GND.n1796 0.165
R6336 GND.n5131 GND.n4747 0.165
R6337 GND.n5949 GND.n1783 0.165
R6338 GND.n5113 GND.n5112 0.165
R6339 GND.n3596 GND.n3581 0.165
R6340 GND.n3228 GND.n3227 0.165
R6341 GND.n5877 GND.n5876 0.165
R6342 GND.n5530 GND.n5529 0.165
R6343 GND.n2020 GND.n2018 0.163
R6344 GND.n5330 GND.n5328 0.163
R6345 GND.n4580 GND.n4578 0.163
R6346 GND.n4951 GND.n4949 0.163
R6347 GND.n3393 GND.n3390 0.163
R6348 GND.n3599 GND.n3596 0.163
R6349 GND.n5695 GND.n5692 0.163
R6350 GND.n3227 GND.n3212 0.163
R6351 GND.n5148 GND.n5143 0.161
R6352 GND.n6327 GND.n491 0.161
R6353 GND.n5398 GND.n5397 0.157
R6354 GND.n2088 GND.n2087 0.157
R6355 GND.n5019 GND.n5018 0.157
R6356 GND.n4839 GND.n4838 0.157
R6357 GND.n4468 GND.n4467 0.157
R6358 GND.n5218 GND.n5217 0.157
R6359 GND.n1908 GND.n1907 0.157
R6360 GND.n3324 GND.n3323 0.157
R6361 GND.n5806 GND.n5805 0.157
R6362 GND.n5626 GND.n5625 0.157
R6363 GND.n3717 GND.n3716 0.157
R6364 GND.n4197 GND.n4196 0.157
R6365 GND.n2792 GND.n2791 0.157
R6366 GND.n3127 GND.n3126 0.157
R6367 GND.n1199 GND.n1198 0.157
R6368 GND.n730 GND.n729 0.157
R6369 GND.n1704 GND.n1703 0.157
R6370 GND.n1364 GND.n1363 0.157
R6371 GND.n1694 GND.n1686 0.15
R6372 GND.n1386 GND.n1378 0.15
R6373 GND.n1189 GND.n1181 0.15
R6374 GND.n752 GND.n744 0.15
R6375 GND.n2814 GND.n2806 0.15
R6376 GND.n3117 GND.n3109 0.15
R6377 GND.n3707 GND.n3699 0.15
R6378 GND.n1930 GND.n1922 0.15
R6379 GND.n2110 GND.n2102 0.15
R6380 GND.n5240 GND.n5232 0.15
R6381 GND.n5420 GND.n5412 0.15
R6382 GND.n4490 GND.n4482 0.15
R6383 GND.n4673 GND.n4664 0.15
R6384 GND.n4861 GND.n4853 0.15
R6385 GND.n5041 GND.n5033 0.15
R6386 GND.n3498 GND.n3490 0.15
R6387 GND.n3314 GND.n3306 0.15
R6388 GND.n5877 GND.n1825 0.15
R6389 GND.n5796 GND.n5788 0.15
R6390 GND.n5616 GND.n5608 0.15
R6391 GND.n5529 GND.n1838 0.15
R6392 GND.n4219 GND.n4211 0.15
R6393 GND.n8075 GND.n8074 0.149
R6394 GND.n2009 GND.n2006 0.146
R6395 GND.n5319 GND.n5316 0.146
R6396 GND.n4569 GND.n4566 0.146
R6397 GND.n4940 GND.n4937 0.146
R6398 GND.n3404 GND.n3402 0.146
R6399 GND.n5706 GND.n5704 0.146
R6400 GND.n2894 GND.n2893 0.146
R6401 GND.n1467 GND.n1466 0.146
R6402 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/SUBSTRATE GND.n1822 0.144
R6403 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/SUBSTRATE GND.n1809 0.144
R6404 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SUBSTRATE GND.n1796 0.144
R6405 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SUBSTRATE GND.n1783 0.144
R6406 GND.n3581 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/SUBSTRATE 0.144
R6407 GND.n5876 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/SUBSTRATE 0.144
R6408 GND.n4388 GND.n4387 0.142
R6409 GND.n4316 GND.n4315 0.142
R6410 GND.n4310 GND.n4309 0.142
R6411 GND.n2239 GND.n2238 0.142
R6412 GND.n6351 GND.n6350 0.142
R6413 GND.n6358 GND.n6357 0.142
R6414 GND.n474 GND.n473 0.142
R6415 GND.n6345 GND.n6344 0.142
R6416 GND.n6326 GND.n651 0.141
R6417 GND.n6138 GND.n944 0.141
R6418 GND.n6122 GND.n6121 0.141
R6419 GND.n3966 GND.n2566 0.141
R6420 GND.n3950 GND.n3949 0.141
R6421 GND.n4307 GND.n2417 0.141
R6422 GND.n3011 GND.n3010 0.141
R6423 GND.n4122 GND.n4121 0.141
R6424 GND.n1590 GND.n1589 0.141
R6425 GND.n6167 GND.n6165 0.141
R6426 GND.n5895 GND.n5894 0.137
R6427 GND.n6131 GND.n6128 0.132
R6428 GND.n6135 GND.n6131 0.132
R6429 GND.n3959 GND.n3956 0.132
R6430 GND.n3963 GND.n3959 0.132
R6431 GND.n2272 GND.n2263 0.132
R6432 GND.n2272 GND.n2269 0.132
R6433 GND.n506 GND.n497 0.132
R6434 GND.n506 GND.n503 0.132
R6435 GND.n3778 GND.n3608 0.128
R6436 GND.n612 GND.n610 0.127
R6437 GND.n619 GND.n617 0.127
R6438 GND.n626 GND.n624 0.127
R6439 GND.n633 GND.n631 0.127
R6440 GND.n640 GND.n638 0.127
R6441 GND.n647 GND.n645 0.127
R6442 GND.n1603 GND.n1601 0.127
R6443 GND.n1592 GND.n1288 0.127
R6444 GND.n6142 GND.n821 0.127
R6445 GND.n6163 GND.n6160 0.127
R6446 GND.n3015 GND.n2712 0.127
R6447 GND.n3026 GND.n3024 0.127
R6448 GND.n3970 GND.n2443 0.127
R6449 GND.n953 GND.n950 0.127
R6450 GND.n960 GND.n957 0.127
R6451 GND.n967 GND.n964 0.127
R6452 GND.n974 GND.n971 0.127
R6453 GND.n981 GND.n978 0.127
R6454 GND.n988 GND.n985 0.127
R6455 GND.n905 GND.n903 0.127
R6456 GND.n912 GND.n910 0.127
R6457 GND.n919 GND.n917 0.127
R6458 GND.n926 GND.n924 0.127
R6459 GND.n933 GND.n931 0.127
R6460 GND.n940 GND.n938 0.127
R6461 GND.n6082 GND.n6080 0.127
R6462 GND.n6089 GND.n6087 0.127
R6463 GND.n6096 GND.n6094 0.127
R6464 GND.n6103 GND.n6101 0.127
R6465 GND.n6110 GND.n6108 0.127
R6466 GND.n6117 GND.n6115 0.127
R6467 GND.n2575 GND.n2572 0.127
R6468 GND.n2582 GND.n2579 0.127
R6469 GND.n2589 GND.n2586 0.127
R6470 GND.n2596 GND.n2593 0.127
R6471 GND.n2603 GND.n2600 0.127
R6472 GND.n2610 GND.n2607 0.127
R6473 GND.n2527 GND.n2525 0.127
R6474 GND.n2534 GND.n2532 0.127
R6475 GND.n2541 GND.n2539 0.127
R6476 GND.n2548 GND.n2546 0.127
R6477 GND.n2555 GND.n2553 0.127
R6478 GND.n2562 GND.n2560 0.127
R6479 GND.n3910 GND.n3908 0.127
R6480 GND.n3917 GND.n3915 0.127
R6481 GND.n3924 GND.n3922 0.127
R6482 GND.n3931 GND.n3929 0.127
R6483 GND.n3938 GND.n3936 0.127
R6484 GND.n3945 GND.n3943 0.127
R6485 GND.n2378 GND.n2376 0.127
R6486 GND.n2385 GND.n2383 0.127
R6487 GND.n2392 GND.n2390 0.127
R6488 GND.n2399 GND.n2397 0.127
R6489 GND.n2406 GND.n2404 0.127
R6490 GND.n2413 GND.n2411 0.127
R6491 GND.n3006 GND.n3004 0.127
R6492 GND.n2999 GND.n2997 0.127
R6493 GND.n2992 GND.n2990 0.127
R6494 GND.n2985 GND.n2983 0.127
R6495 GND.n2978 GND.n2976 0.127
R6496 GND.n2971 GND.n2969 0.127
R6497 GND.n4117 GND.n4115 0.127
R6498 GND.n4110 GND.n4108 0.127
R6499 GND.n4103 GND.n4101 0.127
R6500 GND.n4096 GND.n4094 0.127
R6501 GND.n4089 GND.n4087 0.127
R6502 GND.n4082 GND.n4080 0.127
R6503 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/GATE GND.n4296 0.127
R6504 GND.n4128 GND.n4126 0.127
R6505 GND.n1585 GND.n1583 0.127
R6506 GND.n1578 GND.n1576 0.127
R6507 GND.n1571 GND.n1569 0.127
R6508 GND.n1564 GND.n1562 0.127
R6509 GND.n1557 GND.n1555 0.127
R6510 GND.n1550 GND.n1548 0.127
R6511 GND.n6174 GND.n6171 0.127
R6512 GND.n6181 GND.n6178 0.127
R6513 GND.n6188 GND.n6185 0.127
R6514 GND.n6195 GND.n6192 0.127
R6515 GND.n6202 GND.n6199 0.127
R6516 GND.n6209 GND.n6206 0.127
R6517 GND.n6316 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/GATE 0.127
R6518 GND.n6340 GND.n6339 0.125
R6519 GND.n5913 GND.n5912 0.125
R6520 GND.n2435 GND.n2434 0.118
R6521 GND.n458 GND.n457 0.116
R6522 GND.n2215 GND.n2214 0.114
R6523 GND.n4334 GND.n4333 0.114
R6524 GND.n1766 GND.n1758 0.114
R6525 GND.n1754 GND.n1746 0.114
R6526 GND.n1742 GND.n1734 0.114
R6527 GND.n1730 GND.n1722 0.114
R6528 GND.n1718 GND.n1710 0.114
R6529 GND.n1706 GND.n1698 0.114
R6530 GND.n1676 GND.n1674 0.114
R6531 GND.n1664 GND.n1662 0.114
R6532 GND.n1652 GND.n1650 0.114
R6533 GND.n1640 GND.n1638 0.114
R6534 GND.n1628 GND.n1626 0.114
R6535 GND.n1616 GND.n1614 0.114
R6536 GND.n1308 GND.n1306 0.114
R6537 GND.n1320 GND.n1318 0.114
R6538 GND.n1332 GND.n1330 0.114
R6539 GND.n1344 GND.n1342 0.114
R6540 GND.n1356 GND.n1354 0.114
R6541 GND.n1368 GND.n1366 0.114
R6542 GND.n1398 GND.n1390 0.114
R6543 GND.n1410 GND.n1402 0.114
R6544 GND.n1422 GND.n1414 0.114
R6545 GND.n1434 GND.n1426 0.114
R6546 GND.n1447 GND.n1438 0.114
R6547 GND.n1459 GND.n1451 0.114
R6548 GND.n1254 GND.n1253 0.114
R6549 GND.n1249 GND.n1241 0.114
R6550 GND.n1237 GND.n1229 0.114
R6551 GND.n1225 GND.n1217 0.114
R6552 GND.n1213 GND.n1205 0.114
R6553 GND.n1201 GND.n1193 0.114
R6554 GND.n1171 GND.n1169 0.114
R6555 GND.n1159 GND.n1157 0.114
R6556 GND.n1147 GND.n1145 0.114
R6557 GND.n1135 GND.n1133 0.114
R6558 GND.n1123 GND.n1121 0.114
R6559 GND.n1111 GND.n1109 0.114
R6560 GND.n686 GND.n684 0.114
R6561 GND.n698 GND.n696 0.114
R6562 GND.n710 GND.n708 0.114
R6563 GND.n722 GND.n720 0.114
R6564 GND.n734 GND.n732 0.114
R6565 GND.n764 GND.n756 0.114
R6566 GND.n776 GND.n768 0.114
R6567 GND.n788 GND.n780 0.114
R6568 GND.n800 GND.n792 0.114
R6569 GND.n812 GND.n804 0.114
R6570 GND.n817 GND.n816 0.114
R6571 GND.n2736 GND.n2734 0.114
R6572 GND.n2748 GND.n2746 0.114
R6573 GND.n2760 GND.n2758 0.114
R6574 GND.n2772 GND.n2770 0.114
R6575 GND.n2784 GND.n2782 0.114
R6576 GND.n2796 GND.n2794 0.114
R6577 GND.n2826 GND.n2818 0.114
R6578 GND.n2838 GND.n2830 0.114
R6579 GND.n2850 GND.n2842 0.114
R6580 GND.n2862 GND.n2854 0.114
R6581 GND.n2874 GND.n2866 0.114
R6582 GND.n2886 GND.n2878 0.114
R6583 GND.n3189 GND.n3181 0.114
R6584 GND.n3177 GND.n3169 0.114
R6585 GND.n3165 GND.n3157 0.114
R6586 GND.n3153 GND.n3145 0.114
R6587 GND.n3141 GND.n3133 0.114
R6588 GND.n3129 GND.n3121 0.114
R6589 GND.n3099 GND.n3097 0.114
R6590 GND.n3087 GND.n3085 0.114
R6591 GND.n3075 GND.n3073 0.114
R6592 GND.n3063 GND.n3061 0.114
R6593 GND.n3051 GND.n3049 0.114
R6594 GND.n3039 GND.n3037 0.114
R6595 GND.n3772 GND.n3771 0.114
R6596 GND.n3767 GND.n3759 0.114
R6597 GND.n3755 GND.n3747 0.114
R6598 GND.n3743 GND.n3735 0.114
R6599 GND.n3731 GND.n3723 0.114
R6600 GND.n3719 GND.n3711 0.114
R6601 GND.n3689 GND.n3687 0.114
R6602 GND.n3677 GND.n3675 0.114
R6603 GND.n3665 GND.n3663 0.114
R6604 GND.n3653 GND.n3651 0.114
R6605 GND.n3641 GND.n3639 0.114
R6606 GND.n3629 GND.n3627 0.114
R6607 GND.n1852 GND.n1850 0.114
R6608 GND.n1864 GND.n1862 0.114
R6609 GND.n1876 GND.n1874 0.114
R6610 GND.n1888 GND.n1886 0.114
R6611 GND.n1900 GND.n1898 0.114
R6612 GND.n1912 GND.n1910 0.114
R6613 GND.n1942 GND.n1934 0.114
R6614 GND.n1954 GND.n1946 0.114
R6615 GND.n1966 GND.n1958 0.114
R6616 GND.n1978 GND.n1970 0.114
R6617 GND.n1990 GND.n1982 0.114
R6618 GND.n2002 GND.n1994 0.114
R6619 GND.n2032 GND.n2030 0.114
R6620 GND.n2044 GND.n2042 0.114
R6621 GND.n2056 GND.n2054 0.114
R6622 GND.n2068 GND.n2066 0.114
R6623 GND.n2080 GND.n2078 0.114
R6624 GND.n2092 GND.n2090 0.114
R6625 GND.n2122 GND.n2114 0.114
R6626 GND.n2134 GND.n2126 0.114
R6627 GND.n2146 GND.n2138 0.114
R6628 GND.n2158 GND.n2150 0.114
R6629 GND.n2170 GND.n2162 0.114
R6630 GND.n2175 GND.n2174 0.114
R6631 GND.n5162 GND.n5160 0.114
R6632 GND.n5174 GND.n5172 0.114
R6633 GND.n5186 GND.n5184 0.114
R6634 GND.n5198 GND.n5196 0.114
R6635 GND.n5210 GND.n5208 0.114
R6636 GND.n5222 GND.n5220 0.114
R6637 GND.n5252 GND.n5244 0.114
R6638 GND.n5264 GND.n5256 0.114
R6639 GND.n5276 GND.n5268 0.114
R6640 GND.n5288 GND.n5280 0.114
R6641 GND.n5300 GND.n5292 0.114
R6642 GND.n5312 GND.n5304 0.114
R6643 GND.n5342 GND.n5340 0.114
R6644 GND.n5354 GND.n5352 0.114
R6645 GND.n5366 GND.n5364 0.114
R6646 GND.n5378 GND.n5376 0.114
R6647 GND.n5390 GND.n5388 0.114
R6648 GND.n5402 GND.n5400 0.114
R6649 GND.n5432 GND.n5424 0.114
R6650 GND.n5444 GND.n5436 0.114
R6651 GND.n5456 GND.n5448 0.114
R6652 GND.n5468 GND.n5460 0.114
R6653 GND.n5480 GND.n5472 0.114
R6654 GND.n5485 GND.n5484 0.114
R6655 GND.n4412 GND.n4410 0.114
R6656 GND.n4424 GND.n4422 0.114
R6657 GND.n4436 GND.n4434 0.114
R6658 GND.n4448 GND.n4446 0.114
R6659 GND.n4460 GND.n4458 0.114
R6660 GND.n4472 GND.n4470 0.114
R6661 GND.n4502 GND.n4494 0.114
R6662 GND.n4514 GND.n4506 0.114
R6663 GND.n4526 GND.n4518 0.114
R6664 GND.n4538 GND.n4530 0.114
R6665 GND.n4550 GND.n4542 0.114
R6666 GND.n4562 GND.n4554 0.114
R6667 GND.n4592 GND.n4590 0.114
R6668 GND.n4604 GND.n4602 0.114
R6669 GND.n4616 GND.n4614 0.114
R6670 GND.n4629 GND.n4627 0.114
R6671 GND.n4641 GND.n4639 0.114
R6672 GND.n4654 GND.n4652 0.114
R6673 GND.n4686 GND.n4677 0.114
R6674 GND.n4698 GND.n4690 0.114
R6675 GND.n4711 GND.n4702 0.114
R6676 GND.n4723 GND.n4715 0.114
R6677 GND.n4736 GND.n4727 0.114
R6678 GND.n4741 GND.n4740 0.114
R6679 GND.n4783 GND.n4781 0.114
R6680 GND.n4795 GND.n4793 0.114
R6681 GND.n4807 GND.n4805 0.114
R6682 GND.n4819 GND.n4817 0.114
R6683 GND.n4831 GND.n4829 0.114
R6684 GND.n4843 GND.n4841 0.114
R6685 GND.n4873 GND.n4865 0.114
R6686 GND.n4885 GND.n4877 0.114
R6687 GND.n4897 GND.n4889 0.114
R6688 GND.n4909 GND.n4901 0.114
R6689 GND.n4921 GND.n4913 0.114
R6690 GND.n4933 GND.n4925 0.114
R6691 GND.n4963 GND.n4961 0.114
R6692 GND.n4975 GND.n4973 0.114
R6693 GND.n4987 GND.n4985 0.114
R6694 GND.n4999 GND.n4997 0.114
R6695 GND.n5011 GND.n5009 0.114
R6696 GND.n5023 GND.n5021 0.114
R6697 GND.n5053 GND.n5045 0.114
R6698 GND.n5065 GND.n5057 0.114
R6699 GND.n5077 GND.n5069 0.114
R6700 GND.n5089 GND.n5081 0.114
R6701 GND.n5101 GND.n5093 0.114
R6702 GND.n5106 GND.n5105 0.114
R6703 GND.n3566 GND.n3565 0.114
R6704 GND.n3561 GND.n3552 0.114
R6705 GND.n3548 GND.n3540 0.114
R6706 GND.n3536 GND.n3527 0.114
R6707 GND.n3523 GND.n3515 0.114
R6708 GND.n3511 GND.n3502 0.114
R6709 GND.n3479 GND.n3477 0.114
R6710 GND.n3466 GND.n3464 0.114
R6711 GND.n3454 GND.n3452 0.114
R6712 GND.n3441 GND.n3439 0.114
R6713 GND.n3429 GND.n3427 0.114
R6714 GND.n3416 GND.n3414 0.114
R6715 GND.n3386 GND.n3378 0.114
R6716 GND.n3374 GND.n3366 0.114
R6717 GND.n3362 GND.n3354 0.114
R6718 GND.n3350 GND.n3342 0.114
R6719 GND.n3338 GND.n3330 0.114
R6720 GND.n3326 GND.n3318 0.114
R6721 GND.n3296 GND.n3294 0.114
R6722 GND.n3284 GND.n3282 0.114
R6723 GND.n3272 GND.n3270 0.114
R6724 GND.n3260 GND.n3258 0.114
R6725 GND.n3248 GND.n3246 0.114
R6726 GND.n3235 GND.n3233 0.114
R6727 GND.n5861 GND.n5860 0.114
R6728 GND.n5856 GND.n5848 0.114
R6729 GND.n5844 GND.n5836 0.114
R6730 GND.n5832 GND.n5824 0.114
R6731 GND.n5820 GND.n5812 0.114
R6732 GND.n5808 GND.n5800 0.114
R6733 GND.n5778 GND.n5776 0.114
R6734 GND.n5766 GND.n5764 0.114
R6735 GND.n5754 GND.n5752 0.114
R6736 GND.n5742 GND.n5740 0.114
R6737 GND.n5730 GND.n5728 0.114
R6738 GND.n5718 GND.n5716 0.114
R6739 GND.n5688 GND.n5680 0.114
R6740 GND.n5676 GND.n5668 0.114
R6741 GND.n5664 GND.n5656 0.114
R6742 GND.n5652 GND.n5644 0.114
R6743 GND.n5640 GND.n5632 0.114
R6744 GND.n5628 GND.n5620 0.114
R6745 GND.n5598 GND.n5596 0.114
R6746 GND.n5586 GND.n5584 0.114
R6747 GND.n5574 GND.n5572 0.114
R6748 GND.n5562 GND.n5560 0.114
R6749 GND.n5550 GND.n5548 0.114
R6750 GND.n5537 GND.n5535 0.114
R6751 GND.n4141 GND.n4139 0.114
R6752 GND.n4153 GND.n4151 0.114
R6753 GND.n4165 GND.n4163 0.114
R6754 GND.n4177 GND.n4175 0.114
R6755 GND.n4189 GND.n4187 0.114
R6756 GND.n4201 GND.n4199 0.114
R6757 GND.n4231 GND.n4223 0.114
R6758 GND.n4243 GND.n4235 0.114
R6759 GND.n4255 GND.n4247 0.114
R6760 GND.n4267 GND.n4259 0.114
R6761 GND.n4279 GND.n4271 0.114
R6762 GND.n4291 GND.n4283 0.114
R6763 GND.n5134 GND.n5131 0.112
R6764 GND.n5931 GND.n5930 0.112
R6765 GND.n2181 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SUBSTRATE 0.109
R6766 GND.n5491 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/SUBSTRATE 0.109
R6767 GND.n4747 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SUBSTRATE 0.109
R6768 GND.n5112 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SUBSTRATE 0.109
R6769 GND.n3228 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/SUBSTRATE 0.109
R6770 GND.n5530 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SUBSTRATE 0.109
R6771 GND.n5969 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/SUBSTRATE 0.107
R6772 GND.n1260 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/SUBSTRATE 0.107
R6773 GND.n3196 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/SUBSTRATE 0.107
R6774 GND.n3778 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/SUBSTRATE 0.107
R6775 GND.n507 GND.n506 0.103
R6776 GND.n6131 GND.n1087 0.103
R6777 GND.n5976 GND.n5975 0.103
R6778 GND.n3959 GND.n2709 0.103
R6779 GND.n3804 GND.n3803 0.103
R6780 GND.n2273 GND.n2272 0.103
R6781 GND.n2898 GND.n2897 0.103
R6782 GND.n4298 GND.n2422 0.103
R6783 GND.n1471 GND.n1470 0.103
R6784 GND.n6314 GND.n6311 0.103
R6785 GND.n5116 GND.n5113 0.099
R6786 GND.n5949 GND.n5948 0.099
R6787 GND.n8074 GND.n8073 0.095
R6788 GND.n6611 GND.n6607 0.095
R6789 GND.n8056 GND.n8055 0.095
R6790 GND.n6628 GND.n6624 0.095
R6791 GND.n7829 GND.n7828 0.095
R6792 GND.n6645 GND.n6641 0.095
R6793 GND.n7602 GND.n7601 0.095
R6794 GND.n6662 GND.n6658 0.095
R6795 GND.n7375 GND.n7374 0.095
R6796 GND.n6679 GND.n6675 0.095
R6797 GND.n7148 GND.n7147 0.095
R6798 GND.n6696 GND.n6692 0.095
R6799 GND.n6921 GND.n6920 0.095
R6800 GND.n451 GND.n450 0.095
R6801 GND.n8491 GND.n8490 0.095
R6802 GND.n402 GND.n401 0.095
R6803 GND.n8676 GND.n8675 0.095
R6804 GND.n353 GND.n352 0.095
R6805 GND.n8861 GND.n8860 0.095
R6806 GND.n304 GND.n303 0.095
R6807 GND.n9046 GND.n9045 0.095
R6808 GND.n255 GND.n254 0.095
R6809 GND.n9231 GND.n9230 0.095
R6810 GND.n9252 GND.n9251 0.095
R6811 GND.n228 GND.n225 0.095
R6812 GND.n277 GND.n274 0.095
R6813 GND.n326 GND.n323 0.095
R6814 GND.n375 GND.n372 0.095
R6815 GND.n424 GND.n421 0.095
R6816 GND.n6898 GND.n6897 0.095
R6817 GND.n7125 GND.n7124 0.095
R6818 GND.n7352 GND.n7351 0.095
R6819 GND.n7579 GND.n7578 0.095
R6820 GND.n7806 GND.n7805 0.095
R6821 GND.n8033 GND.n8032 0.095
R6822 GND.n5514 GND.n5511 0.094
R6823 GND.n4307 GND.n2421 0.093
R6824 GND.n4307 GND.n4304 0.093
R6825 GND.n6326 GND.n655 0.093
R6826 GND.n6326 GND.n661 0.093
R6827 GND.n1021 GND.n1000 0.092
R6828 GND.n2643 GND.n2622 0.092
R6829 GND.n1466 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/SUBSTRATE 0.073
R6830 GND.n6316 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/SUBSTRATE 0.073
R6831 GND.n2893 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/SUBSTRATE 0.073
R6832 GND.n5113 GND.n4769 0.073
R6833 GND.n5954 GND.n5949 0.073
R6834 GND.n4296 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/SUBSTRATE 0.073
R6835 GND.n1595 GND.n1592 0.066
R6836 GND.n6163 GND.n6148 0.066
R6837 GND.n3018 GND.n3015 0.066
R6838 GND.n4126 GND.n3976 0.066
R6839 GND.n3786 GND.n3783 0.065
R6840 GND.n4343 GND.n4342 0.063
R6841 GND.n7916 GND.n7915 0.06
R6842 GND.n7689 GND.n7688 0.06
R6843 GND.n7462 GND.n7461 0.06
R6844 GND.n7235 GND.n7234 0.06
R6845 GND.n7008 GND.n7007 0.06
R6846 GND.n6781 GND.n6780 0.06
R6847 GND.n6460 GND.n6459 0.06
R6848 GND.n516 GND.n515 0.06
R6849 GND.n526 GND.n525 0.06
R6850 GND.n537 GND.n536 0.06
R6851 GND.n548 GND.n547 0.06
R6852 GND.n1048 GND.n1046 0.06
R6853 GND.n1059 GND.n1057 0.06
R6854 GND.n1069 GND.n1068 0.06
R6855 GND.n1079 GND.n1078 0.06
R6856 GND.n831 GND.n830 0.06
R6857 GND.n841 GND.n840 0.06
R6858 GND.n852 GND.n851 0.06
R6859 GND.n863 GND.n862 0.06
R6860 GND.n5985 GND.n5984 0.06
R6861 GND.n5995 GND.n5994 0.06
R6862 GND.n6006 GND.n6005 0.06
R6863 GND.n6017 GND.n6016 0.06
R6864 GND.n2670 GND.n2668 0.06
R6865 GND.n2681 GND.n2679 0.06
R6866 GND.n2691 GND.n2690 0.06
R6867 GND.n2701 GND.n2700 0.06
R6868 GND.n2453 GND.n2452 0.06
R6869 GND.n2463 GND.n2462 0.06
R6870 GND.n2474 GND.n2473 0.06
R6871 GND.n2485 GND.n2484 0.06
R6872 GND.n3813 GND.n3812 0.06
R6873 GND.n3823 GND.n3822 0.06
R6874 GND.n3834 GND.n3833 0.06
R6875 GND.n3845 GND.n3844 0.06
R6876 GND.n5131 GND.n5130 0.06
R6877 GND.n5936 GND.n5931 0.06
R6878 GND.n2282 GND.n2281 0.06
R6879 GND.n2292 GND.n2291 0.06
R6880 GND.n2303 GND.n2302 0.06
R6881 GND.n2314 GND.n2313 0.06
R6882 GND.n2935 GND.n2934 0.06
R6883 GND.n2925 GND.n2924 0.06
R6884 GND.n2915 GND.n2914 0.06
R6885 GND.n2906 GND.n2905 0.06
R6886 GND.n4046 GND.n4045 0.06
R6887 GND.n4036 GND.n4035 0.06
R6888 GND.n4026 GND.n4025 0.06
R6889 GND.n4017 GND.n4016 0.06
R6890 GND.n1509 GND.n1508 0.06
R6891 GND.n1498 GND.n1497 0.06
R6892 GND.n1488 GND.n1487 0.06
R6893 GND.n1479 GND.n1478 0.06
R6894 GND.n6249 GND.n6247 0.06
R6895 GND.n6260 GND.n6258 0.06
R6896 GND.n6270 GND.n6269 0.06
R6897 GND.n6280 GND.n6279 0.06
R6898 GND.n8225 GND.n8224 0.06
R6899 GND.n8153 GND.n8152 0.06
R6900 GND.n8332 GND.n8331 0.06
R6901 GND.n8404 GND.n8403 0.06
R6902 GND.n8517 GND.n8516 0.06
R6903 GND.n8589 GND.n8588 0.06
R6904 GND.n8702 GND.n8701 0.06
R6905 GND.n8774 GND.n8773 0.06
R6906 GND.n8887 GND.n8886 0.06
R6907 GND.n8959 GND.n8958 0.06
R6908 GND.n9072 GND.n9071 0.06
R6909 GND.n9144 GND.n9143 0.06
R6910 GND.n33 GND.n32 0.06
R6911 GND.n105 GND.n104 0.06
R6912 GND.n3199 GND.n3196 0.059
R6913 GND.n462 GND.n461 0.059
R6914 GND.n4384 GND.n4383 0.059
R6915 GND.n4355 GND.n4354 0.059
R6916 GND.n6359 GND.n6358 0.059
R6917 GND.n475 GND.n474 0.059
R6918 GND.n2223 GND.n2222 0.059
R6919 GND.n2240 GND.n2239 0.059
R6920 GND.n4317 GND.n4316 0.059
R6921 GND.n4338 GND.n4325 0.059
R6922 GND.n4336 GND.n4335 0.059
R6923 GND.n2217 GND.n2216 0.059
R6924 GND.n5975 GND.n5974 0.057
R6925 GND.n1281 GND.n1277 0.057
R6926 GND.n8076 GND.n8075 0.056
R6927 GND.n1274 GND.n1271 0.055
R6928 GND.n5510 GND.n5505 0.054
R6929 GND.n5505 GND.n5502 0.054
R6930 GND.n5498 GND.n5495 0.054
R6931 GND.n561 GND.n560 0.053
R6932 GND.n566 GND.n561 0.053
R6933 GND.n1033 GND.n1032 0.053
R6934 GND.n1035 GND.n1033 0.053
R6935 GND.n876 GND.n875 0.053
R6936 GND.n881 GND.n876 0.053
R6937 GND.n6030 GND.n6029 0.053
R6938 GND.n6035 GND.n6030 0.053
R6939 GND.n2655 GND.n2654 0.053
R6940 GND.n2657 GND.n2655 0.053
R6941 GND.n2498 GND.n2497 0.053
R6942 GND.n2503 GND.n2498 0.053
R6943 GND.n3858 GND.n3857 0.053
R6944 GND.n3863 GND.n3858 0.053
R6945 GND.n2327 GND.n2326 0.053
R6946 GND.n2332 GND.n2327 0.053
R6947 GND.n2948 GND.n2947 0.053
R6948 GND.n2947 GND.n2946 0.053
R6949 GND.n4059 GND.n4058 0.053
R6950 GND.n4058 GND.n4057 0.053
R6951 GND.n1527 GND.n1521 0.053
R6952 GND.n1521 GND.n1520 0.053
R6953 GND.n6234 GND.n6233 0.053
R6954 GND.n6236 GND.n6234 0.053
R6955 GND.n5410 GND.n5409 0.053
R6956 GND.n2100 GND.n2099 0.053
R6957 GND.n4662 GND.n4661 0.053
R6958 GND.n4671 GND.n4670 0.053
R6959 GND.n5031 GND.n5030 0.053
R6960 GND.n4851 GND.n4850 0.053
R6961 GND.n4480 GND.n4479 0.053
R6962 GND.n5230 GND.n5229 0.053
R6963 GND.n1920 GND.n1919 0.053
R6964 GND.n3496 GND.n3495 0.053
R6965 GND.n3488 GND.n3487 0.053
R6966 GND.n3312 GND.n3311 0.053
R6967 GND.n5794 GND.n5793 0.053
R6968 GND.n5614 GND.n5613 0.053
R6969 GND.n3705 GND.n3704 0.053
R6970 GND.n4209 GND.n4208 0.053
R6971 GND.n2804 GND.n2803 0.053
R6972 GND.n3115 GND.n3114 0.053
R6973 GND.n1187 GND.n1186 0.053
R6974 GND.n742 GND.n741 0.053
R6975 GND.n1692 GND.n1691 0.053
R6976 GND.n1376 GND.n1375 0.053
R6977 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/SUBSTRATE GND.n1463 0.053
R6978 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/SUBSTRATE GND.n819 0.053
R6979 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/SUBSTRATE GND.n2890 0.053
R6980 GND.n2177 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SUBSTRATE 0.053
R6981 GND.n5487 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/SUBSTRATE 0.053
R6982 GND.n4743 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SUBSTRATE 0.053
R6983 GND.n5108 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SUBSTRATE 0.053
R6984 GND.n3231 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/SUBSTRATE 0.053
R6985 GND.n5533 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SUBSTRATE 0.053
R6986 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/SUBSTRATE GND.n4295 0.053
R6987 GND.n8251 GND.n8248 0.052
R6988 GND.n8179 GND.n8176 0.052
R6989 GND.n8358 GND.n8355 0.052
R6990 GND.n8430 GND.n8427 0.052
R6991 GND.n8543 GND.n8540 0.052
R6992 GND.n8615 GND.n8612 0.052
R6993 GND.n8728 GND.n8725 0.052
R6994 GND.n8800 GND.n8797 0.052
R6995 GND.n8913 GND.n8910 0.052
R6996 GND.n8985 GND.n8982 0.052
R6997 GND.n9098 GND.n9095 0.052
R6998 GND.n9170 GND.n9167 0.052
R6999 GND.n59 GND.n56 0.052
R7000 GND.n131 GND.n128 0.052
R7001 GND.n2425 GND.n2252 0.051
R7002 GND.n2435 GND.n2425 0.051
R7003 GND.n598 GND.n595 0.05
R7004 GND.n891 GND.n888 0.05
R7005 GND.n6068 GND.n6065 0.05
R7006 GND.n1261 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/GATE 0.05
R7007 GND.n2513 GND.n2510 0.05
R7008 GND.n3896 GND.n3893 0.05
R7009 GND.n2364 GND.n2361 0.05
R7010 GND.n2957 GND.n2954 0.05
R7011 GND.n4068 GND.n4065 0.05
R7012 GND.n1536 GND.n1533 0.05
R7013 GND.n6222 GND.n6221 0.05
R7014 GND.n8247 GND.n8246 0.05
R7015 GND.n8175 GND.n8174 0.05
R7016 GND.n8354 GND.n8353 0.05
R7017 GND.n8426 GND.n8425 0.05
R7018 GND.n8539 GND.n8538 0.05
R7019 GND.n8611 GND.n8610 0.05
R7020 GND.n8724 GND.n8723 0.05
R7021 GND.n8796 GND.n8795 0.05
R7022 GND.n8909 GND.n8908 0.05
R7023 GND.n8981 GND.n8980 0.05
R7024 GND.n9094 GND.n9093 0.05
R7025 GND.n9166 GND.n9165 0.05
R7026 GND.n55 GND.n54 0.05
R7027 GND.n127 GND.n126 0.05
R7028 GND.n2208 GND.n2207 0.05
R7029 GND.n1601 GND.n1598 0.049
R7030 GND.n6145 GND.n6142 0.049
R7031 GND.n3024 GND.n3021 0.049
R7032 GND.n3973 GND.n3970 0.049
R7033 GND.n7945 GND.n7940 0.048
R7034 GND.n7951 GND.n7950 0.048
R7035 GND.n7718 GND.n7713 0.048
R7036 GND.n7724 GND.n7723 0.048
R7037 GND.n7491 GND.n7486 0.048
R7038 GND.n7497 GND.n7496 0.048
R7039 GND.n7264 GND.n7259 0.048
R7040 GND.n7270 GND.n7269 0.048
R7041 GND.n7037 GND.n7032 0.048
R7042 GND.n7043 GND.n7042 0.048
R7043 GND.n6810 GND.n6805 0.048
R7044 GND.n6816 GND.n6815 0.048
R7045 GND.n6478 GND.n6473 0.048
R7046 GND.n6484 GND.n6483 0.048
R7047 GND.n480 GND.n479 0.048
R7048 GND.n8307 GND.n8306 0.048
R7049 GND.n8066 GND.n8065 0.048
R7050 GND.n4350 GND.n4349 0.048
R7051 GND.n4381 GND.n4380 0.048
R7052 GND.n4376 GND.n486 0.048
R7053 GND.n2224 GND.n2223 0.048
R7054 GND.n4339 GND.n4338 0.048
R7055 GND.n5918 GND.n5913 0.047
R7056 GND.n5969 GND.n5966 0.046
R7057 GND.n7983 GND.n7976 0.043
R7058 GND.n7987 GND.n7986 0.043
R7059 GND.n7756 GND.n7749 0.043
R7060 GND.n7760 GND.n7759 0.043
R7061 GND.n7529 GND.n7522 0.043
R7062 GND.n7533 GND.n7532 0.043
R7063 GND.n7302 GND.n7295 0.043
R7064 GND.n7306 GND.n7305 0.043
R7065 GND.n7075 GND.n7068 0.043
R7066 GND.n7079 GND.n7078 0.043
R7067 GND.n6848 GND.n6841 0.043
R7068 GND.n6852 GND.n6851 0.043
R7069 GND.n6516 GND.n6509 0.043
R7070 GND.n6520 GND.n6519 0.043
R7071 GND.n519 GND.n516 0.043
R7072 GND.n594 GND.n593 0.043
R7073 GND.n1078 GND.n1077 0.043
R7074 GND.n834 GND.n831 0.043
R7075 GND.n887 GND.n886 0.043
R7076 GND.n5988 GND.n5985 0.043
R7077 GND.n6064 GND.n6063 0.043
R7078 GND.n2700 GND.n2699 0.043
R7079 GND.n2456 GND.n2453 0.043
R7080 GND.n2509 GND.n2508 0.043
R7081 GND.n3816 GND.n3813 0.043
R7082 GND.n3892 GND.n3891 0.043
R7083 GND.n2285 GND.n2282 0.043
R7084 GND.n2360 GND.n2359 0.043
R7085 GND.n2953 GND.n2952 0.043
R7086 GND.n2909 GND.n2906 0.043
R7087 GND.n4064 GND.n4063 0.043
R7088 GND.n4020 GND.n4017 0.043
R7089 GND.n1532 GND.n1531 0.043
R7090 GND.n1482 GND.n1479 0.043
R7091 GND.n6225 GND.n6223 0.043
R7092 GND.n6279 GND.n6278 0.043
R7093 GND.n8237 GND.n8236 0.043
R7094 GND.n8165 GND.n8164 0.043
R7095 GND.n8344 GND.n8343 0.043
R7096 GND.n8416 GND.n8415 0.043
R7097 GND.n8529 GND.n8528 0.043
R7098 GND.n8601 GND.n8600 0.043
R7099 GND.n8714 GND.n8713 0.043
R7100 GND.n8786 GND.n8785 0.043
R7101 GND.n8899 GND.n8898 0.043
R7102 GND.n8971 GND.n8970 0.043
R7103 GND.n9084 GND.n9083 0.043
R7104 GND.n9156 GND.n9155 0.043
R7105 GND.n45 GND.n44 0.043
R7106 GND.n117 GND.n116 0.043
R7107 GND.n6328 GND.n6327 0.042
R7108 GND.n8235 GND.n8234 0.041
R7109 GND.n8163 GND.n8162 0.041
R7110 GND.n8342 GND.n8341 0.041
R7111 GND.n8414 GND.n8413 0.041
R7112 GND.n8527 GND.n8526 0.041
R7113 GND.n8599 GND.n8598 0.041
R7114 GND.n8712 GND.n8711 0.041
R7115 GND.n8784 GND.n8783 0.041
R7116 GND.n8897 GND.n8896 0.041
R7117 GND.n8969 GND.n8968 0.041
R7118 GND.n9082 GND.n9081 0.041
R7119 GND.n9154 GND.n9153 0.041
R7120 GND.n43 GND.n42 0.041
R7121 GND.n115 GND.n114 0.041
R7122 GND.n8012 GND.n8011 0.04
R7123 GND.n7999 GND.n7998 0.04
R7124 GND.n7785 GND.n7784 0.04
R7125 GND.n7772 GND.n7771 0.04
R7126 GND.n7558 GND.n7557 0.04
R7127 GND.n7545 GND.n7544 0.04
R7128 GND.n7331 GND.n7330 0.04
R7129 GND.n7318 GND.n7317 0.04
R7130 GND.n7104 GND.n7103 0.04
R7131 GND.n7091 GND.n7090 0.04
R7132 GND.n6877 GND.n6876 0.04
R7133 GND.n6864 GND.n6863 0.04
R7134 GND.n6545 GND.n6544 0.04
R7135 GND.n6532 GND.n6531 0.04
R7136 GND.n552 GND.n549 0.04
R7137 GND.n1045 GND.n1044 0.04
R7138 GND.n867 GND.n864 0.04
R7139 GND.n6021 GND.n6018 0.04
R7140 GND.n2667 GND.n2666 0.04
R7141 GND.n2489 GND.n2486 0.04
R7142 GND.n3849 GND.n3846 0.04
R7143 GND.n5499 GND.n5498 0.04
R7144 GND.n2318 GND.n2315 0.04
R7145 GND.n2939 GND.n2936 0.04
R7146 GND.n4050 GND.n4047 0.04
R7147 GND.n1513 GND.n1510 0.04
R7148 GND.n6246 GND.n6245 0.04
R7149 GND.n8263 GND.n8260 0.04
R7150 GND.n8191 GND.n8188 0.04
R7151 GND.n8370 GND.n8367 0.04
R7152 GND.n8442 GND.n8439 0.04
R7153 GND.n8555 GND.n8552 0.04
R7154 GND.n8627 GND.n8624 0.04
R7155 GND.n8740 GND.n8737 0.04
R7156 GND.n8812 GND.n8809 0.04
R7157 GND.n8925 GND.n8922 0.04
R7158 GND.n8997 GND.n8994 0.04
R7159 GND.n9110 GND.n9107 0.04
R7160 GND.n9182 GND.n9179 0.04
R7161 GND.n71 GND.n68 0.04
R7162 GND.n143 GND.n140 0.04
R7163 GND.n4377 GND 0.04
R7164 GND.n5495 GND.n5492 0.039
R7165 GND.n8019 GND.n8017 0.038
R7166 GND.n7792 GND.n7790 0.038
R7167 GND.n7565 GND.n7563 0.038
R7168 GND.n7338 GND.n7336 0.038
R7169 GND.n7111 GND.n7109 0.038
R7170 GND.n6884 GND.n6882 0.038
R7171 GND.n6552 GND.n6550 0.038
R7172 GND.n509 GND.n507 0.038
R7173 GND.n600 GND.n598 0.038
R7174 GND.n610 GND.n607 0.038
R7175 GND.n990 GND.n988 0.038
R7176 GND.n1000 GND.n997 0.038
R7177 GND.n1087 GND.n1086 0.038
R7178 GND.n824 GND.n822 0.038
R7179 GND.n893 GND.n891 0.038
R7180 GND.n903 GND.n900 0.038
R7181 GND.n5978 GND.n5976 0.038
R7182 GND.n6070 GND.n6068 0.038
R7183 GND.n6080 GND.n6077 0.038
R7184 GND.n2612 GND.n2610 0.038
R7185 GND.n2622 GND.n2619 0.038
R7186 GND.n2709 GND.n2708 0.038
R7187 GND.n2446 GND.n2444 0.038
R7188 GND.n2515 GND.n2513 0.038
R7189 GND.n2525 GND.n2522 0.038
R7190 GND.n3806 GND.n3804 0.038
R7191 GND.n3898 GND.n3896 0.038
R7192 GND.n3908 GND.n3905 0.038
R7193 GND.n2275 GND.n2273 0.038
R7194 GND.n2366 GND.n2364 0.038
R7195 GND.n2376 GND.n2373 0.038
R7196 GND.n2969 GND.n2966 0.038
R7197 GND.n2959 GND.n2957 0.038
R7198 GND.n2900 GND.n2898 0.038
R7199 GND.n4080 GND.n4077 0.038
R7200 GND.n4070 GND.n4068 0.038
R7201 GND.n3988 GND.n2422 0.038
R7202 GND.n1548 GND.n1545 0.038
R7203 GND.n1538 GND.n1536 0.038
R7204 GND.n1473 GND.n1471 0.038
R7205 GND.n6211 GND.n6209 0.038
R7206 GND.n6221 GND.n6218 0.038
R7207 GND.n6311 GND.n6310 0.038
R7208 GND.n8226 GND.n8225 0.038
R7209 GND.n8154 GND.n8153 0.038
R7210 GND.n8333 GND.n8332 0.038
R7211 GND.n8405 GND.n8404 0.038
R7212 GND.n8518 GND.n8517 0.038
R7213 GND.n8590 GND.n8589 0.038
R7214 GND.n8703 GND.n8702 0.038
R7215 GND.n8775 GND.n8774 0.038
R7216 GND.n8888 GND.n8887 0.038
R7217 GND.n8960 GND.n8959 0.038
R7218 GND.n9073 GND.n9072 0.038
R7219 GND.n9145 GND.n9144 0.038
R7220 GND.n34 GND.n33 0.038
R7221 GND.n106 GND.n105 0.038
R7222 GND.n3799 GND.n3796 0.037
R7223 GND.n527 GND.n526 0.036
R7224 GND.n1068 GND.n1067 0.036
R7225 GND.n842 GND.n841 0.036
R7226 GND.n5996 GND.n5995 0.036
R7227 GND.n2690 GND.n2689 0.036
R7228 GND.n2464 GND.n2463 0.036
R7229 GND.n3824 GND.n3823 0.036
R7230 GND.n2293 GND.n2292 0.036
R7231 GND.n2916 GND.n2915 0.036
R7232 GND.n4027 GND.n4026 0.036
R7233 GND.n1489 GND.n1488 0.036
R7234 GND.n6269 GND.n6268 0.036
R7235 GND.n8275 GND.n8274 0.036
R7236 GND.n8273 GND.n8272 0.036
R7237 GND.n8202 GND.n8200 0.036
R7238 GND.n8199 GND.n8198 0.036
R7239 GND.n8382 GND.n8381 0.036
R7240 GND.n8380 GND.n8379 0.036
R7241 GND.n8453 GND.n8452 0.036
R7242 GND.n8451 GND.n8450 0.036
R7243 GND.n8567 GND.n8566 0.036
R7244 GND.n8565 GND.n8564 0.036
R7245 GND.n8638 GND.n8637 0.036
R7246 GND.n8636 GND.n8635 0.036
R7247 GND.n8752 GND.n8751 0.036
R7248 GND.n8750 GND.n8749 0.036
R7249 GND.n8823 GND.n8822 0.036
R7250 GND.n8821 GND.n8820 0.036
R7251 GND.n8937 GND.n8936 0.036
R7252 GND.n8935 GND.n8934 0.036
R7253 GND.n9008 GND.n9007 0.036
R7254 GND.n9006 GND.n9005 0.036
R7255 GND.n9122 GND.n9121 0.036
R7256 GND.n9120 GND.n9119 0.036
R7257 GND.n9193 GND.n9192 0.036
R7258 GND.n9191 GND.n9190 0.036
R7259 GND.n83 GND.n82 0.036
R7260 GND.n81 GND.n80 0.036
R7261 GND.n154 GND.n153 0.036
R7262 GND.n152 GND.n151 0.036
R7263 GND.n1698 GND.n1696 0.034
R7264 GND.n1678 GND.n1676 0.034
R7265 GND.n1370 GND.n1368 0.034
R7266 GND.n1390 GND.n1388 0.034
R7267 GND.n1193 GND.n1191 0.034
R7268 GND.n1173 GND.n1171 0.034
R7269 GND.n736 GND.n734 0.034
R7270 GND.n756 GND.n754 0.034
R7271 GND.n2798 GND.n2796 0.034
R7272 GND.n2818 GND.n2816 0.034
R7273 GND.n3121 GND.n3119 0.034
R7274 GND.n3101 GND.n3099 0.034
R7275 GND.n3711 GND.n3709 0.034
R7276 GND.n3691 GND.n3689 0.034
R7277 GND.n1914 GND.n1912 0.034
R7278 GND.n1934 GND.n1932 0.034
R7279 GND.n2094 GND.n2092 0.034
R7280 GND.n2114 GND.n2112 0.034
R7281 GND.n5224 GND.n5222 0.034
R7282 GND.n5244 GND.n5242 0.034
R7283 GND.n5404 GND.n5402 0.034
R7284 GND.n5424 GND.n5422 0.034
R7285 GND.n4474 GND.n4472 0.034
R7286 GND.n4494 GND.n4492 0.034
R7287 GND.n4656 GND.n4654 0.034
R7288 GND.n4677 GND.n4675 0.034
R7289 GND.n4845 GND.n4843 0.034
R7290 GND.n4865 GND.n4863 0.034
R7291 GND.n5025 GND.n5023 0.034
R7292 GND.n5045 GND.n5043 0.034
R7293 GND.n3502 GND.n3500 0.034
R7294 GND.n3481 GND.n3479 0.034
R7295 GND.n3318 GND.n3316 0.034
R7296 GND.n3298 GND.n3296 0.034
R7297 GND.n5900 GND.n5895 0.034
R7298 GND.n5800 GND.n5798 0.034
R7299 GND.n5780 GND.n5778 0.034
R7300 GND.n5620 GND.n5618 0.034
R7301 GND.n5600 GND.n5598 0.034
R7302 GND.n4203 GND.n4201 0.034
R7303 GND.n4223 GND.n4221 0.034
R7304 GND.n617 GND.n614 0.033
R7305 GND.n983 GND.n981 0.033
R7306 GND.n910 GND.n907 0.033
R7307 GND.n6087 GND.n6084 0.033
R7308 GND.n2605 GND.n2603 0.033
R7309 GND.n2532 GND.n2529 0.033
R7310 GND.n3915 GND.n3912 0.033
R7311 GND.n2383 GND.n2380 0.033
R7312 GND.n2976 GND.n2973 0.033
R7313 GND.n4087 GND.n4084 0.033
R7314 GND.n1555 GND.n1552 0.033
R7315 GND.n6204 GND.n6202 0.033
R7316 GND.n8281 GND.n8280 0.033
R7317 GND.n8208 GND.n8207 0.033
R7318 GND.n8388 GND.n8387 0.033
R7319 GND.n8459 GND.n8458 0.033
R7320 GND.n8573 GND.n8572 0.033
R7321 GND.n8644 GND.n8643 0.033
R7322 GND.n8758 GND.n8757 0.033
R7323 GND.n8829 GND.n8828 0.033
R7324 GND.n8943 GND.n8942 0.033
R7325 GND.n9014 GND.n9013 0.033
R7326 GND.n9128 GND.n9127 0.033
R7327 GND.n9199 GND.n9198 0.033
R7328 GND.n89 GND.n88 0.033
R7329 GND.n160 GND.n159 0.033
R7330 GND.n5974 GND.n5969 0.032
R7331 GND GND.n4376 0.032
R7332 GND.n3793 GND.n3790 0.032
R7333 GND.n7845 GND.n7843 0.031
R7334 GND.n7853 GND.n7852 0.031
R7335 GND.n7852 GND.n7851 0.031
R7336 GND.n7883 GND.n7881 0.031
R7337 GND.n8003 GND.n7996 0.031
R7338 GND.n8029 GND.n8021 0.031
R7339 GND.n8024 GND.n8023 0.031
R7340 GND.n8023 GND.n8022 0.031
R7341 GND.n7875 GND.n7870 0.031
R7342 GND.n7618 GND.n7616 0.031
R7343 GND.n7626 GND.n7625 0.031
R7344 GND.n7625 GND.n7624 0.031
R7345 GND.n7656 GND.n7654 0.031
R7346 GND.n7776 GND.n7769 0.031
R7347 GND.n7802 GND.n7794 0.031
R7348 GND.n7797 GND.n7796 0.031
R7349 GND.n7796 GND.n7795 0.031
R7350 GND.n7648 GND.n7643 0.031
R7351 GND.n7391 GND.n7389 0.031
R7352 GND.n7399 GND.n7398 0.031
R7353 GND.n7398 GND.n7397 0.031
R7354 GND.n7429 GND.n7427 0.031
R7355 GND.n7549 GND.n7542 0.031
R7356 GND.n7575 GND.n7567 0.031
R7357 GND.n7570 GND.n7569 0.031
R7358 GND.n7569 GND.n7568 0.031
R7359 GND.n7421 GND.n7416 0.031
R7360 GND.n7164 GND.n7162 0.031
R7361 GND.n7172 GND.n7171 0.031
R7362 GND.n7171 GND.n7170 0.031
R7363 GND.n7202 GND.n7200 0.031
R7364 GND.n7322 GND.n7315 0.031
R7365 GND.n7348 GND.n7340 0.031
R7366 GND.n7343 GND.n7342 0.031
R7367 GND.n7342 GND.n7341 0.031
R7368 GND.n7194 GND.n7189 0.031
R7369 GND.n6937 GND.n6935 0.031
R7370 GND.n6945 GND.n6944 0.031
R7371 GND.n6944 GND.n6943 0.031
R7372 GND.n6975 GND.n6973 0.031
R7373 GND.n7095 GND.n7088 0.031
R7374 GND.n7121 GND.n7113 0.031
R7375 GND.n7116 GND.n7115 0.031
R7376 GND.n7115 GND.n7114 0.031
R7377 GND.n6967 GND.n6962 0.031
R7378 GND.n6710 GND.n6708 0.031
R7379 GND.n6718 GND.n6717 0.031
R7380 GND.n6717 GND.n6716 0.031
R7381 GND.n6748 GND.n6746 0.031
R7382 GND.n6868 GND.n6861 0.031
R7383 GND.n6894 GND.n6886 0.031
R7384 GND.n6889 GND.n6888 0.031
R7385 GND.n6888 GND.n6887 0.031
R7386 GND.n6740 GND.n6735 0.031
R7387 GND.n6378 GND.n6376 0.031
R7388 GND.n6386 GND.n6385 0.031
R7389 GND.n6385 GND.n6384 0.031
R7390 GND.n6428 GND.n6426 0.031
R7391 GND.n6536 GND.n6529 0.031
R7392 GND.n6562 GND.n6554 0.031
R7393 GND.n6557 GND.n6556 0.031
R7394 GND.n6556 GND.n6555 0.031
R7395 GND.n6420 GND.n6415 0.031
R7396 GND.n545 GND.n543 0.031
R7397 GND.n556 GND.n554 0.031
R7398 GND.n649 GND.n647 0.031
R7399 GND.n950 GND.n948 0.031
R7400 GND.n1041 GND.n1039 0.031
R7401 GND.n1052 GND.n1050 0.031
R7402 GND.n860 GND.n858 0.031
R7403 GND.n871 GND.n869 0.031
R7404 GND.n942 GND.n940 0.031
R7405 GND.n6014 GND.n6012 0.031
R7406 GND.n6025 GND.n6023 0.031
R7407 GND.n6119 GND.n6117 0.031
R7408 GND.n2572 GND.n2570 0.031
R7409 GND.n2663 GND.n2661 0.031
R7410 GND.n2674 GND.n2672 0.031
R7411 GND.n2482 GND.n2480 0.031
R7412 GND.n2493 GND.n2491 0.031
R7413 GND.n2564 GND.n2562 0.031
R7414 GND.n3842 GND.n3840 0.031
R7415 GND.n3853 GND.n3851 0.031
R7416 GND.n3947 GND.n3945 0.031
R7417 GND.n3803 GND.n3199 0.031
R7418 GND.n2311 GND.n2309 0.031
R7419 GND.n2322 GND.n2320 0.031
R7420 GND.n2415 GND.n2413 0.031
R7421 GND.n3008 GND.n3006 0.031
R7422 GND.n2943 GND.n2941 0.031
R7423 GND.n2932 GND.n2930 0.031
R7424 GND.n4119 GND.n4117 0.031
R7425 GND.n4054 GND.n4052 0.031
R7426 GND.n4043 GND.n4041 0.031
R7427 GND.n1587 GND.n1585 0.031
R7428 GND.n1517 GND.n1515 0.031
R7429 GND.n1506 GND.n1504 0.031
R7430 GND.n6171 GND.n6169 0.031
R7431 GND.n6242 GND.n6240 0.031
R7432 GND.n6253 GND.n6251 0.031
R7433 GND.n8255 GND.n8253 0.031
R7434 GND.n8258 GND.n8257 0.031
R7435 GND.n8288 GND.n8287 0.031
R7436 GND.n8183 GND.n8181 0.031
R7437 GND.n8186 GND.n8185 0.031
R7438 GND.n8216 GND.n8214 0.031
R7439 GND.n8362 GND.n8360 0.031
R7440 GND.n8365 GND.n8364 0.031
R7441 GND.n8395 GND.n8394 0.031
R7442 GND.n8434 GND.n8432 0.031
R7443 GND.n8437 GND.n8436 0.031
R7444 GND.n8467 GND.n8465 0.031
R7445 GND.n8547 GND.n8545 0.031
R7446 GND.n8550 GND.n8549 0.031
R7447 GND.n8580 GND.n8579 0.031
R7448 GND.n8619 GND.n8617 0.031
R7449 GND.n8622 GND.n8621 0.031
R7450 GND.n8652 GND.n8650 0.031
R7451 GND.n8732 GND.n8730 0.031
R7452 GND.n8735 GND.n8734 0.031
R7453 GND.n8765 GND.n8764 0.031
R7454 GND.n8804 GND.n8802 0.031
R7455 GND.n8807 GND.n8806 0.031
R7456 GND.n8837 GND.n8835 0.031
R7457 GND.n8917 GND.n8915 0.031
R7458 GND.n8920 GND.n8919 0.031
R7459 GND.n8950 GND.n8949 0.031
R7460 GND.n8989 GND.n8987 0.031
R7461 GND.n8992 GND.n8991 0.031
R7462 GND.n9022 GND.n9020 0.031
R7463 GND.n9102 GND.n9100 0.031
R7464 GND.n9105 GND.n9104 0.031
R7465 GND.n9135 GND.n9134 0.031
R7466 GND.n9174 GND.n9172 0.031
R7467 GND.n9177 GND.n9176 0.031
R7468 GND.n9207 GND.n9205 0.031
R7469 GND.n63 GND.n61 0.031
R7470 GND.n66 GND.n65 0.031
R7471 GND.n96 GND.n95 0.031
R7472 GND.n135 GND.n133 0.031
R7473 GND.n138 GND.n137 0.031
R7474 GND.n168 GND.n166 0.031
R7475 GND.n1710 GND.n1708 0.03
R7476 GND.n1666 GND.n1664 0.03
R7477 GND.n1358 GND.n1356 0.03
R7478 GND.n1402 GND.n1400 0.03
R7479 GND.n1205 GND.n1203 0.03
R7480 GND.n1161 GND.n1159 0.03
R7481 GND.n724 GND.n722 0.03
R7482 GND.n768 GND.n766 0.03
R7483 GND.n2786 GND.n2784 0.03
R7484 GND.n2830 GND.n2828 0.03
R7485 GND.n3133 GND.n3131 0.03
R7486 GND.n3089 GND.n3087 0.03
R7487 GND.n3723 GND.n3721 0.03
R7488 GND.n3679 GND.n3677 0.03
R7489 GND.n1902 GND.n1900 0.03
R7490 GND.n1946 GND.n1944 0.03
R7491 GND.n2082 GND.n2080 0.03
R7492 GND.n2126 GND.n2124 0.03
R7493 GND.n5212 GND.n5210 0.03
R7494 GND.n5256 GND.n5254 0.03
R7495 GND.n5392 GND.n5390 0.03
R7496 GND.n5436 GND.n5434 0.03
R7497 GND.n4462 GND.n4460 0.03
R7498 GND.n4506 GND.n4504 0.03
R7499 GND.n4643 GND.n4641 0.03
R7500 GND.n4690 GND.n4688 0.03
R7501 GND.n4833 GND.n4831 0.03
R7502 GND.n4877 GND.n4875 0.03
R7503 GND.n5013 GND.n5011 0.03
R7504 GND.n5057 GND.n5055 0.03
R7505 GND.n3515 GND.n3513 0.03
R7506 GND.n3468 GND.n3466 0.03
R7507 GND.n3330 GND.n3328 0.03
R7508 GND.n3286 GND.n3284 0.03
R7509 GND.n5812 GND.n5810 0.03
R7510 GND.n5768 GND.n5766 0.03
R7511 GND.n5632 GND.n5630 0.03
R7512 GND.n5588 GND.n5586 0.03
R7513 GND.n4191 GND.n4189 0.03
R7514 GND.n4235 GND.n4233 0.03
R7515 GND.n7851 GND.n7850 0.028
R7516 GND.n7624 GND.n7623 0.028
R7517 GND.n7397 GND.n7396 0.028
R7518 GND.n7170 GND.n7169 0.028
R7519 GND.n6943 GND.n6942 0.028
R7520 GND.n6716 GND.n6715 0.028
R7521 GND.n6384 GND.n6383 0.028
R7522 GND.n624 GND.n621 0.028
R7523 GND.n1768 GND.n1766 0.028
R7524 GND.n1614 GND.n1605 0.028
R7525 GND.n1306 GND.n1297 0.028
R7526 GND.n1461 GND.n1459 0.028
R7527 GND.n1255 GND.n1254 0.028
R7528 GND.n1109 GND.n1101 0.028
R7529 GND.n6158 GND.n6156 0.028
R7530 GND.n818 GND.n817 0.028
R7531 GND.n2734 GND.n2725 0.028
R7532 GND.n2888 GND.n2886 0.028
R7533 GND.n3191 GND.n3189 0.028
R7534 GND.n3037 GND.n3028 0.028
R7535 GND.n3773 GND.n3772 0.028
R7536 GND.n3627 GND.n3619 0.028
R7537 GND.n976 GND.n974 0.028
R7538 GND.n917 GND.n914 0.028
R7539 GND.n6094 GND.n6091 0.028
R7540 GND.n2598 GND.n2596 0.028
R7541 GND.n2539 GND.n2536 0.028
R7542 GND.n3922 GND.n3919 0.028
R7543 GND.n3796 GND.n3793 0.028
R7544 GND.n1850 GND.n1849 0.028
R7545 GND.n2004 GND.n2002 0.028
R7546 GND.n2030 GND.n2022 0.028
R7547 GND.n2176 GND.n2175 0.028
R7548 GND.n5160 GND.n5159 0.028
R7549 GND.n5314 GND.n5312 0.028
R7550 GND.n5340 GND.n5332 0.028
R7551 GND.n5486 GND.n5485 0.028
R7552 GND.n4410 GND.n4409 0.028
R7553 GND.n4564 GND.n4562 0.028
R7554 GND.n4590 GND.n4582 0.028
R7555 GND.n4742 GND.n4741 0.028
R7556 GND.n4781 GND.n4780 0.028
R7557 GND.n4935 GND.n4933 0.028
R7558 GND.n4961 GND.n4953 0.028
R7559 GND.n5107 GND.n5106 0.028
R7560 GND.n3567 GND.n3566 0.028
R7561 GND.n3414 GND.n3406 0.028
R7562 GND.n3388 GND.n3386 0.028
R7563 GND.n3233 GND.n3232 0.028
R7564 GND.n5862 GND.n5861 0.028
R7565 GND.n5716 GND.n5708 0.028
R7566 GND.n5690 GND.n5688 0.028
R7567 GND.n5535 GND.n5534 0.028
R7568 GND.n2390 GND.n2387 0.028
R7569 GND.n2983 GND.n2980 0.028
R7570 GND.n4094 GND.n4091 0.028
R7571 GND.n4139 GND.n4130 0.028
R7572 GND.n4293 GND.n4291 0.028
R7573 GND.n1562 GND.n1559 0.028
R7574 GND.n6197 GND.n6195 0.028
R7575 GND.n8259 GND.n8258 0.028
R7576 GND.n8282 GND.n8281 0.028
R7577 GND.n8187 GND.n8186 0.028
R7578 GND.n8209 GND.n8208 0.028
R7579 GND.n8366 GND.n8365 0.028
R7580 GND.n8389 GND.n8388 0.028
R7581 GND.n8438 GND.n8437 0.028
R7582 GND.n8460 GND.n8459 0.028
R7583 GND.n8551 GND.n8550 0.028
R7584 GND.n8574 GND.n8573 0.028
R7585 GND.n8623 GND.n8622 0.028
R7586 GND.n8645 GND.n8644 0.028
R7587 GND.n8736 GND.n8735 0.028
R7588 GND.n8759 GND.n8758 0.028
R7589 GND.n8808 GND.n8807 0.028
R7590 GND.n8830 GND.n8829 0.028
R7591 GND.n8921 GND.n8920 0.028
R7592 GND.n8944 GND.n8943 0.028
R7593 GND.n8993 GND.n8992 0.028
R7594 GND.n9015 GND.n9014 0.028
R7595 GND.n9106 GND.n9105 0.028
R7596 GND.n9129 GND.n9128 0.028
R7597 GND.n9178 GND.n9177 0.028
R7598 GND.n9200 GND.n9199 0.028
R7599 GND.n67 GND.n66 0.028
R7600 GND.n90 GND.n89 0.028
R7601 GND.n139 GND.n138 0.028
R7602 GND.n161 GND.n160 0.028
R7603 GND.n8074 GND.n8072 0.028
R7604 GND.n1261 GND.n1260 0.027
R7605 GND.n7911 GND.n7909 0.026
R7606 GND.n7917 GND.n7916 0.026
R7607 GND.n7863 GND.n7861 0.026
R7608 GND.n7929 GND.n7922 0.026
R7609 GND.n7925 GND.n7924 0.026
R7610 GND.n7900 GND.n7897 0.026
R7611 GND.n7684 GND.n7682 0.026
R7612 GND.n7690 GND.n7689 0.026
R7613 GND.n7636 GND.n7634 0.026
R7614 GND.n7702 GND.n7695 0.026
R7615 GND.n7698 GND.n7697 0.026
R7616 GND.n7673 GND.n7670 0.026
R7617 GND.n7457 GND.n7455 0.026
R7618 GND.n7463 GND.n7462 0.026
R7619 GND.n7409 GND.n7407 0.026
R7620 GND.n7475 GND.n7468 0.026
R7621 GND.n7471 GND.n7470 0.026
R7622 GND.n7446 GND.n7443 0.026
R7623 GND.n7230 GND.n7228 0.026
R7624 GND.n7236 GND.n7235 0.026
R7625 GND.n7182 GND.n7180 0.026
R7626 GND.n7248 GND.n7241 0.026
R7627 GND.n7244 GND.n7243 0.026
R7628 GND.n7219 GND.n7216 0.026
R7629 GND.n7003 GND.n7001 0.026
R7630 GND.n7009 GND.n7008 0.026
R7631 GND.n6955 GND.n6953 0.026
R7632 GND.n7021 GND.n7014 0.026
R7633 GND.n7017 GND.n7016 0.026
R7634 GND.n6992 GND.n6989 0.026
R7635 GND.n6776 GND.n6774 0.026
R7636 GND.n6782 GND.n6781 0.026
R7637 GND.n6728 GND.n6726 0.026
R7638 GND.n6794 GND.n6787 0.026
R7639 GND.n6790 GND.n6789 0.026
R7640 GND.n6765 GND.n6762 0.026
R7641 GND.n6455 GND.n6453 0.026
R7642 GND.n6461 GND.n6460 0.026
R7643 GND.n6444 GND.n6442 0.026
R7644 GND.n6397 GND.n6390 0.026
R7645 GND.n6393 GND.n6392 0.026
R7646 GND.n6407 GND.n6404 0.026
R7647 GND.n590 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/DRAIN 0.026
R7648 GND.n524 GND.n522 0.026
R7649 GND.n534 GND.n532 0.026
R7650 GND.n538 GND.n537 0.026
R7651 GND.n541 GND.n538 0.026
R7652 GND.n642 GND.n640 0.026
R7653 GND.n957 GND.n955 0.026
R7654 GND.n1056 GND.n1055 0.026
R7655 GND.n1057 GND.n1056 0.026
R7656 GND.n1063 GND.n1061 0.026
R7657 GND.n1073 GND.n1071 0.026
R7658 GND.n6060 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/SOURCE 0.026
R7659 GND.n839 GND.n837 0.026
R7660 GND.n849 GND.n847 0.026
R7661 GND.n853 GND.n852 0.026
R7662 GND.n856 GND.n853 0.026
R7663 GND.n935 GND.n933 0.026
R7664 GND.n6124 GND.n6122 0.026
R7665 GND.n6138 GND.n6137 0.026
R7666 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/GATE GND.n6139 0.026
R7667 GND.n5993 GND.n5991 0.026
R7668 GND.n6003 GND.n6001 0.026
R7669 GND.n6007 GND.n6006 0.026
R7670 GND.n6010 GND.n6007 0.026
R7671 GND.n6112 GND.n6110 0.026
R7672 GND.n2579 GND.n2577 0.026
R7673 GND.n2678 GND.n2677 0.026
R7674 GND.n2679 GND.n2678 0.026
R7675 GND.n2685 GND.n2683 0.026
R7676 GND.n2695 GND.n2693 0.026
R7677 GND.n3888 GND 0.026
R7678 GND.n2461 GND.n2459 0.026
R7679 GND.n2471 GND.n2469 0.026
R7680 GND.n2475 GND.n2474 0.026
R7681 GND.n2478 GND.n2475 0.026
R7682 GND.n2557 GND.n2555 0.026
R7683 GND.n3952 GND.n3950 0.026
R7684 GND.n3966 GND.n3965 0.026
R7685 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/GATE GND.n3967 0.026
R7686 GND.n3821 GND.n3819 0.026
R7687 GND.n3831 GND.n3829 0.026
R7688 GND.n3835 GND.n3834 0.026
R7689 GND.n3838 GND.n3835 0.026
R7690 GND.n3940 GND.n3938 0.026
R7691 GND.n2356 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/DRAIN 0.026
R7692 GND.n2290 GND.n2288 0.026
R7693 GND.n2300 GND.n2298 0.026
R7694 GND.n2304 GND.n2303 0.026
R7695 GND.n2307 GND.n2304 0.026
R7696 GND.n2408 GND.n2406 0.026
R7697 GND.n3001 GND.n2999 0.026
R7698 GND.n2929 GND.n2926 0.026
R7699 GND.n2926 GND.n2925 0.026
R7700 GND.n2922 GND.n2920 0.026
R7701 GND.n2913 GND.n2911 0.026
R7702 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/GATE GND.n4123 0.026
R7703 GND.n4112 GND.n4110 0.026
R7704 GND.n4040 GND.n4037 0.026
R7705 GND.n4037 GND.n4036 0.026
R7706 GND.n4033 GND.n4031 0.026
R7707 GND.n4024 GND.n4022 0.026
R7708 GND.n1580 GND.n1578 0.026
R7709 GND.n1502 GND.n1499 0.026
R7710 GND.n1499 GND.n1498 0.026
R7711 GND.n1495 GND.n1493 0.026
R7712 GND.n1486 GND.n1484 0.026
R7713 GND.n6164 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/GATE 0.026
R7714 GND.n6178 GND.n6176 0.026
R7715 GND.n6257 GND.n6256 0.026
R7716 GND.n6258 GND.n6257 0.026
R7717 GND.n6264 GND.n6262 0.026
R7718 GND.n6274 GND.n6272 0.026
R7719 GND.n8233 GND.n8231 0.026
R7720 GND.n8244 GND.n8242 0.026
R7721 GND.n8283 GND.n8282 0.026
R7722 GND.n8274 GND.n8273 0.026
R7723 GND.n8161 GND.n8159 0.026
R7724 GND.n8172 GND.n8170 0.026
R7725 GND.n8210 GND.n8209 0.026
R7726 GND.n8200 GND.n8199 0.026
R7727 GND.n8340 GND.n8338 0.026
R7728 GND.n8351 GND.n8349 0.026
R7729 GND.n8390 GND.n8389 0.026
R7730 GND.n8381 GND.n8380 0.026
R7731 GND.n8412 GND.n8410 0.026
R7732 GND.n8423 GND.n8421 0.026
R7733 GND.n8461 GND.n8460 0.026
R7734 GND.n8452 GND.n8451 0.026
R7735 GND.n8525 GND.n8523 0.026
R7736 GND.n8536 GND.n8534 0.026
R7737 GND.n8575 GND.n8574 0.026
R7738 GND.n8566 GND.n8565 0.026
R7739 GND.n8597 GND.n8595 0.026
R7740 GND.n8608 GND.n8606 0.026
R7741 GND.n8646 GND.n8645 0.026
R7742 GND.n8637 GND.n8636 0.026
R7743 GND.n8710 GND.n8708 0.026
R7744 GND.n8721 GND.n8719 0.026
R7745 GND.n8760 GND.n8759 0.026
R7746 GND.n8751 GND.n8750 0.026
R7747 GND.n8782 GND.n8780 0.026
R7748 GND.n8793 GND.n8791 0.026
R7749 GND.n8831 GND.n8830 0.026
R7750 GND.n8822 GND.n8821 0.026
R7751 GND.n8895 GND.n8893 0.026
R7752 GND.n8906 GND.n8904 0.026
R7753 GND.n8945 GND.n8944 0.026
R7754 GND.n8936 GND.n8935 0.026
R7755 GND.n8967 GND.n8965 0.026
R7756 GND.n8978 GND.n8976 0.026
R7757 GND.n9016 GND.n9015 0.026
R7758 GND.n9007 GND.n9006 0.026
R7759 GND.n9080 GND.n9078 0.026
R7760 GND.n9091 GND.n9089 0.026
R7761 GND.n9130 GND.n9129 0.026
R7762 GND.n9121 GND.n9120 0.026
R7763 GND.n9152 GND.n9150 0.026
R7764 GND.n9163 GND.n9161 0.026
R7765 GND.n9201 GND.n9200 0.026
R7766 GND.n9192 GND.n9191 0.026
R7767 GND.n41 GND.n39 0.026
R7768 GND.n52 GND.n50 0.026
R7769 GND.n91 GND.n90 0.026
R7770 GND.n82 GND.n81 0.026
R7771 GND.n113 GND.n111 0.026
R7772 GND.n124 GND.n122 0.026
R7773 GND.n162 GND.n161 0.026
R7774 GND.n153 GND.n152 0.026
R7775 GND.n1722 GND.n1720 0.025
R7776 GND.n1654 GND.n1652 0.025
R7777 GND.n1346 GND.n1344 0.025
R7778 GND.n1414 GND.n1412 0.025
R7779 GND.n1217 GND.n1215 0.025
R7780 GND.n1149 GND.n1147 0.025
R7781 GND.n712 GND.n710 0.025
R7782 GND.n780 GND.n778 0.025
R7783 GND.n2774 GND.n2772 0.025
R7784 GND.n2842 GND.n2840 0.025
R7785 GND.n3145 GND.n3143 0.025
R7786 GND.n3077 GND.n3075 0.025
R7787 GND.n3735 GND.n3733 0.025
R7788 GND.n3667 GND.n3665 0.025
R7789 GND.n1890 GND.n1888 0.025
R7790 GND.n1958 GND.n1956 0.025
R7791 GND.n2070 GND.n2068 0.025
R7792 GND.n2138 GND.n2136 0.025
R7793 GND.n5200 GND.n5198 0.025
R7794 GND.n5268 GND.n5266 0.025
R7795 GND.n5380 GND.n5378 0.025
R7796 GND.n5448 GND.n5446 0.025
R7797 GND.n4450 GND.n4448 0.025
R7798 GND.n4518 GND.n4516 0.025
R7799 GND.n4631 GND.n4629 0.025
R7800 GND.n4702 GND.n4700 0.025
R7801 GND.n4821 GND.n4819 0.025
R7802 GND.n4889 GND.n4887 0.025
R7803 GND.n5001 GND.n4999 0.025
R7804 GND.n5069 GND.n5067 0.025
R7805 GND.n3527 GND.n3525 0.025
R7806 GND.n3456 GND.n3454 0.025
R7807 GND.n3342 GND.n3340 0.025
R7808 GND.n3274 GND.n3272 0.025
R7809 GND.n5824 GND.n5822 0.025
R7810 GND.n5756 GND.n5754 0.025
R7811 GND.n5644 GND.n5642 0.025
R7812 GND.n5576 GND.n5574 0.025
R7813 GND.n4179 GND.n4177 0.025
R7814 GND.n4247 GND.n4245 0.025
R7815 GND.n514 GND.n512 0.024
R7816 GND.n515 GND.n514 0.024
R7817 GND.n631 GND.n628 0.024
R7818 GND.n969 GND.n967 0.024
R7819 GND.n1081 GND.n1079 0.024
R7820 GND.n1082 GND.n1081 0.024
R7821 GND.n829 GND.n827 0.024
R7822 GND.n830 GND.n829 0.024
R7823 GND.n924 GND.n921 0.024
R7824 GND.n5983 GND.n5981 0.024
R7825 GND.n5984 GND.n5983 0.024
R7826 GND.n6101 GND.n6098 0.024
R7827 GND.n2591 GND.n2589 0.024
R7828 GND.n2703 GND.n2701 0.024
R7829 GND.n2704 GND.n2703 0.024
R7830 GND.n2451 GND.n2449 0.024
R7831 GND.n2452 GND.n2451 0.024
R7832 GND.n2546 GND.n2543 0.024
R7833 GND.n3811 GND.n3809 0.024
R7834 GND.n3812 GND.n3811 0.024
R7835 GND.n3929 GND.n3926 0.024
R7836 GND.n2280 GND.n2278 0.024
R7837 GND.n2281 GND.n2280 0.024
R7838 GND.n2397 GND.n2394 0.024
R7839 GND.n2990 GND.n2987 0.024
R7840 GND.n2905 GND.n2904 0.024
R7841 GND.n2904 GND.n2902 0.024
R7842 GND.n4101 GND.n4098 0.024
R7843 GND.n4016 GND.n4015 0.024
R7844 GND.n4015 GND.n4013 0.024
R7845 GND.n1569 GND.n1566 0.024
R7846 GND.n1478 GND.n1477 0.024
R7847 GND.n1477 GND.n1475 0.024
R7848 GND.n6190 GND.n6188 0.024
R7849 GND.n6282 GND.n6280 0.024
R7850 GND.n6283 GND.n6282 0.024
R7851 GND.n8223 GND.n8221 0.024
R7852 GND.n8224 GND.n8223 0.024
R7853 GND.n8151 GND.n8149 0.024
R7854 GND.n8152 GND.n8151 0.024
R7855 GND.n8330 GND.n8328 0.024
R7856 GND.n8331 GND.n8330 0.024
R7857 GND.n8402 GND.n8400 0.024
R7858 GND.n8403 GND.n8402 0.024
R7859 GND.n8515 GND.n8513 0.024
R7860 GND.n8516 GND.n8515 0.024
R7861 GND.n8587 GND.n8585 0.024
R7862 GND.n8588 GND.n8587 0.024
R7863 GND.n8700 GND.n8698 0.024
R7864 GND.n8701 GND.n8700 0.024
R7865 GND.n8772 GND.n8770 0.024
R7866 GND.n8773 GND.n8772 0.024
R7867 GND.n8885 GND.n8883 0.024
R7868 GND.n8886 GND.n8885 0.024
R7869 GND.n8957 GND.n8955 0.024
R7870 GND.n8958 GND.n8957 0.024
R7871 GND.n9070 GND.n9068 0.024
R7872 GND.n9071 GND.n9070 0.024
R7873 GND.n9142 GND.n9140 0.024
R7874 GND.n9143 GND.n9142 0.024
R7875 GND.n31 GND.n29 0.024
R7876 GND.n32 GND.n31 0.024
R7877 GND.n103 GND.n101 0.024
R7878 GND.n104 GND.n103 0.024
R7879 GND.n3802 GND.n3799 0.024
R7880 GND.n581 GND.n580 0.023
R7881 GND.n584 GND.n583 0.023
R7882 GND.n1756 GND.n1754 0.023
R7883 GND.n1626 GND.n1618 0.023
R7884 GND.n1318 GND.n1310 0.023
R7885 GND.n1449 GND.n1447 0.023
R7886 GND.n1251 GND.n1249 0.023
R7887 GND.n1121 GND.n1113 0.023
R7888 GND.n684 GND.n676 0.023
R7889 GND.n814 GND.n812 0.023
R7890 GND.n2746 GND.n2738 0.023
R7891 GND.n2876 GND.n2874 0.023
R7892 GND.n3179 GND.n3177 0.023
R7893 GND.n3049 GND.n3041 0.023
R7894 GND.n3769 GND.n3767 0.023
R7895 GND.n3639 GND.n3631 0.023
R7896 GND.n1015 GND.n1014 0.023
R7897 GND.n1012 GND.n1011 0.023
R7898 GND.n6051 GND.n6050 0.023
R7899 GND.n6054 GND.n6053 0.023
R7900 GND.n2637 GND.n2636 0.023
R7901 GND.n2634 GND.n2633 0.023
R7902 GND.n3879 GND.n3878 0.023
R7903 GND.n3882 GND.n3881 0.023
R7904 GND.n1862 GND.n1854 0.023
R7905 GND.n1992 GND.n1990 0.023
R7906 GND.n2042 GND.n2034 0.023
R7907 GND.n2172 GND.n2170 0.023
R7908 GND.n5172 GND.n5164 0.023
R7909 GND.n5302 GND.n5300 0.023
R7910 GND.n5352 GND.n5344 0.023
R7911 GND.n5482 GND.n5480 0.023
R7912 GND.n4422 GND.n4414 0.023
R7913 GND.n4552 GND.n4550 0.023
R7914 GND.n4602 GND.n4594 0.023
R7915 GND.n4738 GND.n4736 0.023
R7916 GND.n4793 GND.n4785 0.023
R7917 GND.n4923 GND.n4921 0.023
R7918 GND.n4973 GND.n4965 0.023
R7919 GND.n5103 GND.n5101 0.023
R7920 GND.n3563 GND.n3561 0.023
R7921 GND.n3427 GND.n3418 0.023
R7922 GND.n3376 GND.n3374 0.023
R7923 GND.n3246 GND.n3237 0.023
R7924 GND.n5858 GND.n5856 0.023
R7925 GND.n5728 GND.n5720 0.023
R7926 GND.n5678 GND.n5676 0.023
R7927 GND.n5548 GND.n5539 0.023
R7928 GND.n2347 GND.n2346 0.023
R7929 GND.n2350 GND.n2349 0.023
R7930 GND.n3998 GND.n3997 0.023
R7931 GND.n4001 GND.n4000 0.023
R7932 GND.n4151 GND.n4143 0.023
R7933 GND.n4281 GND.n4279 0.023
R7934 GND.n6294 GND.n6293 0.023
R7935 GND.n6297 GND.n6296 0.023
R7936 GND.n1023 GND.n1021 0.022
R7937 GND.n2645 GND.n2643 0.022
R7938 GND.n7970 GND.n7966 0.021
R7939 GND.n8011 GND.n8010 0.021
R7940 GND.n7853 GND.n7848 0.021
R7941 GND.n7917 GND.n7914 0.021
R7942 GND.n7858 GND.n7856 0.021
R7943 GND.n7964 GND.n7959 0.021
R7944 GND.n8027 GND.n8024 0.021
R7945 GND.n7928 GND.n7925 0.021
R7946 GND.n7901 GND.n7894 0.021
R7947 GND.n7743 GND.n7739 0.021
R7948 GND.n7784 GND.n7783 0.021
R7949 GND.n7626 GND.n7621 0.021
R7950 GND.n7690 GND.n7687 0.021
R7951 GND.n7631 GND.n7629 0.021
R7952 GND.n7737 GND.n7732 0.021
R7953 GND.n7800 GND.n7797 0.021
R7954 GND.n7701 GND.n7698 0.021
R7955 GND.n7674 GND.n7667 0.021
R7956 GND.n7516 GND.n7512 0.021
R7957 GND.n7557 GND.n7556 0.021
R7958 GND.n7399 GND.n7394 0.021
R7959 GND.n7463 GND.n7460 0.021
R7960 GND.n7404 GND.n7402 0.021
R7961 GND.n7510 GND.n7505 0.021
R7962 GND.n7573 GND.n7570 0.021
R7963 GND.n7474 GND.n7471 0.021
R7964 GND.n7447 GND.n7440 0.021
R7965 GND.n7289 GND.n7285 0.021
R7966 GND.n7330 GND.n7329 0.021
R7967 GND.n7172 GND.n7167 0.021
R7968 GND.n7236 GND.n7233 0.021
R7969 GND.n7177 GND.n7175 0.021
R7970 GND.n7283 GND.n7278 0.021
R7971 GND.n7346 GND.n7343 0.021
R7972 GND.n7247 GND.n7244 0.021
R7973 GND.n7220 GND.n7213 0.021
R7974 GND.n7062 GND.n7058 0.021
R7975 GND.n7103 GND.n7102 0.021
R7976 GND.n6945 GND.n6940 0.021
R7977 GND.n7009 GND.n7006 0.021
R7978 GND.n6950 GND.n6948 0.021
R7979 GND.n7056 GND.n7051 0.021
R7980 GND.n7119 GND.n7116 0.021
R7981 GND.n7020 GND.n7017 0.021
R7982 GND.n6993 GND.n6986 0.021
R7983 GND.n6835 GND.n6831 0.021
R7984 GND.n6876 GND.n6875 0.021
R7985 GND.n6718 GND.n6713 0.021
R7986 GND.n6782 GND.n6779 0.021
R7987 GND.n6723 GND.n6721 0.021
R7988 GND.n6829 GND.n6824 0.021
R7989 GND.n6892 GND.n6889 0.021
R7990 GND.n6793 GND.n6790 0.021
R7991 GND.n6766 GND.n6759 0.021
R7992 GND.n6503 GND.n6499 0.021
R7993 GND.n6544 GND.n6543 0.021
R7994 GND.n6386 GND.n6381 0.021
R7995 GND.n6461 GND.n6458 0.021
R7996 GND.n6439 GND.n6437 0.021
R7997 GND.n6497 GND.n6492 0.021
R7998 GND.n6560 GND.n6557 0.021
R7999 GND.n6396 GND.n6393 0.021
R8000 GND.n6408 GND.n6401 0.021
R8001 GND.n567 GND.n566 0.021
R8002 GND.n635 GND.n633 0.021
R8003 GND.n1734 GND.n1732 0.021
R8004 GND.n1642 GND.n1640 0.021
R8005 GND.n1334 GND.n1332 0.021
R8006 GND.n1426 GND.n1424 0.021
R8007 GND.n1229 GND.n1227 0.021
R8008 GND.n1137 GND.n1135 0.021
R8009 GND.n700 GND.n698 0.021
R8010 GND.n792 GND.n790 0.021
R8011 GND.n2762 GND.n2760 0.021
R8012 GND.n2854 GND.n2852 0.021
R8013 GND.n3157 GND.n3155 0.021
R8014 GND.n3065 GND.n3063 0.021
R8015 GND.n3747 GND.n3745 0.021
R8016 GND.n3655 GND.n3653 0.021
R8017 GND.n964 GND.n962 0.021
R8018 GND.n1032 GND.n1026 0.021
R8019 GND.n882 GND.n881 0.021
R8020 GND.n928 GND.n926 0.021
R8021 GND.n6036 GND.n6035 0.021
R8022 GND.n6105 GND.n6103 0.021
R8023 GND.n2586 GND.n2584 0.021
R8024 GND.n2654 GND.n2648 0.021
R8025 GND.n2504 GND.n2503 0.021
R8026 GND.n2550 GND.n2548 0.021
R8027 GND.n3864 GND.n3863 0.021
R8028 GND.n3933 GND.n3931 0.021
R8029 GND.n1878 GND.n1876 0.021
R8030 GND.n1970 GND.n1968 0.021
R8031 GND.n2058 GND.n2056 0.021
R8032 GND.n2150 GND.n2148 0.021
R8033 GND.n5188 GND.n5186 0.021
R8034 GND.n5280 GND.n5278 0.021
R8035 GND.n5368 GND.n5366 0.021
R8036 GND.n5460 GND.n5458 0.021
R8037 GND.n4438 GND.n4436 0.021
R8038 GND.n4530 GND.n4528 0.021
R8039 GND.n4618 GND.n4616 0.021
R8040 GND.n4715 GND.n4713 0.021
R8041 GND.n4809 GND.n4807 0.021
R8042 GND.n4901 GND.n4899 0.021
R8043 GND.n4989 GND.n4987 0.021
R8044 GND.n5081 GND.n5079 0.021
R8045 GND.n3540 GND.n3538 0.021
R8046 GND.n3443 GND.n3441 0.021
R8047 GND.n3354 GND.n3352 0.021
R8048 GND.n3262 GND.n3260 0.021
R8049 GND.n5882 GND.n5877 0.021
R8050 GND.n5836 GND.n5834 0.021
R8051 GND.n5744 GND.n5742 0.021
R8052 GND.n5656 GND.n5654 0.021
R8053 GND.n5564 GND.n5562 0.021
R8054 GND.n5529 GND.n5528 0.021
R8055 GND.n4308 GND.n2252 0.021
R8056 GND.n2333 GND.n2332 0.021
R8057 GND.n2401 GND.n2399 0.021
R8058 GND.n2994 GND.n2992 0.021
R8059 GND.n2949 GND.n2948 0.021
R8060 GND.n4105 GND.n4103 0.021
R8061 GND.n4060 GND.n4059 0.021
R8062 GND.n4167 GND.n4165 0.021
R8063 GND.n4259 GND.n4257 0.021
R8064 GND.n1573 GND.n1571 0.021
R8065 GND.n1528 GND.n1527 0.021
R8066 GND.n6185 GND.n6183 0.021
R8067 GND.n6233 GND.n6228 0.021
R8068 GND.n8279 GND.n8278 0.021
R8069 GND.n8206 GND.n8205 0.021
R8070 GND.n8386 GND.n8385 0.021
R8071 GND.n8457 GND.n8456 0.021
R8072 GND.n8571 GND.n8570 0.021
R8073 GND.n8642 GND.n8641 0.021
R8074 GND.n8756 GND.n8755 0.021
R8075 GND.n8827 GND.n8826 0.021
R8076 GND.n8941 GND.n8940 0.021
R8077 GND.n9012 GND.n9011 0.021
R8078 GND.n9126 GND.n9125 0.021
R8079 GND.n9197 GND.n9196 0.021
R8080 GND.n87 GND.n86 0.021
R8081 GND.n158 GND.n157 0.021
R8082 GND.n2190 GND.n2182 0.02
R8083 GND.n5499 GND.n2190 0.02
R8084 GND.n5499 GND.n4397 0.02
R8085 GND.n4397 GND.n4389 0.02
R8086 GND.n7982 GND.n7981 0.019
R8087 GND.n7884 GND.n7883 0.019
R8088 GND.n7991 GND.n7990 0.019
R8089 GND.n7893 GND.n7891 0.019
R8090 GND.n7870 GND.n7868 0.019
R8091 GND.n7755 GND.n7754 0.019
R8092 GND.n7657 GND.n7656 0.019
R8093 GND.n7764 GND.n7763 0.019
R8094 GND.n7666 GND.n7664 0.019
R8095 GND.n7643 GND.n7641 0.019
R8096 GND.n7528 GND.n7527 0.019
R8097 GND.n7430 GND.n7429 0.019
R8098 GND.n7537 GND.n7536 0.019
R8099 GND.n7439 GND.n7437 0.019
R8100 GND.n7416 GND.n7414 0.019
R8101 GND.n7301 GND.n7300 0.019
R8102 GND.n7203 GND.n7202 0.019
R8103 GND.n7310 GND.n7309 0.019
R8104 GND.n7212 GND.n7210 0.019
R8105 GND.n7189 GND.n7187 0.019
R8106 GND.n7074 GND.n7073 0.019
R8107 GND.n6976 GND.n6975 0.019
R8108 GND.n7083 GND.n7082 0.019
R8109 GND.n6985 GND.n6983 0.019
R8110 GND.n6962 GND.n6960 0.019
R8111 GND.n6847 GND.n6846 0.019
R8112 GND.n6749 GND.n6748 0.019
R8113 GND.n6856 GND.n6855 0.019
R8114 GND.n6758 GND.n6756 0.019
R8115 GND.n6735 GND.n6733 0.019
R8116 GND.n6515 GND.n6514 0.019
R8117 GND.n6429 GND.n6428 0.019
R8118 GND.n6524 GND.n6523 0.019
R8119 GND.n6400 GND.n6398 0.019
R8120 GND.n6415 GND.n6413 0.019
R8121 GND.n525 GND.n524 0.019
R8122 GND.n560 GND.n558 0.019
R8123 GND.n569 GND.n567 0.019
R8124 GND.n595 GND.n594 0.019
R8125 GND.n638 GND.n635 0.019
R8126 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/SUBSTRATE GND.n1770 0.019
R8127 GND.n1744 GND.n1742 0.019
R8128 GND.n1638 GND.n1630 0.019
R8129 GND.n1330 GND.n1322 0.019
R8130 GND.n1436 GND.n1434 0.019
R8131 GND.n1256 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/SUBSTRATE 0.019
R8132 GND.n1239 GND.n1237 0.019
R8133 GND.n1133 GND.n1125 0.019
R8134 GND.n696 GND.n688 0.019
R8135 GND.n802 GND.n800 0.019
R8136 GND.n2758 GND.n2750 0.019
R8137 GND.n2864 GND.n2862 0.019
R8138 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/SUBSTRATE GND.n3193 0.019
R8139 GND.n3167 GND.n3165 0.019
R8140 GND.n3061 GND.n3053 0.019
R8141 GND.n3774 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/SUBSTRATE 0.019
R8142 GND.n3757 GND.n3755 0.019
R8143 GND.n3651 GND.n3643 0.019
R8144 GND.n962 GND.n960 0.019
R8145 GND.n1026 GND.n1025 0.019
R8146 GND.n1037 GND.n1035 0.019
R8147 GND.n1071 GND.n1069 0.019
R8148 GND.n840 GND.n839 0.019
R8149 GND.n875 GND.n873 0.019
R8150 GND.n884 GND.n882 0.019
R8151 GND.n888 GND.n887 0.019
R8152 GND.n931 GND.n928 0.019
R8153 GND.n5994 GND.n5993 0.019
R8154 GND.n6029 GND.n6027 0.019
R8155 GND.n6038 GND.n6036 0.019
R8156 GND.n6065 GND.n6064 0.019
R8157 GND.n6108 GND.n6105 0.019
R8158 GND.n2584 GND.n2582 0.019
R8159 GND.n2648 GND.n2647 0.019
R8160 GND.n2659 GND.n2657 0.019
R8161 GND.n2693 GND.n2691 0.019
R8162 GND.n2462 GND.n2461 0.019
R8163 GND.n2497 GND.n2495 0.019
R8164 GND.n2506 GND.n2504 0.019
R8165 GND.n2510 GND.n2509 0.019
R8166 GND.n2553 GND.n2550 0.019
R8167 GND.n3822 GND.n3821 0.019
R8168 GND.n3857 GND.n3855 0.019
R8169 GND.n3866 GND.n3864 0.019
R8170 GND.n3893 GND.n3892 0.019
R8171 GND.n3936 GND.n3933 0.019
R8172 GND.n1848 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/SUBSTRATE 0.019
R8173 GND.n1874 GND.n1866 0.019
R8174 GND.n1980 GND.n1978 0.019
R8175 GND.n2054 GND.n2046 0.019
R8176 GND.n2160 GND.n2158 0.019
R8177 GND.n5158 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/SUBSTRATE 0.019
R8178 GND.n5184 GND.n5176 0.019
R8179 GND.n5290 GND.n5288 0.019
R8180 GND.n5364 GND.n5356 0.019
R8181 GND.n5470 GND.n5468 0.019
R8182 GND.n4408 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SUBSTRATE 0.019
R8183 GND.n4434 GND.n4426 0.019
R8184 GND.n4540 GND.n4538 0.019
R8185 GND.n4614 GND.n4606 0.019
R8186 GND.n4725 GND.n4723 0.019
R8187 GND.n4779 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SUBSTRATE 0.019
R8188 GND.n4805 GND.n4797 0.019
R8189 GND.n4911 GND.n4909 0.019
R8190 GND.n4985 GND.n4977 0.019
R8191 GND.n5091 GND.n5089 0.019
R8192 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/SUBSTRATE GND.n3568 0.019
R8193 GND.n3550 GND.n3548 0.019
R8194 GND.n3439 GND.n3431 0.019
R8195 GND.n3364 GND.n3362 0.019
R8196 GND.n3258 GND.n3250 0.019
R8197 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/SUBSTRATE GND.n5863 0.019
R8198 GND.n5846 GND.n5844 0.019
R8199 GND.n5740 GND.n5732 0.019
R8200 GND.n5666 GND.n5664 0.019
R8201 GND.n5560 GND.n5552 0.019
R8202 GND.n2291 GND.n2290 0.019
R8203 GND.n2326 GND.n2324 0.019
R8204 GND.n2335 GND.n2333 0.019
R8205 GND.n2361 GND.n2360 0.019
R8206 GND.n2404 GND.n2401 0.019
R8207 GND.n2997 GND.n2994 0.019
R8208 GND.n2954 GND.n2953 0.019
R8209 GND.n2951 GND.n2949 0.019
R8210 GND.n2946 GND.n2945 0.019
R8211 GND.n2914 GND.n2913 0.019
R8212 GND.n4108 GND.n4105 0.019
R8213 GND.n4065 GND.n4064 0.019
R8214 GND.n4062 GND.n4060 0.019
R8215 GND.n4057 GND.n4056 0.019
R8216 GND.n4025 GND.n4024 0.019
R8217 GND.n4163 GND.n4155 0.019
R8218 GND.n4269 GND.n4267 0.019
R8219 GND.n1576 GND.n1573 0.019
R8220 GND.n1533 GND.n1532 0.019
R8221 GND.n1530 GND.n1528 0.019
R8222 GND.n1520 GND.n1519 0.019
R8223 GND.n1487 GND.n1486 0.019
R8224 GND.n6183 GND.n6181 0.019
R8225 GND.n6223 GND.n6222 0.019
R8226 GND.n6228 GND.n6227 0.019
R8227 GND.n6238 GND.n6236 0.019
R8228 GND.n6272 GND.n6270 0.019
R8229 GND.n8236 GND.n8235 0.019
R8230 GND.n8285 GND.n8283 0.019
R8231 GND.n8280 GND.n8279 0.019
R8232 GND.n8278 GND.n8277 0.019
R8233 GND.n8164 GND.n8163 0.019
R8234 GND.n8212 GND.n8210 0.019
R8235 GND.n8207 GND.n8206 0.019
R8236 GND.n8205 GND.n8204 0.019
R8237 GND.n8343 GND.n8342 0.019
R8238 GND.n8392 GND.n8390 0.019
R8239 GND.n8387 GND.n8386 0.019
R8240 GND.n8385 GND.n8384 0.019
R8241 GND.n8415 GND.n8414 0.019
R8242 GND.n8463 GND.n8461 0.019
R8243 GND.n8458 GND.n8457 0.019
R8244 GND.n8456 GND.n8455 0.019
R8245 GND.n8528 GND.n8527 0.019
R8246 GND.n8577 GND.n8575 0.019
R8247 GND.n8572 GND.n8571 0.019
R8248 GND.n8570 GND.n8569 0.019
R8249 GND.n8600 GND.n8599 0.019
R8250 GND.n8648 GND.n8646 0.019
R8251 GND.n8643 GND.n8642 0.019
R8252 GND.n8641 GND.n8640 0.019
R8253 GND.n8713 GND.n8712 0.019
R8254 GND.n8762 GND.n8760 0.019
R8255 GND.n8757 GND.n8756 0.019
R8256 GND.n8755 GND.n8754 0.019
R8257 GND.n8785 GND.n8784 0.019
R8258 GND.n8833 GND.n8831 0.019
R8259 GND.n8828 GND.n8827 0.019
R8260 GND.n8826 GND.n8825 0.019
R8261 GND.n8898 GND.n8897 0.019
R8262 GND.n8947 GND.n8945 0.019
R8263 GND.n8942 GND.n8941 0.019
R8264 GND.n8940 GND.n8939 0.019
R8265 GND.n8970 GND.n8969 0.019
R8266 GND.n9018 GND.n9016 0.019
R8267 GND.n9013 GND.n9012 0.019
R8268 GND.n9011 GND.n9010 0.019
R8269 GND.n9083 GND.n9082 0.019
R8270 GND.n9132 GND.n9130 0.019
R8271 GND.n9127 GND.n9126 0.019
R8272 GND.n9125 GND.n9124 0.019
R8273 GND.n9155 GND.n9154 0.019
R8274 GND.n9203 GND.n9201 0.019
R8275 GND.n9198 GND.n9197 0.019
R8276 GND.n9196 GND.n9195 0.019
R8277 GND.n44 GND.n43 0.019
R8278 GND.n93 GND.n91 0.019
R8279 GND.n88 GND.n87 0.019
R8280 GND.n86 GND.n85 0.019
R8281 GND.n116 GND.n115 0.019
R8282 GND.n164 GND.n162 0.019
R8283 GND.n159 GND.n158 0.019
R8284 GND.n157 GND.n156 0.019
R8285 GND.n2897 GND.n2896 0.018
R8286 GND.n4300 GND.n4298 0.018
R8287 GND.n4297 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/GATE 0.018
R8288 GND.n1470 GND.n1469 0.018
R8289 GND.n6314 GND.n6313 0.018
R8290 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/GATE GND.n6315 0.018
R8291 GND.n8125 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE 0.018
R8292 GND.n8476 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/SOURCE 0.018
R8293 GND.n8661 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/SOURCE 0.018
R8294 GND.n8846 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/SOURCE 0.018
R8295 GND.n9031 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/SOURCE 0.018
R8296 GND.n9216 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/SOURCE 0.018
R8297 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6/SOURCE GND.n9262 0.018
R8298 GND.n8234 GND.n8233 0.017
R8299 GND.n8162 GND.n8161 0.017
R8300 GND.n8341 GND.n8340 0.017
R8301 GND.n8413 GND.n8412 0.017
R8302 GND.n8526 GND.n8525 0.017
R8303 GND.n8598 GND.n8597 0.017
R8304 GND.n8711 GND.n8710 0.017
R8305 GND.n8783 GND.n8782 0.017
R8306 GND.n8896 GND.n8895 0.017
R8307 GND.n8968 GND.n8967 0.017
R8308 GND.n9081 GND.n9080 0.017
R8309 GND.n9153 GND.n9152 0.017
R8310 GND.n42 GND.n41 0.017
R8311 GND.n114 GND.n113 0.017
R8312 GND.n1746 GND.n1744 0.017
R8313 GND.n1630 GND.n1628 0.017
R8314 GND.n1322 GND.n1320 0.017
R8315 GND.n1438 GND.n1436 0.017
R8316 GND.n1241 GND.n1239 0.017
R8317 GND.n1125 GND.n1123 0.017
R8318 GND.n688 GND.n686 0.017
R8319 GND.n804 GND.n802 0.017
R8320 GND.n2750 GND.n2748 0.017
R8321 GND.n2866 GND.n2864 0.017
R8322 GND.n3169 GND.n3167 0.017
R8323 GND.n3053 GND.n3051 0.017
R8324 GND.n3759 GND.n3757 0.017
R8325 GND.n3643 GND.n3641 0.017
R8326 GND.n1866 GND.n1864 0.017
R8327 GND.n1982 GND.n1980 0.017
R8328 GND.n2046 GND.n2044 0.017
R8329 GND.n2162 GND.n2160 0.017
R8330 GND.n5176 GND.n5174 0.017
R8331 GND.n5292 GND.n5290 0.017
R8332 GND.n5356 GND.n5354 0.017
R8333 GND.n5472 GND.n5470 0.017
R8334 GND.n4426 GND.n4424 0.017
R8335 GND.n4542 GND.n4540 0.017
R8336 GND.n4606 GND.n4604 0.017
R8337 GND.n4727 GND.n4725 0.017
R8338 GND.n4797 GND.n4795 0.017
R8339 GND.n4913 GND.n4911 0.017
R8340 GND.n4977 GND.n4975 0.017
R8341 GND.n5093 GND.n5091 0.017
R8342 GND.n3552 GND.n3550 0.017
R8343 GND.n3431 GND.n3429 0.017
R8344 GND.n3366 GND.n3364 0.017
R8345 GND.n3250 GND.n3248 0.017
R8346 GND.n5848 GND.n5846 0.017
R8347 GND.n5732 GND.n5730 0.017
R8348 GND.n5668 GND.n5666 0.017
R8349 GND.n5552 GND.n5550 0.017
R8350 GND.n4155 GND.n4153 0.017
R8351 GND.n4271 GND.n4269 0.017
R8352 GND.n8074 GND.n6362 0.017
R8353 GND.n8012 GND.n8009 0.016
R8354 GND.n7863 GND.n7862 0.016
R8355 GND.n8002 GND.n7999 0.016
R8356 GND.n7897 GND.n7896 0.016
R8357 GND.n7785 GND.n7782 0.016
R8358 GND.n7636 GND.n7635 0.016
R8359 GND.n7775 GND.n7772 0.016
R8360 GND.n7670 GND.n7669 0.016
R8361 GND.n7558 GND.n7555 0.016
R8362 GND.n7409 GND.n7408 0.016
R8363 GND.n7548 GND.n7545 0.016
R8364 GND.n7443 GND.n7442 0.016
R8365 GND.n7331 GND.n7328 0.016
R8366 GND.n7182 GND.n7181 0.016
R8367 GND.n7321 GND.n7318 0.016
R8368 GND.n7216 GND.n7215 0.016
R8369 GND.n7104 GND.n7101 0.016
R8370 GND.n6955 GND.n6954 0.016
R8371 GND.n7094 GND.n7091 0.016
R8372 GND.n6989 GND.n6988 0.016
R8373 GND.n6877 GND.n6874 0.016
R8374 GND.n6728 GND.n6727 0.016
R8375 GND.n6867 GND.n6864 0.016
R8376 GND.n6762 GND.n6761 0.016
R8377 GND.n6545 GND.n6542 0.016
R8378 GND.n6444 GND.n6443 0.016
R8379 GND.n6535 GND.n6532 0.016
R8380 GND.n6404 GND.n6403 0.016
R8381 GND.n549 GND.n548 0.016
R8382 GND.n628 GND.n626 0.016
R8383 GND.n971 GND.n969 0.016
R8384 GND.n1046 GND.n1045 0.016
R8385 GND.n864 GND.n863 0.016
R8386 GND.n921 GND.n919 0.016
R8387 GND.n6018 GND.n6017 0.016
R8388 GND.n6098 GND.n6096 0.016
R8389 GND.n2593 GND.n2591 0.016
R8390 GND.n2668 GND.n2667 0.016
R8391 GND.n2486 GND.n2485 0.016
R8392 GND.n2543 GND.n2541 0.016
R8393 GND.n3846 GND.n3845 0.016
R8394 GND.n3926 GND.n3924 0.016
R8395 GND.n2315 GND.n2314 0.016
R8396 GND.n2394 GND.n2392 0.016
R8397 GND.n2987 GND.n2985 0.016
R8398 GND.n2936 GND.n2935 0.016
R8399 GND.n4098 GND.n4096 0.016
R8400 GND.n4047 GND.n4046 0.016
R8401 GND.n1566 GND.n1564 0.016
R8402 GND.n1510 GND.n1509 0.016
R8403 GND.n6192 GND.n6190 0.016
R8404 GND.n6247 GND.n6246 0.016
R8405 GND.n8260 GND.n8259 0.016
R8406 GND.n8188 GND.n8187 0.016
R8407 GND.n8367 GND.n8366 0.016
R8408 GND.n8439 GND.n8438 0.016
R8409 GND.n8552 GND.n8551 0.016
R8410 GND.n8624 GND.n8623 0.016
R8411 GND.n8737 GND.n8736 0.016
R8412 GND.n8809 GND.n8808 0.016
R8413 GND.n8922 GND.n8921 0.016
R8414 GND.n8994 GND.n8993 0.016
R8415 GND.n9107 GND.n9106 0.016
R8416 GND.n9179 GND.n9178 0.016
R8417 GND.n68 GND.n67 0.016
R8418 GND.n140 GND.n139 0.016
R8419 GND.n1732 GND.n1730 0.015
R8420 GND.n1650 GND.n1642 0.015
R8421 GND.n1342 GND.n1334 0.015
R8422 GND.n1424 GND.n1422 0.015
R8423 GND.n1227 GND.n1225 0.015
R8424 GND.n1145 GND.n1137 0.015
R8425 GND.n708 GND.n700 0.015
R8426 GND.n790 GND.n788 0.015
R8427 GND.n2770 GND.n2762 0.015
R8428 GND.n2852 GND.n2850 0.015
R8429 GND.n3155 GND.n3153 0.015
R8430 GND.n3073 GND.n3065 0.015
R8431 GND.n3745 GND.n3743 0.015
R8432 GND.n3663 GND.n3655 0.015
R8433 GND.n1886 GND.n1878 0.015
R8434 GND.n1968 GND.n1966 0.015
R8435 GND.n2066 GND.n2058 0.015
R8436 GND.n2148 GND.n2146 0.015
R8437 GND.n5492 GND.n5148 0.015
R8438 GND.n5196 GND.n5188 0.015
R8439 GND.n5278 GND.n5276 0.015
R8440 GND.n5376 GND.n5368 0.015
R8441 GND.n5458 GND.n5456 0.015
R8442 GND.n4446 GND.n4438 0.015
R8443 GND.n4528 GND.n4526 0.015
R8444 GND.n4627 GND.n4618 0.015
R8445 GND.n4713 GND.n4711 0.015
R8446 GND.n4817 GND.n4809 0.015
R8447 GND.n4899 GND.n4897 0.015
R8448 GND.n4997 GND.n4989 0.015
R8449 GND.n5079 GND.n5077 0.015
R8450 GND.n3538 GND.n3536 0.015
R8451 GND.n3452 GND.n3443 0.015
R8452 GND.n3352 GND.n3350 0.015
R8453 GND.n3270 GND.n3262 0.015
R8454 GND.n5834 GND.n5832 0.015
R8455 GND.n5752 GND.n5744 0.015
R8456 GND.n5654 GND.n5652 0.015
R8457 GND.n5572 GND.n5564 0.015
R8458 GND.n4175 GND.n4167 0.015
R8459 GND.n4257 GND.n4255 0.015
R8460 GND.n7940 GND.n7939 0.014
R8461 GND.n7945 GND.n7944 0.014
R8462 GND.n7944 GND.n7943 0.014
R8463 GND.n7914 GND.n7911 0.014
R8464 GND.n7861 GND.n7858 0.014
R8465 GND.n7950 GND.n7949 0.014
R8466 GND.n7955 GND.n7951 0.014
R8467 GND.n7955 GND.n7954 0.014
R8468 GND.n7922 GND.n7920 0.014
R8469 GND.n7929 GND.n7928 0.014
R8470 GND.n7901 GND.n7900 0.014
R8471 GND.n7713 GND.n7712 0.014
R8472 GND.n7718 GND.n7717 0.014
R8473 GND.n7717 GND.n7716 0.014
R8474 GND.n7687 GND.n7684 0.014
R8475 GND.n7634 GND.n7631 0.014
R8476 GND.n7723 GND.n7722 0.014
R8477 GND.n7728 GND.n7724 0.014
R8478 GND.n7728 GND.n7727 0.014
R8479 GND.n7695 GND.n7693 0.014
R8480 GND.n7702 GND.n7701 0.014
R8481 GND.n7674 GND.n7673 0.014
R8482 GND.n7486 GND.n7485 0.014
R8483 GND.n7491 GND.n7490 0.014
R8484 GND.n7490 GND.n7489 0.014
R8485 GND.n7460 GND.n7457 0.014
R8486 GND.n7407 GND.n7404 0.014
R8487 GND.n7496 GND.n7495 0.014
R8488 GND.n7501 GND.n7497 0.014
R8489 GND.n7501 GND.n7500 0.014
R8490 GND.n7468 GND.n7466 0.014
R8491 GND.n7475 GND.n7474 0.014
R8492 GND.n7447 GND.n7446 0.014
R8493 GND.n7259 GND.n7258 0.014
R8494 GND.n7264 GND.n7263 0.014
R8495 GND.n7263 GND.n7262 0.014
R8496 GND.n7233 GND.n7230 0.014
R8497 GND.n7180 GND.n7177 0.014
R8498 GND.n7269 GND.n7268 0.014
R8499 GND.n7274 GND.n7270 0.014
R8500 GND.n7274 GND.n7273 0.014
R8501 GND.n7241 GND.n7239 0.014
R8502 GND.n7248 GND.n7247 0.014
R8503 GND.n7220 GND.n7219 0.014
R8504 GND.n7032 GND.n7031 0.014
R8505 GND.n7037 GND.n7036 0.014
R8506 GND.n7036 GND.n7035 0.014
R8507 GND.n7006 GND.n7003 0.014
R8508 GND.n6953 GND.n6950 0.014
R8509 GND.n7042 GND.n7041 0.014
R8510 GND.n7047 GND.n7043 0.014
R8511 GND.n7047 GND.n7046 0.014
R8512 GND.n7014 GND.n7012 0.014
R8513 GND.n7021 GND.n7020 0.014
R8514 GND.n6993 GND.n6992 0.014
R8515 GND.n6805 GND.n6804 0.014
R8516 GND.n6810 GND.n6809 0.014
R8517 GND.n6809 GND.n6808 0.014
R8518 GND.n6779 GND.n6776 0.014
R8519 GND.n6726 GND.n6723 0.014
R8520 GND.n6815 GND.n6814 0.014
R8521 GND.n6820 GND.n6816 0.014
R8522 GND.n6820 GND.n6819 0.014
R8523 GND.n6787 GND.n6785 0.014
R8524 GND.n6794 GND.n6793 0.014
R8525 GND.n6766 GND.n6765 0.014
R8526 GND.n6473 GND.n6472 0.014
R8527 GND.n6478 GND.n6477 0.014
R8528 GND.n6477 GND.n6476 0.014
R8529 GND.n6458 GND.n6455 0.014
R8530 GND.n6442 GND.n6439 0.014
R8531 GND.n6483 GND.n6482 0.014
R8532 GND.n6488 GND.n6484 0.014
R8533 GND.n6488 GND.n6487 0.014
R8534 GND.n6390 GND.n6388 0.014
R8535 GND.n6397 GND.n6396 0.014
R8536 GND.n6408 GND.n6407 0.014
R8537 GND.n532 GND.n530 0.014
R8538 GND.n536 GND.n534 0.014
R8539 GND.n593 GND.n569 0.014
R8540 GND.n645 GND.n642 0.014
R8541 GND.n955 GND.n953 0.014
R8542 GND.n1025 GND.n1023 0.014
R8543 GND.n1061 GND.n1059 0.014
R8544 GND.n1066 GND.n1063 0.014
R8545 GND.n847 GND.n845 0.014
R8546 GND.n851 GND.n849 0.014
R8547 GND.n886 GND.n884 0.014
R8548 GND.n938 GND.n935 0.014
R8549 GND.n6001 GND.n5999 0.014
R8550 GND.n6005 GND.n6003 0.014
R8551 GND.n6063 GND.n6038 0.014
R8552 GND.n6115 GND.n6112 0.014
R8553 GND.n2577 GND.n2575 0.014
R8554 GND.n2647 GND.n2645 0.014
R8555 GND.n2683 GND.n2681 0.014
R8556 GND.n2688 GND.n2685 0.014
R8557 GND.n2469 GND.n2467 0.014
R8558 GND.n2473 GND.n2471 0.014
R8559 GND.n2508 GND.n2506 0.014
R8560 GND.n2560 GND.n2557 0.014
R8561 GND.n3829 GND.n3827 0.014
R8562 GND.n3833 GND.n3831 0.014
R8563 GND.n3891 GND.n3866 0.014
R8564 GND.n3943 GND.n3940 0.014
R8565 GND.n5502 GND.n5499 0.014
R8566 GND.n2298 GND.n2296 0.014
R8567 GND.n2302 GND.n2300 0.014
R8568 GND.n2359 GND.n2335 0.014
R8569 GND.n2411 GND.n2408 0.014
R8570 GND.n3004 GND.n3001 0.014
R8571 GND.n2952 GND.n2951 0.014
R8572 GND.n2924 GND.n2922 0.014
R8573 GND.n2920 GND.n2919 0.014
R8574 GND.n4115 GND.n4112 0.014
R8575 GND.n4063 GND.n4062 0.014
R8576 GND.n4035 GND.n4033 0.014
R8577 GND.n4031 GND.n4030 0.014
R8578 GND.n1583 GND.n1580 0.014
R8579 GND.n1531 GND.n1530 0.014
R8580 GND.n1497 GND.n1495 0.014
R8581 GND.n1493 GND.n1492 0.014
R8582 GND.n6176 GND.n6174 0.014
R8583 GND.n6227 GND.n6225 0.014
R8584 GND.n6262 GND.n6260 0.014
R8585 GND.n6267 GND.n6264 0.014
R8586 GND.n8231 GND.n8229 0.014
R8587 GND.n8242 GND.n8240 0.014
R8588 GND.n8246 GND.n8244 0.014
R8589 GND.n8277 GND.n8275 0.014
R8590 GND.n8159 GND.n8157 0.014
R8591 GND.n8170 GND.n8168 0.014
R8592 GND.n8174 GND.n8172 0.014
R8593 GND.n8204 GND.n8202 0.014
R8594 GND.n8338 GND.n8336 0.014
R8595 GND.n8349 GND.n8347 0.014
R8596 GND.n8353 GND.n8351 0.014
R8597 GND.n8384 GND.n8382 0.014
R8598 GND.n8410 GND.n8408 0.014
R8599 GND.n8421 GND.n8419 0.014
R8600 GND.n8425 GND.n8423 0.014
R8601 GND.n8455 GND.n8453 0.014
R8602 GND.n8523 GND.n8521 0.014
R8603 GND.n8534 GND.n8532 0.014
R8604 GND.n8538 GND.n8536 0.014
R8605 GND.n8569 GND.n8567 0.014
R8606 GND.n8595 GND.n8593 0.014
R8607 GND.n8606 GND.n8604 0.014
R8608 GND.n8610 GND.n8608 0.014
R8609 GND.n8640 GND.n8638 0.014
R8610 GND.n8708 GND.n8706 0.014
R8611 GND.n8719 GND.n8717 0.014
R8612 GND.n8723 GND.n8721 0.014
R8613 GND.n8754 GND.n8752 0.014
R8614 GND.n8780 GND.n8778 0.014
R8615 GND.n8791 GND.n8789 0.014
R8616 GND.n8795 GND.n8793 0.014
R8617 GND.n8825 GND.n8823 0.014
R8618 GND.n8893 GND.n8891 0.014
R8619 GND.n8904 GND.n8902 0.014
R8620 GND.n8908 GND.n8906 0.014
R8621 GND.n8939 GND.n8937 0.014
R8622 GND.n8965 GND.n8963 0.014
R8623 GND.n8976 GND.n8974 0.014
R8624 GND.n8980 GND.n8978 0.014
R8625 GND.n9010 GND.n9008 0.014
R8626 GND.n9078 GND.n9076 0.014
R8627 GND.n9089 GND.n9087 0.014
R8628 GND.n9093 GND.n9091 0.014
R8629 GND.n9124 GND.n9122 0.014
R8630 GND.n9150 GND.n9148 0.014
R8631 GND.n9161 GND.n9159 0.014
R8632 GND.n9165 GND.n9163 0.014
R8633 GND.n9195 GND.n9193 0.014
R8634 GND.n39 GND.n37 0.014
R8635 GND.n50 GND.n48 0.014
R8636 GND.n54 GND.n52 0.014
R8637 GND.n85 GND.n83 0.014
R8638 GND.n111 GND.n109 0.014
R8639 GND.n122 GND.n120 0.014
R8640 GND.n126 GND.n124 0.014
R8641 GND.n156 GND.n154 0.014
R8642 GND.n574 GND.n573 0.013
R8643 GND.n578 GND.n577 0.013
R8644 GND.n1009 GND.n1008 0.013
R8645 GND.n1005 GND.n1004 0.013
R8646 GND.n6044 GND.n6043 0.013
R8647 GND.n6048 GND.n6047 0.013
R8648 GND.n2631 GND.n2630 0.013
R8649 GND.n2627 GND.n2626 0.013
R8650 GND.n3872 GND.n3871 0.013
R8651 GND.n3876 GND.n3875 0.013
R8652 GND.n2340 GND.n2339 0.013
R8653 GND.n2344 GND.n2343 0.013
R8654 GND.n4004 GND.n4003 0.013
R8655 GND.n4008 GND.n4007 0.013
R8656 GND.n6300 GND.n6299 0.013
R8657 GND.n6304 GND.n6303 0.013
R8658 GND.n6362 GND.n6361 0.013
R8659 GND.n7971 GND.n7970 0.012
R8660 GND.n7964 GND.n7963 0.012
R8661 GND.n7744 GND.n7743 0.012
R8662 GND.n7737 GND.n7736 0.012
R8663 GND.n7517 GND.n7516 0.012
R8664 GND.n7510 GND.n7509 0.012
R8665 GND.n7290 GND.n7289 0.012
R8666 GND.n7283 GND.n7282 0.012
R8667 GND.n7063 GND.n7062 0.012
R8668 GND.n7056 GND.n7055 0.012
R8669 GND.n6836 GND.n6835 0.012
R8670 GND.n6829 GND.n6828 0.012
R8671 GND.n6504 GND.n6503 0.012
R8672 GND.n6497 GND.n6496 0.012
R8673 GND.n587 GND.n586 0.012
R8674 GND.n588 GND.n587 0.012
R8675 GND.n589 GND.n588 0.012
R8676 GND.n592 GND.n589 0.012
R8677 GND.n522 GND.n520 0.012
R8678 GND.n530 GND.n527 0.012
R8679 GND.n621 GND.n619 0.012
R8680 GND.n1758 GND.n1756 0.012
R8681 GND.n1618 GND.n1616 0.012
R8682 GND.n1310 GND.n1308 0.012
R8683 GND.n1451 GND.n1449 0.012
R8684 GND.n1253 GND.n1251 0.012
R8685 GND.n1113 GND.n1111 0.012
R8686 GND.n676 GND.n674 0.012
R8687 GND.n816 GND.n814 0.012
R8688 GND.n2738 GND.n2736 0.012
R8689 GND.n2878 GND.n2876 0.012
R8690 GND.n3181 GND.n3179 0.012
R8691 GND.n3041 GND.n3039 0.012
R8692 GND.n3771 GND.n3769 0.012
R8693 GND.n3631 GND.n3629 0.012
R8694 GND.n1020 GND.n1019 0.012
R8695 GND.n1019 GND.n1018 0.012
R8696 GND.n1018 GND.n1017 0.012
R8697 GND.n978 GND.n976 0.012
R8698 GND.n1067 GND.n1066 0.012
R8699 GND.n1074 GND.n1073 0.012
R8700 GND.n6057 GND.n6056 0.012
R8701 GND.n6058 GND.n6057 0.012
R8702 GND.n6059 GND.n6058 0.012
R8703 GND.n6062 GND.n6059 0.012
R8704 GND.n837 GND.n835 0.012
R8705 GND.n845 GND.n842 0.012
R8706 GND.n914 GND.n912 0.012
R8707 GND.n5991 GND.n5989 0.012
R8708 GND.n5999 GND.n5996 0.012
R8709 GND.n6091 GND.n6089 0.012
R8710 GND.n2642 GND.n2641 0.012
R8711 GND.n2641 GND.n2640 0.012
R8712 GND.n2640 GND.n2639 0.012
R8713 GND.n2600 GND.n2598 0.012
R8714 GND.n2689 GND.n2688 0.012
R8715 GND.n2696 GND.n2695 0.012
R8716 GND.n3885 GND.n3884 0.012
R8717 GND.n3886 GND.n3885 0.012
R8718 GND.n3887 GND.n3886 0.012
R8719 GND.n3890 GND.n3887 0.012
R8720 GND.n2459 GND.n2457 0.012
R8721 GND.n2467 GND.n2464 0.012
R8722 GND.n2536 GND.n2534 0.012
R8723 GND.n3819 GND.n3817 0.012
R8724 GND.n3827 GND.n3824 0.012
R8725 GND.n3919 GND.n3917 0.012
R8726 GND.n1854 GND.n1852 0.012
R8727 GND.n1994 GND.n1992 0.012
R8728 GND.n2034 GND.n2032 0.012
R8729 GND.n2174 GND.n2172 0.012
R8730 GND.n5164 GND.n5162 0.012
R8731 GND.n5304 GND.n5302 0.012
R8732 GND.n5344 GND.n5342 0.012
R8733 GND.n5484 GND.n5482 0.012
R8734 GND.n4414 GND.n4412 0.012
R8735 GND.n4554 GND.n4552 0.012
R8736 GND.n4594 GND.n4592 0.012
R8737 GND.n4740 GND.n4738 0.012
R8738 GND.n4785 GND.n4783 0.012
R8739 GND.n4925 GND.n4923 0.012
R8740 GND.n4965 GND.n4963 0.012
R8741 GND.n5105 GND.n5103 0.012
R8742 GND.n3565 GND.n3563 0.012
R8743 GND.n3418 GND.n3416 0.012
R8744 GND.n3378 GND.n3376 0.012
R8745 GND.n3237 GND.n3235 0.012
R8746 GND.n5860 GND.n5858 0.012
R8747 GND.n5720 GND.n5718 0.012
R8748 GND.n5680 GND.n5678 0.012
R8749 GND.n5539 GND.n5537 0.012
R8750 GND.n2353 GND.n2352 0.012
R8751 GND.n2354 GND.n2353 0.012
R8752 GND.n2355 GND.n2354 0.012
R8753 GND.n2358 GND.n2355 0.012
R8754 GND.n2288 GND.n2286 0.012
R8755 GND.n2296 GND.n2293 0.012
R8756 GND.n2387 GND.n2385 0.012
R8757 GND.n3992 GND.n3991 0.012
R8758 GND.n3993 GND.n3992 0.012
R8759 GND.n3994 GND.n3993 0.012
R8760 GND.n3995 GND.n3994 0.012
R8761 GND.n2980 GND.n2978 0.012
R8762 GND.n2919 GND.n2916 0.012
R8763 GND.n2911 GND.n2910 0.012
R8764 GND.n4091 GND.n4089 0.012
R8765 GND.n4030 GND.n4027 0.012
R8766 GND.n4022 GND.n4021 0.012
R8767 GND.n4143 GND.n4141 0.012
R8768 GND.n4283 GND.n4281 0.012
R8769 GND.n6288 GND.n6287 0.012
R8770 GND.n6289 GND.n6288 0.012
R8771 GND.n6290 GND.n6289 0.012
R8772 GND.n6291 GND.n6290 0.012
R8773 GND.n1559 GND.n1557 0.012
R8774 GND.n1492 GND.n1489 0.012
R8775 GND.n1484 GND.n1483 0.012
R8776 GND.n6199 GND.n6197 0.012
R8777 GND.n6268 GND.n6267 0.012
R8778 GND.n6275 GND.n6274 0.012
R8779 GND.n6338 GND.n6332 0.012
R8780 GND.n8120 GND.n8119 0.012
R8781 GND.n410 GND.n409 0.012
R8782 GND.n361 GND.n360 0.012
R8783 GND.n312 GND.n311 0.012
R8784 GND.n263 GND.n262 0.012
R8785 GND.n214 GND.n213 0.012
R8786 GND.n18 GND.n17 0.012
R8787 GND.n6335 GND.n6334 0.012
R8788 GND.n6330 GND.n6329 0.012
R8789 GND.n6331 GND.n6330 0.012
R8790 GND.n6337 GND.n6336 0.012
R8791 GND.n6332 GND.n6331 0.011
R8792 GND.n6336 GND.n6335 0.011
R8793 GND.n6329 GND.n6328 0.011
R8794 GND.n6334 GND.n6333 0.011
R8795 GND.n7946 GND.n7936 0.011
R8796 GND.n7885 GND.n7876 0.011
R8797 GND.n7719 GND.n7709 0.011
R8798 GND.n7658 GND.n7649 0.011
R8799 GND.n7492 GND.n7482 0.011
R8800 GND.n7431 GND.n7422 0.011
R8801 GND.n7265 GND.n7255 0.011
R8802 GND.n7204 GND.n7195 0.011
R8803 GND.n7038 GND.n7028 0.011
R8804 GND.n6977 GND.n6968 0.011
R8805 GND.n6811 GND.n6801 0.011
R8806 GND.n6750 GND.n6741 0.011
R8807 GND.n6430 GND.n6421 0.011
R8808 GND.n6041 GND.n6040 0.011
R8809 GND.n6043 GND.n6042 0.011
R8810 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/GATE GND.n1089 0.011
R8811 GND.n3869 GND.n3868 0.011
R8812 GND.n3871 GND.n3870 0.011
R8813 GND.n3787 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/GATE 0.011
R8814 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/GATE GND.n3786 0.011
R8815 GND.n4009 GND.n4008 0.011
R8816 GND.n4011 GND.n4010 0.011
R8817 GND.n6305 GND.n6304 0.011
R8818 GND.n6307 GND.n6306 0.011
R8819 GND.n8092 GND.n8091 0.011
R8820 GND.n8094 GND.n8093 0.011
R8821 GND.n429 GND.n428 0.011
R8822 GND.n431 GND.n430 0.011
R8823 GND.n447 GND.n446 0.011
R8824 GND.n380 GND.n379 0.011
R8825 GND.n382 GND.n381 0.011
R8826 GND.n398 GND.n397 0.011
R8827 GND.n331 GND.n330 0.011
R8828 GND.n333 GND.n332 0.011
R8829 GND.n349 GND.n348 0.011
R8830 GND.n282 GND.n281 0.011
R8831 GND.n284 GND.n283 0.011
R8832 GND.n300 GND.n299 0.011
R8833 GND.n233 GND.n232 0.011
R8834 GND.n235 GND.n234 0.011
R8835 GND.n251 GND.n250 0.011
R8836 GND.n1 GND.n0 0.011
R8837 GND.n3 GND.n2 0.011
R8838 GND.n15 GND.n14 0.011
R8839 GND.n3803 GND.n3802 0.01
R8840 GND.n3790 GND.n3787 0.01
R8841 GND.n6479 GND.n6469 0.01
R8842 GND.n573 GND.n572 0.01
R8843 GND.n575 GND.n574 0.01
R8844 GND.n577 GND.n576 0.01
R8845 GND.n586 GND.n585 0.01
R8846 GND.n1720 GND.n1718 0.01
R8847 GND.n1662 GND.n1654 0.01
R8848 GND.n1354 GND.n1346 0.01
R8849 GND.n1412 GND.n1410 0.01
R8850 GND.n1215 GND.n1213 0.01
R8851 GND.n1157 GND.n1149 0.01
R8852 GND.n720 GND.n712 0.01
R8853 GND.n778 GND.n776 0.01
R8854 GND.n2782 GND.n2774 0.01
R8855 GND.n2840 GND.n2838 0.01
R8856 GND.n3143 GND.n3141 0.01
R8857 GND.n3085 GND.n3077 0.01
R8858 GND.n3733 GND.n3731 0.01
R8859 GND.n3675 GND.n3667 0.01
R8860 GND.n1017 GND.n1016 0.01
R8861 GND.n1008 GND.n1007 0.01
R8862 GND.n1006 GND.n1005 0.01
R8863 GND.n1004 GND.n1003 0.01
R8864 GND.n1002 GND.n1001 0.01
R8865 GND.n6045 GND.n6044 0.01
R8866 GND.n6047 GND.n6046 0.01
R8867 GND.n6056 GND.n6055 0.01
R8868 GND.n2639 GND.n2638 0.01
R8869 GND.n2630 GND.n2629 0.01
R8870 GND.n2628 GND.n2627 0.01
R8871 GND.n2626 GND.n2625 0.01
R8872 GND.n2624 GND.n2623 0.01
R8873 GND.n3873 GND.n3872 0.01
R8874 GND.n3875 GND.n3874 0.01
R8875 GND.n3884 GND.n3883 0.01
R8876 GND.n1898 GND.n1890 0.01
R8877 GND.n1956 GND.n1954 0.01
R8878 GND.n2078 GND.n2070 0.01
R8879 GND.n2136 GND.n2134 0.01
R8880 GND.n5511 GND.n5510 0.01
R8881 GND.n5208 GND.n5200 0.01
R8882 GND.n5266 GND.n5264 0.01
R8883 GND.n5388 GND.n5380 0.01
R8884 GND.n5446 GND.n5444 0.01
R8885 GND.n4458 GND.n4450 0.01
R8886 GND.n4516 GND.n4514 0.01
R8887 GND.n4639 GND.n4631 0.01
R8888 GND.n4700 GND.n4698 0.01
R8889 GND.n4829 GND.n4821 0.01
R8890 GND.n4887 GND.n4885 0.01
R8891 GND.n5009 GND.n5001 0.01
R8892 GND.n5067 GND.n5065 0.01
R8893 GND.n3525 GND.n3523 0.01
R8894 GND.n3464 GND.n3456 0.01
R8895 GND.n3340 GND.n3338 0.01
R8896 GND.n3282 GND.n3274 0.01
R8897 GND.n5822 GND.n5820 0.01
R8898 GND.n5764 GND.n5756 0.01
R8899 GND.n5642 GND.n5640 0.01
R8900 GND.n5584 GND.n5576 0.01
R8901 GND.n2339 GND.n2338 0.01
R8902 GND.n2341 GND.n2340 0.01
R8903 GND.n2343 GND.n2342 0.01
R8904 GND.n2352 GND.n2351 0.01
R8905 GND.n3996 GND.n3995 0.01
R8906 GND.n4005 GND.n4004 0.01
R8907 GND.n4007 GND.n4006 0.01
R8908 GND.n4187 GND.n4179 0.01
R8909 GND.n4245 GND.n4243 0.01
R8910 GND.n6292 GND.n6291 0.01
R8911 GND.n6301 GND.n6300 0.01
R8912 GND.n6303 GND.n6302 0.01
R8913 GND.n169 GND.n24 0.01
R8914 GND.n9236 GND.n9235 0.01
R8915 GND.n9051 GND.n9050 0.01
R8916 GND.n8866 GND.n8865 0.01
R8917 GND.n8681 GND.n8680 0.01
R8918 GND.n8496 GND.n8495 0.01
R8919 GND.n8311 GND.n8310 0.01
R8920 GND.n6924 GND.n6923 0.01
R8921 GND.n7151 GND.n7150 0.01
R8922 GND.n7378 GND.n7377 0.01
R8923 GND.n7605 GND.n7604 0.01
R8924 GND.n7832 GND.n7831 0.01
R8925 GND.n8059 GND.n8058 0.01
R8926 GND.n7843 GND.n7841 0.009
R8927 GND.n7848 GND.n7845 0.009
R8928 GND.n7881 GND.n7880 0.009
R8929 GND.n8021 GND.n8019 0.009
R8930 GND.n8029 GND.n8027 0.009
R8931 GND.n7875 GND.n7873 0.009
R8932 GND.n7973 GND.n7972 0.009
R8933 GND.n7984 GND.n7974 0.009
R8934 GND.n8014 GND.n8013 0.009
R8935 GND.n8016 GND.n8015 0.009
R8936 GND.n7932 GND.n7931 0.009
R8937 GND.n7906 GND.n7905 0.009
R8938 GND.n7902 GND.n7890 0.009
R8939 GND.n7616 GND.n7614 0.009
R8940 GND.n7621 GND.n7618 0.009
R8941 GND.n7654 GND.n7653 0.009
R8942 GND.n7794 GND.n7792 0.009
R8943 GND.n7802 GND.n7800 0.009
R8944 GND.n7648 GND.n7646 0.009
R8945 GND.n7746 GND.n7745 0.009
R8946 GND.n7757 GND.n7747 0.009
R8947 GND.n7787 GND.n7786 0.009
R8948 GND.n7789 GND.n7788 0.009
R8949 GND.n7705 GND.n7704 0.009
R8950 GND.n7679 GND.n7678 0.009
R8951 GND.n7675 GND.n7663 0.009
R8952 GND.n7389 GND.n7387 0.009
R8953 GND.n7394 GND.n7391 0.009
R8954 GND.n7427 GND.n7426 0.009
R8955 GND.n7567 GND.n7565 0.009
R8956 GND.n7575 GND.n7573 0.009
R8957 GND.n7421 GND.n7419 0.009
R8958 GND.n7519 GND.n7518 0.009
R8959 GND.n7530 GND.n7520 0.009
R8960 GND.n7560 GND.n7559 0.009
R8961 GND.n7562 GND.n7561 0.009
R8962 GND.n7478 GND.n7477 0.009
R8963 GND.n7452 GND.n7451 0.009
R8964 GND.n7448 GND.n7436 0.009
R8965 GND.n7162 GND.n7160 0.009
R8966 GND.n7167 GND.n7164 0.009
R8967 GND.n7200 GND.n7199 0.009
R8968 GND.n7340 GND.n7338 0.009
R8969 GND.n7348 GND.n7346 0.009
R8970 GND.n7194 GND.n7192 0.009
R8971 GND.n7292 GND.n7291 0.009
R8972 GND.n7303 GND.n7293 0.009
R8973 GND.n7333 GND.n7332 0.009
R8974 GND.n7335 GND.n7334 0.009
R8975 GND.n7251 GND.n7250 0.009
R8976 GND.n7225 GND.n7224 0.009
R8977 GND.n7221 GND.n7209 0.009
R8978 GND.n6935 GND.n6933 0.009
R8979 GND.n6940 GND.n6937 0.009
R8980 GND.n6973 GND.n6972 0.009
R8981 GND.n7113 GND.n7111 0.009
R8982 GND.n7121 GND.n7119 0.009
R8983 GND.n6967 GND.n6965 0.009
R8984 GND.n7065 GND.n7064 0.009
R8985 GND.n7076 GND.n7066 0.009
R8986 GND.n7106 GND.n7105 0.009
R8987 GND.n7108 GND.n7107 0.009
R8988 GND.n7024 GND.n7023 0.009
R8989 GND.n6998 GND.n6997 0.009
R8990 GND.n6994 GND.n6982 0.009
R8991 GND.n6708 GND.n6706 0.009
R8992 GND.n6713 GND.n6710 0.009
R8993 GND.n6746 GND.n6745 0.009
R8994 GND.n6886 GND.n6884 0.009
R8995 GND.n6894 GND.n6892 0.009
R8996 GND.n6740 GND.n6738 0.009
R8997 GND.n6838 GND.n6837 0.009
R8998 GND.n6849 GND.n6839 0.009
R8999 GND.n6879 GND.n6878 0.009
R9000 GND.n6881 GND.n6880 0.009
R9001 GND.n6797 GND.n6796 0.009
R9002 GND.n6771 GND.n6770 0.009
R9003 GND.n6767 GND.n6755 0.009
R9004 GND.n6376 GND.n6374 0.009
R9005 GND.n6381 GND.n6378 0.009
R9006 GND.n6426 GND.n6425 0.009
R9007 GND.n6554 GND.n6552 0.009
R9008 GND.n6562 GND.n6560 0.009
R9009 GND.n6420 GND.n6419 0.009
R9010 GND.n6506 GND.n6505 0.009
R9011 GND.n6517 GND.n6507 0.009
R9012 GND.n6547 GND.n6546 0.009
R9013 GND.n6549 GND.n6548 0.009
R9014 GND.n6465 GND.n6464 0.009
R9015 GND.n6450 GND.n6449 0.009
R9016 GND.n6446 GND.n6445 0.009
R9017 GND.n592 GND.n591 0.009
R9018 GND.n511 GND.n509 0.009
R9019 GND.n543 GND.n541 0.009
R9020 GND.n547 GND.n545 0.009
R9021 GND.n651 GND.n649 0.009
R9022 GND.n948 GND.n946 0.009
R9023 GND.n1050 GND.n1048 0.009
R9024 GND.n1055 GND.n1052 0.009
R9025 GND.n1086 GND.n1084 0.009
R9026 GND.n6062 GND.n6061 0.009
R9027 GND.n826 GND.n824 0.009
R9028 GND.n858 GND.n856 0.009
R9029 GND.n862 GND.n860 0.009
R9030 GND.n944 GND.n942 0.009
R9031 GND.n5980 GND.n5978 0.009
R9032 GND.n6012 GND.n6010 0.009
R9033 GND.n6016 GND.n6014 0.009
R9034 GND.n6121 GND.n6119 0.009
R9035 GND.n1267 GND.n1265 0.009
R9036 GND.n2570 GND.n2568 0.009
R9037 GND.n2672 GND.n2670 0.009
R9038 GND.n2677 GND.n2674 0.009
R9039 GND.n2708 GND.n2706 0.009
R9040 GND.n3890 GND.n3889 0.009
R9041 GND.n2448 GND.n2446 0.009
R9042 GND.n2480 GND.n2478 0.009
R9043 GND.n2484 GND.n2482 0.009
R9044 GND.n2566 GND.n2564 0.009
R9045 GND.n3808 GND.n3806 0.009
R9046 GND.n3840 GND.n3838 0.009
R9047 GND.n3844 GND.n3842 0.009
R9048 GND.n3949 GND.n3947 0.009
R9049 GND.n2358 GND.n2357 0.009
R9050 GND.n2277 GND.n2275 0.009
R9051 GND.n2309 GND.n2307 0.009
R9052 GND.n2313 GND.n2311 0.009
R9053 GND.n2417 GND.n2415 0.009
R9054 GND.n3991 GND.n3990 0.009
R9055 GND.n3010 GND.n3008 0.009
R9056 GND.n2934 GND.n2932 0.009
R9057 GND.n2930 GND.n2929 0.009
R9058 GND.n2901 GND.n2900 0.009
R9059 GND.n4121 GND.n4119 0.009
R9060 GND.n4045 GND.n4043 0.009
R9061 GND.n4041 GND.n4040 0.009
R9062 GND.n4012 GND.n3988 0.009
R9063 GND.n6287 GND.n6286 0.009
R9064 GND.n1589 GND.n1587 0.009
R9065 GND.n1508 GND.n1506 0.009
R9066 GND.n1504 GND.n1502 0.009
R9067 GND.n1474 GND.n1473 0.009
R9068 GND.n6169 GND.n6167 0.009
R9069 GND.n6251 GND.n6249 0.009
R9070 GND.n6256 GND.n6253 0.009
R9071 GND.n6310 GND.n6308 0.009
R9072 GND.n8220 GND.n8218 0.009
R9073 GND.n8248 GND.n8247 0.009
R9074 GND.n8253 GND.n8251 0.009
R9075 GND.n8257 GND.n8255 0.009
R9076 GND.n8148 GND.n8146 0.009
R9077 GND.n8176 GND.n8175 0.009
R9078 GND.n8181 GND.n8179 0.009
R9079 GND.n8185 GND.n8183 0.009
R9080 GND.n8106 GND.n8105 0.009
R9081 GND.n8108 GND.n8107 0.009
R9082 GND.n8118 GND.n8117 0.009
R9083 GND.n8327 GND.n8325 0.009
R9084 GND.n8355 GND.n8354 0.009
R9085 GND.n8360 GND.n8358 0.009
R9086 GND.n8364 GND.n8362 0.009
R9087 GND.n8399 GND.n8397 0.009
R9088 GND.n8427 GND.n8426 0.009
R9089 GND.n8432 GND.n8430 0.009
R9090 GND.n8436 GND.n8434 0.009
R9091 GND.n442 GND.n441 0.009
R9092 GND.n444 GND.n443 0.009
R9093 GND.n8512 GND.n8510 0.009
R9094 GND.n8540 GND.n8539 0.009
R9095 GND.n8545 GND.n8543 0.009
R9096 GND.n8549 GND.n8547 0.009
R9097 GND.n8584 GND.n8582 0.009
R9098 GND.n8612 GND.n8611 0.009
R9099 GND.n8617 GND.n8615 0.009
R9100 GND.n8621 GND.n8619 0.009
R9101 GND.n393 GND.n392 0.009
R9102 GND.n395 GND.n394 0.009
R9103 GND.n8697 GND.n8695 0.009
R9104 GND.n8725 GND.n8724 0.009
R9105 GND.n8730 GND.n8728 0.009
R9106 GND.n8734 GND.n8732 0.009
R9107 GND.n8769 GND.n8767 0.009
R9108 GND.n8797 GND.n8796 0.009
R9109 GND.n8802 GND.n8800 0.009
R9110 GND.n8806 GND.n8804 0.009
R9111 GND.n344 GND.n343 0.009
R9112 GND.n346 GND.n345 0.009
R9113 GND.n8882 GND.n8880 0.009
R9114 GND.n8910 GND.n8909 0.009
R9115 GND.n8915 GND.n8913 0.009
R9116 GND.n8919 GND.n8917 0.009
R9117 GND.n8954 GND.n8952 0.009
R9118 GND.n8982 GND.n8981 0.009
R9119 GND.n8987 GND.n8985 0.009
R9120 GND.n8991 GND.n8989 0.009
R9121 GND.n295 GND.n294 0.009
R9122 GND.n297 GND.n296 0.009
R9123 GND.n9067 GND.n9065 0.009
R9124 GND.n9095 GND.n9094 0.009
R9125 GND.n9100 GND.n9098 0.009
R9126 GND.n9104 GND.n9102 0.009
R9127 GND.n9139 GND.n9137 0.009
R9128 GND.n9167 GND.n9166 0.009
R9129 GND.n9172 GND.n9170 0.009
R9130 GND.n9176 GND.n9174 0.009
R9131 GND.n246 GND.n245 0.009
R9132 GND.n248 GND.n247 0.009
R9133 GND.n28 GND.n26 0.009
R9134 GND.n56 GND.n55 0.009
R9135 GND.n61 GND.n59 0.009
R9136 GND.n65 GND.n63 0.009
R9137 GND.n100 GND.n98 0.009
R9138 GND.n128 GND.n127 0.009
R9139 GND.n133 GND.n131 0.009
R9140 GND.n137 GND.n135 0.009
R9141 GND.n9 GND.n8 0.009
R9142 GND.n10 GND.n9 0.009
R9143 GND.n12 GND.n11 0.009
R9144 GND.n16 GND.n15 0.009
R9145 GND.n8030 GND.n8016 0.008
R9146 GND.n7930 GND.n7918 0.008
R9147 GND.n7803 GND.n7789 0.008
R9148 GND.n7703 GND.n7691 0.008
R9149 GND.n7576 GND.n7562 0.008
R9150 GND.n7476 GND.n7464 0.008
R9151 GND.n7349 GND.n7335 0.008
R9152 GND.n7249 GND.n7237 0.008
R9153 GND.n7122 GND.n7108 0.008
R9154 GND.n7022 GND.n7010 0.008
R9155 GND.n6895 GND.n6881 0.008
R9156 GND.n6795 GND.n6783 0.008
R9157 GND.n6563 GND.n6549 0.008
R9158 GND.n6463 GND.n6462 0.008
R9159 GND.n579 GND.n578 0.008
R9160 GND.n583 GND.n582 0.008
R9161 GND.n1770 GND.n1768 0.008
R9162 GND.n1605 GND.n1603 0.008
R9163 GND.n1297 GND.n1288 0.008
R9164 GND.n1463 GND.n1461 0.008
R9165 GND.n1256 GND.n1255 0.008
R9166 GND.n1101 GND.n821 0.008
R9167 GND.n6160 GND.n6158 0.008
R9168 GND.n819 GND.n818 0.008
R9169 GND.n2725 GND.n2712 0.008
R9170 GND.n2890 GND.n2888 0.008
R9171 GND.n3193 GND.n3191 0.008
R9172 GND.n3028 GND.n3026 0.008
R9173 GND.n3774 GND.n3773 0.008
R9174 GND.n3619 GND.n2443 0.008
R9175 GND.n1014 GND.n1013 0.008
R9176 GND.n1010 GND.n1009 0.008
R9177 GND.n6049 GND.n6048 0.008
R9178 GND.n6053 GND.n6052 0.008
R9179 GND.n2636 GND.n2635 0.008
R9180 GND.n2632 GND.n2631 0.008
R9181 GND.n3877 GND.n3876 0.008
R9182 GND.n3881 GND.n3880 0.008
R9183 GND.n1849 GND.n1848 0.008
R9184 GND.n2006 GND.n2004 0.008
R9185 GND.n2022 GND.n2020 0.008
R9186 GND.n2177 GND.n2176 0.008
R9187 GND.n5159 GND.n5158 0.008
R9188 GND.n5316 GND.n5314 0.008
R9189 GND.n5332 GND.n5330 0.008
R9190 GND.n5487 GND.n5486 0.008
R9191 GND.n4409 GND.n4408 0.008
R9192 GND.n4566 GND.n4564 0.008
R9193 GND.n4582 GND.n4580 0.008
R9194 GND.n4743 GND.n4742 0.008
R9195 GND.n4780 GND.n4779 0.008
R9196 GND.n4937 GND.n4935 0.008
R9197 GND.n4953 GND.n4951 0.008
R9198 GND.n5108 GND.n5107 0.008
R9199 GND.n3568 GND.n3567 0.008
R9200 GND.n3406 GND.n3404 0.008
R9201 GND.n3390 GND.n3388 0.008
R9202 GND.n3232 GND.n3231 0.008
R9203 GND.n3596 GND.n3595 0.008
R9204 GND.n5863 GND.n5862 0.008
R9205 GND.n5708 GND.n5706 0.008
R9206 GND.n5692 GND.n5690 0.008
R9207 GND.n5534 GND.n5533 0.008
R9208 GND.n3227 GND.n3226 0.008
R9209 GND.n2345 GND.n2344 0.008
R9210 GND.n2349 GND.n2348 0.008
R9211 GND.n3999 GND.n3998 0.008
R9212 GND.n4003 GND.n4002 0.008
R9213 GND.n4130 GND.n4128 0.008
R9214 GND.n4295 GND.n4293 0.008
R9215 GND.n6295 GND.n6294 0.008
R9216 GND.n6299 GND.n6298 0.008
R9217 GND.n6338 GND.n6337 0.008
R9218 GND.n8126 GND.n8125 0.008
R9219 GND.n8477 GND.n8476 0.008
R9220 GND.n8662 GND.n8661 0.008
R9221 GND.n8847 GND.n8846 0.008
R9222 GND.n9032 GND.n9031 0.008
R9223 GND.n9217 GND.n9216 0.008
R9224 GND.n9262 GND.n9261 0.008
R9225 GND.n479 GND.n478 0.008
R9226 GND.n2196 GND.n2195 0.008
R9227 GND.n4359 GND.n4358 0.008
R9228 GND.n7976 GND.n7975 0.007
R9229 GND.n7986 GND.n7985 0.007
R9230 GND.n7934 GND.n7933 0.007
R9231 GND.n7933 GND.n7932 0.007
R9232 GND.n7749 GND.n7748 0.007
R9233 GND.n7759 GND.n7758 0.007
R9234 GND.n7707 GND.n7706 0.007
R9235 GND.n7706 GND.n7705 0.007
R9236 GND.n7522 GND.n7521 0.007
R9237 GND.n7532 GND.n7531 0.007
R9238 GND.n7480 GND.n7479 0.007
R9239 GND.n7479 GND.n7478 0.007
R9240 GND.n7295 GND.n7294 0.007
R9241 GND.n7305 GND.n7304 0.007
R9242 GND.n7253 GND.n7252 0.007
R9243 GND.n7252 GND.n7251 0.007
R9244 GND.n7068 GND.n7067 0.007
R9245 GND.n7078 GND.n7077 0.007
R9246 GND.n7026 GND.n7025 0.007
R9247 GND.n7025 GND.n7024 0.007
R9248 GND.n6841 GND.n6840 0.007
R9249 GND.n6851 GND.n6850 0.007
R9250 GND.n6799 GND.n6798 0.007
R9251 GND.n6798 GND.n6797 0.007
R9252 GND.n6509 GND.n6508 0.007
R9253 GND.n6519 GND.n6518 0.007
R9254 GND.n6467 GND.n6466 0.007
R9255 GND.n6466 GND.n6465 0.007
R9256 GND.n512 GND.n511 0.007
R9257 GND.n614 GND.n612 0.007
R9258 GND.n985 GND.n983 0.007
R9259 GND.n1084 GND.n1082 0.007
R9260 GND.n827 GND.n826 0.007
R9261 GND.n907 GND.n905 0.007
R9262 GND.n5981 GND.n5980 0.007
R9263 GND.n6084 GND.n6082 0.007
R9264 GND.n5975 GND.n1286 0.007
R9265 GND.n2607 GND.n2605 0.007
R9266 GND.n2706 GND.n2704 0.007
R9267 GND.n2449 GND.n2448 0.007
R9268 GND.n2529 GND.n2527 0.007
R9269 GND.n3809 GND.n3808 0.007
R9270 GND.n3912 GND.n3910 0.007
R9271 GND.n2184 GND.n2183 0.007
R9272 GND.n2186 GND.n2185 0.007
R9273 GND.n2187 GND.n2186 0.007
R9274 GND.n2189 GND.n2188 0.007
R9275 GND.n4388 GND.n2192 0.007
R9276 GND.n4388 GND.n2194 0.007
R9277 GND.n4396 GND.n4395 0.007
R9278 GND.n4394 GND.n4393 0.007
R9279 GND.n4393 GND.n4392 0.007
R9280 GND.n4391 GND.n4390 0.007
R9281 GND.n2214 GND.n2213 0.007
R9282 GND.n2212 GND.n2211 0.007
R9283 GND.n2211 GND.n2209 0.007
R9284 GND.n2238 GND.n2235 0.007
R9285 GND.n2238 GND.n2236 0.007
R9286 GND.n4309 GND.n2248 0.007
R9287 GND.n4309 GND.n2249 0.007
R9288 GND.n4315 GND.n4313 0.007
R9289 GND.n4330 GND.n4328 0.007
R9290 GND.n4331 GND.n4330 0.007
R9291 GND.n4333 GND.n4332 0.007
R9292 GND.n2278 GND.n2277 0.007
R9293 GND.n2380 GND.n2378 0.007
R9294 GND.n2973 GND.n2971 0.007
R9295 GND.n2902 GND.n2901 0.007
R9296 GND.n4084 GND.n4082 0.007
R9297 GND.n4013 GND.n4012 0.007
R9298 GND.n1552 GND.n1550 0.007
R9299 GND.n1475 GND.n1474 0.007
R9300 GND.n6206 GND.n6204 0.007
R9301 GND.n6308 GND.n6283 0.007
R9302 GND.n6339 GND.n488 0.007
R9303 GND.n6344 GND.n6343 0.007
R9304 GND.n6350 GND.n6348 0.007
R9305 GND.n6350 GND.n6349 0.007
R9306 GND.n6357 GND.n6355 0.007
R9307 GND.n6357 GND.n6356 0.007
R9308 GND.n473 GND.n471 0.007
R9309 GND.n473 GND.n472 0.007
R9310 GND.n454 GND.n453 0.007
R9311 GND.n455 GND.n454 0.007
R9312 GND.n457 GND.n456 0.007
R9313 GND.n8221 GND.n8220 0.007
R9314 GND.n8149 GND.n8148 0.007
R9315 GND.n8095 GND.n8094 0.007
R9316 GND.n8289 GND.n8144 0.007
R9317 GND.n8139 GND.n8138 0.007
R9318 GND.n8328 GND.n8327 0.007
R9319 GND.n8400 GND.n8399 0.007
R9320 GND.n432 GND.n431 0.007
R9321 GND.n8487 GND.n8486 0.007
R9322 GND.n8513 GND.n8512 0.007
R9323 GND.n8585 GND.n8584 0.007
R9324 GND.n383 GND.n382 0.007
R9325 GND.n8672 GND.n8671 0.007
R9326 GND.n8698 GND.n8697 0.007
R9327 GND.n8770 GND.n8769 0.007
R9328 GND.n334 GND.n333 0.007
R9329 GND.n8857 GND.n8856 0.007
R9330 GND.n8883 GND.n8882 0.007
R9331 GND.n8955 GND.n8954 0.007
R9332 GND.n285 GND.n284 0.007
R9333 GND.n9042 GND.n9041 0.007
R9334 GND.n9068 GND.n9067 0.007
R9335 GND.n9140 GND.n9139 0.007
R9336 GND.n236 GND.n235 0.007
R9337 GND.n9227 GND.n9226 0.007
R9338 GND.n29 GND.n28 0.007
R9339 GND.n101 GND.n100 0.007
R9340 GND.n4 GND.n3 0.007
R9341 GND.n22 GND.n21 0.007
R9342 GND.n170 GND.n169 0.007
R9343 GND.n175 GND.n174 0.007
R9344 GND.n178 GND.n177 0.007
R9345 GND.n7931 GND.n7930 0.006
R9346 GND.n7887 GND.n7886 0.006
R9347 GND.n7704 GND.n7703 0.006
R9348 GND.n7660 GND.n7659 0.006
R9349 GND.n7477 GND.n7476 0.006
R9350 GND.n7433 GND.n7432 0.006
R9351 GND.n7250 GND.n7249 0.006
R9352 GND.n7206 GND.n7205 0.006
R9353 GND.n7023 GND.n7022 0.006
R9354 GND.n6979 GND.n6978 0.006
R9355 GND.n6796 GND.n6795 0.006
R9356 GND.n6752 GND.n6751 0.006
R9357 GND.n6464 GND.n6463 0.006
R9358 GND.n6432 GND.n6431 0.006
R9359 GND.n580 GND.n579 0.006
R9360 GND.n582 GND.n581 0.006
R9361 GND.n1708 GND.n1706 0.006
R9362 GND.n1674 GND.n1666 0.006
R9363 GND.n1366 GND.n1358 0.006
R9364 GND.n1400 GND.n1398 0.006
R9365 GND.n1203 GND.n1201 0.006
R9366 GND.n1169 GND.n1161 0.006
R9367 GND.n732 GND.n724 0.006
R9368 GND.n766 GND.n764 0.006
R9369 GND.n2794 GND.n2786 0.006
R9370 GND.n2828 GND.n2826 0.006
R9371 GND.n3131 GND.n3129 0.006
R9372 GND.n3097 GND.n3089 0.006
R9373 GND.n3721 GND.n3719 0.006
R9374 GND.n3687 GND.n3679 0.006
R9375 GND.n1013 GND.n1012 0.006
R9376 GND.n1011 GND.n1010 0.006
R9377 GND.n6050 GND.n6049 0.006
R9378 GND.n6052 GND.n6051 0.006
R9379 GND.n2635 GND.n2634 0.006
R9380 GND.n2633 GND.n2632 0.006
R9381 GND.n3878 GND.n3877 0.006
R9382 GND.n3880 GND.n3879 0.006
R9383 GND.n1910 GND.n1902 0.006
R9384 GND.n1944 GND.n1942 0.006
R9385 GND.n2090 GND.n2082 0.006
R9386 GND.n2124 GND.n2122 0.006
R9387 GND.n2185 GND.n2184 0.006
R9388 GND.n2188 GND.n2187 0.006
R9389 GND.n2192 GND.n2191 0.006
R9390 GND.n2194 GND.n2193 0.006
R9391 GND.n4395 GND.n4394 0.006
R9392 GND.n4392 GND.n4391 0.006
R9393 GND.n5220 GND.n5212 0.006
R9394 GND.n5254 GND.n5252 0.006
R9395 GND.n5400 GND.n5392 0.006
R9396 GND.n5434 GND.n5432 0.006
R9397 GND.n4470 GND.n4462 0.006
R9398 GND.n4504 GND.n4502 0.006
R9399 GND.n4652 GND.n4643 0.006
R9400 GND.n4688 GND.n4686 0.006
R9401 GND.n4841 GND.n4833 0.006
R9402 GND.n4875 GND.n4873 0.006
R9403 GND.n5021 GND.n5013 0.006
R9404 GND.n5055 GND.n5053 0.006
R9405 GND.n3513 GND.n3511 0.006
R9406 GND.n3477 GND.n3468 0.006
R9407 GND.n3328 GND.n3326 0.006
R9408 GND.n3294 GND.n3286 0.006
R9409 GND.n5810 GND.n5808 0.006
R9410 GND.n5776 GND.n5768 0.006
R9411 GND.n5630 GND.n5628 0.006
R9412 GND.n5596 GND.n5588 0.006
R9413 GND.n2213 GND.n2212 0.006
R9414 GND.n4328 GND.n4327 0.006
R9415 GND.n4332 GND.n4331 0.006
R9416 GND.n2346 GND.n2345 0.006
R9417 GND.n2348 GND.n2347 0.006
R9418 GND.n4000 GND.n3999 0.006
R9419 GND.n4002 GND.n4001 0.006
R9420 GND.n4199 GND.n4191 0.006
R9421 GND.n4233 GND.n4231 0.006
R9422 GND.n6296 GND.n6295 0.006
R9423 GND.n6298 GND.n6297 0.006
R9424 GND.n6326 GND.n6325 0.006
R9425 GND.n488 GND.n487 0.006
R9426 GND.n456 GND.n455 0.006
R9427 GND.n8096 GND.n8095 0.006
R9428 GND.n8097 GND.n8096 0.006
R9429 GND.n8296 GND.n8295 0.006
R9430 GND.n8140 GND.n8139 0.006
R9431 GND.n8127 GND.n8126 0.006
R9432 GND.n433 GND.n432 0.006
R9433 GND.n434 GND.n433 0.006
R9434 GND.n418 GND.n417 0.006
R9435 GND.n8488 GND.n8487 0.006
R9436 GND.n8478 GND.n8477 0.006
R9437 GND.n384 GND.n383 0.006
R9438 GND.n385 GND.n384 0.006
R9439 GND.n369 GND.n368 0.006
R9440 GND.n8673 GND.n8672 0.006
R9441 GND.n8663 GND.n8662 0.006
R9442 GND.n335 GND.n334 0.006
R9443 GND.n336 GND.n335 0.006
R9444 GND.n320 GND.n319 0.006
R9445 GND.n8858 GND.n8857 0.006
R9446 GND.n8848 GND.n8847 0.006
R9447 GND.n286 GND.n285 0.006
R9448 GND.n287 GND.n286 0.006
R9449 GND.n271 GND.n270 0.006
R9450 GND.n9043 GND.n9042 0.006
R9451 GND.n9033 GND.n9032 0.006
R9452 GND.n237 GND.n236 0.006
R9453 GND.n238 GND.n237 0.006
R9454 GND.n222 GND.n221 0.006
R9455 GND.n9228 GND.n9227 0.006
R9456 GND.n9218 GND.n9217 0.006
R9457 GND.n5 GND.n4 0.006
R9458 GND.n6 GND.n5 0.006
R9459 GND.n23 GND.n22 0.006
R9460 GND.n173 GND.n172 0.006
R9461 GND.n174 GND.n173 0.006
R9462 GND.n9261 GND.n9260 0.006
R9463 GND.n6579 GND.n6578 0.006
R9464 GND.n8031 GND.n8030 0.006
R9465 GND.n7804 GND.n7803 0.006
R9466 GND.n7577 GND.n7576 0.006
R9467 GND.n7350 GND.n7349 0.006
R9468 GND.n7123 GND.n7122 0.006
R9469 GND.n6896 GND.n6895 0.006
R9470 GND.n6564 GND.n6563 0.006
R9471 GND.n7993 GND.n7992 0.005
R9472 GND.n7994 GND.n7993 0.005
R9473 GND.n7904 GND.n7903 0.005
R9474 GND.n7766 GND.n7765 0.005
R9475 GND.n7767 GND.n7766 0.005
R9476 GND.n7677 GND.n7676 0.005
R9477 GND.n7539 GND.n7538 0.005
R9478 GND.n7540 GND.n7539 0.005
R9479 GND.n7450 GND.n7449 0.005
R9480 GND.n7312 GND.n7311 0.005
R9481 GND.n7313 GND.n7312 0.005
R9482 GND.n7223 GND.n7222 0.005
R9483 GND.n7085 GND.n7084 0.005
R9484 GND.n7086 GND.n7085 0.005
R9485 GND.n6996 GND.n6995 0.005
R9486 GND.n6858 GND.n6857 0.005
R9487 GND.n6859 GND.n6858 0.005
R9488 GND.n6769 GND.n6768 0.005
R9489 GND.n6526 GND.n6525 0.005
R9490 GND.n6527 GND.n6526 0.005
R9491 GND.n6448 GND.n6447 0.005
R9492 GND.n8137 GND.n8136 0.005
R9493 GND.n8130 GND.n8129 0.005
R9494 GND.n8102 GND.n8101 0.005
R9495 GND.n8109 GND.n8104 0.005
R9496 GND.n8128 GND.n8124 0.005
R9497 GND.n8485 GND.n8484 0.005
R9498 GND.n8479 GND.n8475 0.005
R9499 GND.n439 GND.n438 0.005
R9500 GND.n445 GND.n440 0.005
R9501 GND.n8670 GND.n8669 0.005
R9502 GND.n8664 GND.n8660 0.005
R9503 GND.n390 GND.n389 0.005
R9504 GND.n396 GND.n391 0.005
R9505 GND.n8855 GND.n8854 0.005
R9506 GND.n8849 GND.n8845 0.005
R9507 GND.n341 GND.n340 0.005
R9508 GND.n347 GND.n342 0.005
R9509 GND.n9040 GND.n9039 0.005
R9510 GND.n9034 GND.n9030 0.005
R9511 GND.n292 GND.n291 0.005
R9512 GND.n298 GND.n293 0.005
R9513 GND.n9225 GND.n9224 0.005
R9514 GND.n9219 GND.n9215 0.005
R9515 GND.n243 GND.n242 0.005
R9516 GND.n249 GND.n244 0.005
R9517 GND.n177 GND.n176 0.005
R9518 GND.n9259 GND.n178 0.005
R9519 GND.n182 GND.n181 0.005
R9520 GND.n184 GND.n183 0.005
R9521 GND.n2228 GND.n2227 0.005
R9522 GND.n435 GND.n427 0.005
R9523 GND.n386 GND.n378 0.005
R9524 GND.n337 GND.n329 0.005
R9525 GND.n288 GND.n280 0.005
R9526 GND.n239 GND.n231 0.005
R9527 GND.n180 GND.n179 0.005
R9528 GND.n7865 GND.n7864 0.005
R9529 GND.n7638 GND.n7637 0.005
R9530 GND.n7411 GND.n7410 0.005
R9531 GND.n7184 GND.n7183 0.005
R9532 GND.n6957 GND.n6956 0.005
R9533 GND.n6730 GND.n6729 0.005
R9534 GND.n6410 GND.n6409 0.005
R9535 GND.n7866 GND.n7865 0.004
R9536 GND.n7639 GND.n7638 0.004
R9537 GND.n7412 GND.n7411 0.004
R9538 GND.n7185 GND.n7184 0.004
R9539 GND.n6958 GND.n6957 0.004
R9540 GND.n6731 GND.n6730 0.004
R9541 GND.n6411 GND.n6410 0.004
R9542 GND.n6598 GND.n6597 0.004
R9543 GND.n6615 GND.n6614 0.004
R9544 GND.n6632 GND.n6631 0.004
R9545 GND.n6649 GND.n6648 0.004
R9546 GND.n6666 GND.n6665 0.004
R9547 GND.n6683 GND.n6682 0.004
R9548 GND.n7983 GND.n7982 0.004
R9549 GND.n7981 GND.n7979 0.004
R9550 GND.n8009 GND.n8006 0.004
R9551 GND.n7856 GND.n7855 0.004
R9552 GND.n7884 GND.n7877 0.004
R9553 GND.n7991 GND.n7987 0.004
R9554 GND.n8003 GND.n8002 0.004
R9555 GND.n7894 GND.n7893 0.004
R9556 GND.n7868 GND.n7867 0.004
R9557 GND.n7957 GND.n7956 0.004
R9558 GND.n7965 GND.n7958 0.004
R9559 GND.n8013 GND.n8004 0.004
R9560 GND.n8015 GND.n8014 0.004
R9561 GND.n7905 GND.n7904 0.004
R9562 GND.n7903 GND.n7902 0.004
R9563 GND.n7864 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/SOURCE 0.004
R9564 GND.n6602 GND.n6601 0.004
R9565 GND.n8032 GND.n7839 0.004
R9566 GND.n8046 GND.n8045 0.004
R9567 GND.n8047 GND.n8046 0.004
R9568 GND.n8055 GND.n8054 0.004
R9569 GND.n8053 GND.n8052 0.004
R9570 GND.n6611 GND.n6596 0.004
R9571 GND.n6611 GND.n6610 0.004
R9572 GND.n8056 GND.n8041 0.004
R9573 GND.n8056 GND.n8044 0.004
R9574 GND.n8043 GND.n8042 0.004
R9575 GND.n7756 GND.n7755 0.004
R9576 GND.n7754 GND.n7752 0.004
R9577 GND.n7782 GND.n7779 0.004
R9578 GND.n7629 GND.n7628 0.004
R9579 GND.n7657 GND.n7650 0.004
R9580 GND.n7764 GND.n7760 0.004
R9581 GND.n7776 GND.n7775 0.004
R9582 GND.n7667 GND.n7666 0.004
R9583 GND.n7641 GND.n7640 0.004
R9584 GND.n7730 GND.n7729 0.004
R9585 GND.n7738 GND.n7731 0.004
R9586 GND.n7786 GND.n7777 0.004
R9587 GND.n7788 GND.n7787 0.004
R9588 GND.n7678 GND.n7677 0.004
R9589 GND.n7676 GND.n7675 0.004
R9590 GND.n7637 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/SOURCE 0.004
R9591 GND.n6619 GND.n6618 0.004
R9592 GND.n7805 GND.n7612 0.004
R9593 GND.n7819 GND.n7818 0.004
R9594 GND.n7820 GND.n7819 0.004
R9595 GND.n7828 GND.n7827 0.004
R9596 GND.n7826 GND.n7825 0.004
R9597 GND.n6628 GND.n6613 0.004
R9598 GND.n6628 GND.n6627 0.004
R9599 GND.n7829 GND.n7814 0.004
R9600 GND.n7829 GND.n7817 0.004
R9601 GND.n7816 GND.n7815 0.004
R9602 GND.n7529 GND.n7528 0.004
R9603 GND.n7527 GND.n7525 0.004
R9604 GND.n7555 GND.n7552 0.004
R9605 GND.n7402 GND.n7401 0.004
R9606 GND.n7430 GND.n7423 0.004
R9607 GND.n7537 GND.n7533 0.004
R9608 GND.n7549 GND.n7548 0.004
R9609 GND.n7440 GND.n7439 0.004
R9610 GND.n7414 GND.n7413 0.004
R9611 GND.n7503 GND.n7502 0.004
R9612 GND.n7511 GND.n7504 0.004
R9613 GND.n7559 GND.n7550 0.004
R9614 GND.n7561 GND.n7560 0.004
R9615 GND.n7451 GND.n7450 0.004
R9616 GND.n7449 GND.n7448 0.004
R9617 GND.n7410 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/SOURCE 0.004
R9618 GND.n6636 GND.n6635 0.004
R9619 GND.n7578 GND.n7385 0.004
R9620 GND.n7592 GND.n7591 0.004
R9621 GND.n7593 GND.n7592 0.004
R9622 GND.n7601 GND.n7600 0.004
R9623 GND.n7599 GND.n7598 0.004
R9624 GND.n6645 GND.n6630 0.004
R9625 GND.n6645 GND.n6644 0.004
R9626 GND.n7602 GND.n7587 0.004
R9627 GND.n7602 GND.n7590 0.004
R9628 GND.n7589 GND.n7588 0.004
R9629 GND.n7302 GND.n7301 0.004
R9630 GND.n7300 GND.n7298 0.004
R9631 GND.n7328 GND.n7325 0.004
R9632 GND.n7175 GND.n7174 0.004
R9633 GND.n7203 GND.n7196 0.004
R9634 GND.n7310 GND.n7306 0.004
R9635 GND.n7322 GND.n7321 0.004
R9636 GND.n7213 GND.n7212 0.004
R9637 GND.n7187 GND.n7186 0.004
R9638 GND.n7276 GND.n7275 0.004
R9639 GND.n7284 GND.n7277 0.004
R9640 GND.n7332 GND.n7323 0.004
R9641 GND.n7334 GND.n7333 0.004
R9642 GND.n7224 GND.n7223 0.004
R9643 GND.n7222 GND.n7221 0.004
R9644 GND.n7183 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/SOURCE 0.004
R9645 GND.n6653 GND.n6652 0.004
R9646 GND.n7351 GND.n7158 0.004
R9647 GND.n7365 GND.n7364 0.004
R9648 GND.n7366 GND.n7365 0.004
R9649 GND.n7374 GND.n7373 0.004
R9650 GND.n7372 GND.n7371 0.004
R9651 GND.n6662 GND.n6647 0.004
R9652 GND.n6662 GND.n6661 0.004
R9653 GND.n7375 GND.n7360 0.004
R9654 GND.n7375 GND.n7363 0.004
R9655 GND.n7362 GND.n7361 0.004
R9656 GND.n7075 GND.n7074 0.004
R9657 GND.n7073 GND.n7071 0.004
R9658 GND.n7101 GND.n7098 0.004
R9659 GND.n6948 GND.n6947 0.004
R9660 GND.n6976 GND.n6969 0.004
R9661 GND.n7083 GND.n7079 0.004
R9662 GND.n7095 GND.n7094 0.004
R9663 GND.n6986 GND.n6985 0.004
R9664 GND.n6960 GND.n6959 0.004
R9665 GND.n7049 GND.n7048 0.004
R9666 GND.n7057 GND.n7050 0.004
R9667 GND.n7105 GND.n7096 0.004
R9668 GND.n7107 GND.n7106 0.004
R9669 GND.n6997 GND.n6996 0.004
R9670 GND.n6995 GND.n6994 0.004
R9671 GND.n6956 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/SOURCE 0.004
R9672 GND.n6670 GND.n6669 0.004
R9673 GND.n7124 GND.n6931 0.004
R9674 GND.n7138 GND.n7137 0.004
R9675 GND.n7139 GND.n7138 0.004
R9676 GND.n7147 GND.n7146 0.004
R9677 GND.n7145 GND.n7144 0.004
R9678 GND.n6679 GND.n6664 0.004
R9679 GND.n6679 GND.n6678 0.004
R9680 GND.n7148 GND.n7133 0.004
R9681 GND.n7148 GND.n7136 0.004
R9682 GND.n7135 GND.n7134 0.004
R9683 GND.n6848 GND.n6847 0.004
R9684 GND.n6846 GND.n6844 0.004
R9685 GND.n6874 GND.n6871 0.004
R9686 GND.n6721 GND.n6720 0.004
R9687 GND.n6749 GND.n6742 0.004
R9688 GND.n6856 GND.n6852 0.004
R9689 GND.n6868 GND.n6867 0.004
R9690 GND.n6759 GND.n6758 0.004
R9691 GND.n6733 GND.n6732 0.004
R9692 GND.n6822 GND.n6821 0.004
R9693 GND.n6830 GND.n6823 0.004
R9694 GND.n6878 GND.n6869 0.004
R9695 GND.n6880 GND.n6879 0.004
R9696 GND.n6770 GND.n6769 0.004
R9697 GND.n6768 GND.n6767 0.004
R9698 GND.n6729 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/SOURCE 0.004
R9699 GND.n6687 GND.n6686 0.004
R9700 GND.n6897 GND.n6704 0.004
R9701 GND.n6911 GND.n6910 0.004
R9702 GND.n6912 GND.n6911 0.004
R9703 GND.n6920 GND.n6919 0.004
R9704 GND.n6918 GND.n6917 0.004
R9705 GND.n6696 GND.n6681 0.004
R9706 GND.n6696 GND.n6695 0.004
R9707 GND.n6921 GND.n6906 0.004
R9708 GND.n6921 GND.n6909 0.004
R9709 GND.n6908 GND.n6907 0.004
R9710 GND.n6516 GND.n6515 0.004
R9711 GND.n6514 GND.n6512 0.004
R9712 GND.n6542 GND.n6539 0.004
R9713 GND.n6437 GND.n6436 0.004
R9714 GND.n6429 GND.n6422 0.004
R9715 GND.n6524 GND.n6520 0.004
R9716 GND.n6536 GND.n6535 0.004
R9717 GND.n6401 GND.n6400 0.004
R9718 GND.n6413 GND.n6412 0.004
R9719 GND.n6490 GND.n6489 0.004
R9720 GND.n6498 GND.n6491 0.004
R9721 GND.n6546 GND.n6537 0.004
R9722 GND.n6548 GND.n6547 0.004
R9723 GND.n6449 GND.n6448 0.004
R9724 GND.n6447 GND.n6446 0.004
R9725 GND.n6409 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/SOURCE 0.004
R9726 GND.n6581 GND.n6580 0.004
R9727 GND.n6576 GND.n6575 0.004
R9728 GND.n6574 GND.n6573 0.004
R9729 GND.n591 GND.n590 0.004
R9730 GND.n554 GND.n552 0.004
R9731 GND.n558 GND.n556 0.004
R9732 GND.n1001 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13/DRAIN 0.004
R9733 GND.n1039 GND.n1037 0.004
R9734 GND.n1044 GND.n1041 0.004
R9735 GND.n6061 GND.n6060 0.004
R9736 GND.n869 GND.n867 0.004
R9737 GND.n873 GND.n871 0.004
R9738 GND.n6023 GND.n6021 0.004
R9739 GND.n6027 GND.n6025 0.004
R9740 GND.n1286 GND.n1283 0.004
R9741 GND.n2623 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14/DRAIN 0.004
R9742 GND.n2661 GND.n2659 0.004
R9743 GND.n2666 GND.n2663 0.004
R9744 GND.n3889 GND.n3888 0.004
R9745 GND.n2491 GND.n2489 0.004
R9746 GND.n2495 GND.n2493 0.004
R9747 GND.n3851 GND.n3849 0.004
R9748 GND.n3855 GND.n3853 0.004
R9749 GND.n2357 GND.n2356 0.004
R9750 GND.n2320 GND.n2318 0.004
R9751 GND.n2324 GND.n2322 0.004
R9752 GND.n3990 GND.n3989 0.004
R9753 GND.n4010 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15/SOURCE 0.004
R9754 GND.n2945 GND.n2943 0.004
R9755 GND.n2941 GND.n2939 0.004
R9756 GND.n4056 GND.n4054 0.004
R9757 GND.n4052 GND.n4050 0.004
R9758 GND.n6286 GND.n6285 0.004
R9759 GND.n6306 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16/SOURCE 0.004
R9760 GND.n1519 GND.n1517 0.004
R9761 GND.n1515 GND.n1513 0.004
R9762 GND.n6240 GND.n6238 0.004
R9763 GND.n6245 GND.n6242 0.004
R9764 GND.n6327 GND.n6326 0.004
R9765 GND.n8229 GND.n8226 0.004
R9766 GND.n8240 GND.n8237 0.004
R9767 GND.n8288 GND.n8263 0.004
R9768 GND.n8287 GND.n8285 0.004
R9769 GND.n8157 GND.n8154 0.004
R9770 GND.n8168 GND.n8165 0.004
R9771 GND.n8216 GND.n8191 0.004
R9772 GND.n8214 GND.n8212 0.004
R9773 GND.n8100 GND.n8099 0.004
R9774 GND.n8107 GND.n8106 0.004
R9775 GND.n8301 GND.n8299 0.004
R9776 GND.n8301 GND.n8300 0.004
R9777 GND.n8138 GND.n8137 0.004
R9778 GND.n8098 GND.n8090 0.004
R9779 GND.n8113 GND.n8112 0.004
R9780 GND.n8132 GND.n8131 0.004
R9781 GND.n8336 GND.n8333 0.004
R9782 GND.n8347 GND.n8344 0.004
R9783 GND.n8395 GND.n8370 0.004
R9784 GND.n8394 GND.n8392 0.004
R9785 GND.n8408 GND.n8405 0.004
R9786 GND.n8419 GND.n8416 0.004
R9787 GND.n8467 GND.n8442 0.004
R9788 GND.n8465 GND.n8463 0.004
R9789 GND.n437 GND.n436 0.004
R9790 GND.n443 GND.n442 0.004
R9791 GND.n414 GND.n412 0.004
R9792 GND.n414 GND.n413 0.004
R9793 GND.n8473 GND.n8471 0.004
R9794 GND.n8486 GND.n8485 0.004
R9795 GND.n440 GND.n439 0.004
R9796 GND.n450 GND.n449 0.004
R9797 GND.n407 GND.n406 0.004
R9798 GND.n8483 GND.n8482 0.004
R9799 GND.n8481 GND.n8480 0.004
R9800 GND.n451 GND.n426 0.004
R9801 GND.n424 GND.n405 0.004
R9802 GND.n424 GND.n423 0.004
R9803 GND.n8491 GND.n8320 0.004
R9804 GND.n8491 GND.n8322 0.004
R9805 GND.n8521 GND.n8518 0.004
R9806 GND.n8532 GND.n8529 0.004
R9807 GND.n8580 GND.n8555 0.004
R9808 GND.n8579 GND.n8577 0.004
R9809 GND.n8593 GND.n8590 0.004
R9810 GND.n8604 GND.n8601 0.004
R9811 GND.n8652 GND.n8627 0.004
R9812 GND.n8650 GND.n8648 0.004
R9813 GND.n388 GND.n387 0.004
R9814 GND.n394 GND.n393 0.004
R9815 GND.n365 GND.n363 0.004
R9816 GND.n365 GND.n364 0.004
R9817 GND.n8658 GND.n8656 0.004
R9818 GND.n8671 GND.n8670 0.004
R9819 GND.n391 GND.n390 0.004
R9820 GND.n401 GND.n400 0.004
R9821 GND.n358 GND.n357 0.004
R9822 GND.n8668 GND.n8667 0.004
R9823 GND.n8666 GND.n8665 0.004
R9824 GND.n402 GND.n377 0.004
R9825 GND.n375 GND.n356 0.004
R9826 GND.n375 GND.n374 0.004
R9827 GND.n8676 GND.n8505 0.004
R9828 GND.n8676 GND.n8507 0.004
R9829 GND.n8706 GND.n8703 0.004
R9830 GND.n8717 GND.n8714 0.004
R9831 GND.n8765 GND.n8740 0.004
R9832 GND.n8764 GND.n8762 0.004
R9833 GND.n8778 GND.n8775 0.004
R9834 GND.n8789 GND.n8786 0.004
R9835 GND.n8837 GND.n8812 0.004
R9836 GND.n8835 GND.n8833 0.004
R9837 GND.n339 GND.n338 0.004
R9838 GND.n345 GND.n344 0.004
R9839 GND.n316 GND.n314 0.004
R9840 GND.n316 GND.n315 0.004
R9841 GND.n8843 GND.n8841 0.004
R9842 GND.n8856 GND.n8855 0.004
R9843 GND.n342 GND.n341 0.004
R9844 GND.n352 GND.n351 0.004
R9845 GND.n309 GND.n308 0.004
R9846 GND.n8853 GND.n8852 0.004
R9847 GND.n8851 GND.n8850 0.004
R9848 GND.n353 GND.n328 0.004
R9849 GND.n326 GND.n307 0.004
R9850 GND.n326 GND.n325 0.004
R9851 GND.n8861 GND.n8690 0.004
R9852 GND.n8861 GND.n8692 0.004
R9853 GND.n8891 GND.n8888 0.004
R9854 GND.n8902 GND.n8899 0.004
R9855 GND.n8950 GND.n8925 0.004
R9856 GND.n8949 GND.n8947 0.004
R9857 GND.n8963 GND.n8960 0.004
R9858 GND.n8974 GND.n8971 0.004
R9859 GND.n9022 GND.n8997 0.004
R9860 GND.n9020 GND.n9018 0.004
R9861 GND.n290 GND.n289 0.004
R9862 GND.n296 GND.n295 0.004
R9863 GND.n267 GND.n265 0.004
R9864 GND.n267 GND.n266 0.004
R9865 GND.n9028 GND.n9026 0.004
R9866 GND.n9041 GND.n9040 0.004
R9867 GND.n293 GND.n292 0.004
R9868 GND.n303 GND.n302 0.004
R9869 GND.n260 GND.n259 0.004
R9870 GND.n9038 GND.n9037 0.004
R9871 GND.n9036 GND.n9035 0.004
R9872 GND.n304 GND.n279 0.004
R9873 GND.n277 GND.n258 0.004
R9874 GND.n277 GND.n276 0.004
R9875 GND.n9046 GND.n8875 0.004
R9876 GND.n9046 GND.n8877 0.004
R9877 GND.n9076 GND.n9073 0.004
R9878 GND.n9087 GND.n9084 0.004
R9879 GND.n9135 GND.n9110 0.004
R9880 GND.n9134 GND.n9132 0.004
R9881 GND.n9148 GND.n9145 0.004
R9882 GND.n9159 GND.n9156 0.004
R9883 GND.n9207 GND.n9182 0.004
R9884 GND.n9205 GND.n9203 0.004
R9885 GND.n241 GND.n240 0.004
R9886 GND.n247 GND.n246 0.004
R9887 GND.n218 GND.n216 0.004
R9888 GND.n218 GND.n217 0.004
R9889 GND.n9213 GND.n9211 0.004
R9890 GND.n9226 GND.n9225 0.004
R9891 GND.n244 GND.n243 0.004
R9892 GND.n254 GND.n253 0.004
R9893 GND.n211 GND.n210 0.004
R9894 GND.n9223 GND.n9222 0.004
R9895 GND.n9221 GND.n9220 0.004
R9896 GND.n255 GND.n230 0.004
R9897 GND.n228 GND.n209 0.004
R9898 GND.n228 GND.n227 0.004
R9899 GND.n9231 GND.n9060 0.004
R9900 GND.n9231 GND.n9062 0.004
R9901 GND.n37 GND.n34 0.004
R9902 GND.n48 GND.n45 0.004
R9903 GND.n96 GND.n71 0.004
R9904 GND.n95 GND.n93 0.004
R9905 GND.n109 GND.n106 0.004
R9906 GND.n120 GND.n117 0.004
R9907 GND.n168 GND.n143 0.004
R9908 GND.n166 GND.n164 0.004
R9909 GND.n8 GND.n7 0.004
R9910 GND.n11 GND.n10 0.004
R9911 GND.n20 GND.n19 0.004
R9912 GND.n21 GND.n20 0.004
R9913 GND.n171 GND.n170 0.004
R9914 GND.n176 GND.n175 0.004
R9915 GND.n183 GND.n182 0.004
R9916 GND.n186 GND.n185 0.004
R9917 GND.n188 GND.n187 0.004
R9918 GND.n194 GND.n193 0.004
R9919 GND.n9255 GND.n9254 0.004
R9920 GND.n9258 GND.n9256 0.004
R9921 GND.n199 GND.n198 0.004
R9922 GND.n200 GND.n199 0.004
R9923 GND.n203 GND.n202 0.004
R9924 GND.n204 GND.n203 0.004
R9925 GND.n9251 GND.n206 0.004
R9926 GND.n9251 GND.n9250 0.004
R9927 GND.n8480 GND.n8474 0.004
R9928 GND.n8665 GND.n8659 0.004
R9929 GND.n8850 GND.n8844 0.004
R9930 GND.n9035 GND.n9029 0.004
R9931 GND.n9220 GND.n9214 0.004
R9932 GND.n9258 GND.n9257 0.004
R9933 GND.n6341 GND.n6340 0.004
R9934 GND.n7936 GND.n7935 0.003
R9935 GND.n7956 GND.n7946 0.003
R9936 GND.n7958 GND.n7957 0.003
R9937 GND.n7918 GND.n7907 0.003
R9938 GND.n7890 GND.n7889 0.003
R9939 GND.n7889 GND.n7888 0.003
R9940 GND.n7888 GND.n7887 0.003
R9941 GND.n6606 GND.n6605 0.003
R9942 GND.n8052 GND.n8051 0.003
R9943 GND.n7709 GND.n7708 0.003
R9944 GND.n7729 GND.n7719 0.003
R9945 GND.n7731 GND.n7730 0.003
R9946 GND.n7691 GND.n7680 0.003
R9947 GND.n7663 GND.n7662 0.003
R9948 GND.n7662 GND.n7661 0.003
R9949 GND.n7661 GND.n7660 0.003
R9950 GND.n6623 GND.n6622 0.003
R9951 GND.n7825 GND.n7824 0.003
R9952 GND.n7482 GND.n7481 0.003
R9953 GND.n7502 GND.n7492 0.003
R9954 GND.n7504 GND.n7503 0.003
R9955 GND.n7464 GND.n7453 0.003
R9956 GND.n7436 GND.n7435 0.003
R9957 GND.n7435 GND.n7434 0.003
R9958 GND.n7434 GND.n7433 0.003
R9959 GND.n6640 GND.n6639 0.003
R9960 GND.n7598 GND.n7597 0.003
R9961 GND.n7255 GND.n7254 0.003
R9962 GND.n7275 GND.n7265 0.003
R9963 GND.n7277 GND.n7276 0.003
R9964 GND.n7237 GND.n7226 0.003
R9965 GND.n7209 GND.n7208 0.003
R9966 GND.n7208 GND.n7207 0.003
R9967 GND.n7207 GND.n7206 0.003
R9968 GND.n6657 GND.n6656 0.003
R9969 GND.n7371 GND.n7370 0.003
R9970 GND.n7028 GND.n7027 0.003
R9971 GND.n7048 GND.n7038 0.003
R9972 GND.n7050 GND.n7049 0.003
R9973 GND.n7010 GND.n6999 0.003
R9974 GND.n6982 GND.n6981 0.003
R9975 GND.n6981 GND.n6980 0.003
R9976 GND.n6980 GND.n6979 0.003
R9977 GND.n6674 GND.n6673 0.003
R9978 GND.n7144 GND.n7143 0.003
R9979 GND.n6801 GND.n6800 0.003
R9980 GND.n6821 GND.n6811 0.003
R9981 GND.n6823 GND.n6822 0.003
R9982 GND.n6783 GND.n6772 0.003
R9983 GND.n6755 GND.n6754 0.003
R9984 GND.n6754 GND.n6753 0.003
R9985 GND.n6753 GND.n6752 0.003
R9986 GND.n6691 GND.n6690 0.003
R9987 GND.n6917 GND.n6916 0.003
R9988 GND.n6469 GND.n6468 0.003
R9989 GND.n6489 GND.n6479 0.003
R9990 GND.n6491 GND.n6490 0.003
R9991 GND.n6462 GND.n6451 0.003
R9992 GND.n6445 GND.n6434 0.003
R9993 GND.n6434 GND.n6433 0.003
R9994 GND.n6433 GND.n6432 0.003
R9995 GND.n6364 GND.n6363 0.003
R9996 GND.n6585 GND.n6584 0.003
R9997 GND.n6570 GND.n6569 0.003
R9998 GND.n585 GND.n584 0.003
R9999 GND.n1016 GND.n1015 0.003
R10000 GND.n6055 GND.n6054 0.003
R10001 GND.n6128 GND.n6124 0.003
R10002 GND.n6137 GND.n6135 0.003
R10003 GND.n2638 GND.n2637 0.003
R10004 GND.n3883 GND.n3882 0.003
R10005 GND.n3956 GND.n3952 0.003
R10006 GND.n3965 GND.n3963 0.003
R10007 GND.n2351 GND.n2350 0.003
R10008 GND.n3997 GND.n3996 0.003
R10009 GND.n2263 GND.n2259 0.003
R10010 GND.n2269 GND.n2265 0.003
R10011 GND.n6293 GND.n6292 0.003
R10012 GND.n497 GND.n493 0.003
R10013 GND.n503 GND.n499 0.003
R10014 GND.n8295 GND.n8294 0.003
R10015 GND.n8121 GND.n8116 0.003
R10016 GND.n8141 GND.n8135 0.003
R10017 GND.n417 GND.n416 0.003
R10018 GND.n411 GND.n407 0.003
R10019 GND.n8489 GND.n8483 0.003
R10020 GND.n368 GND.n367 0.003
R10021 GND.n362 GND.n358 0.003
R10022 GND.n8674 GND.n8668 0.003
R10023 GND.n319 GND.n318 0.003
R10024 GND.n313 GND.n309 0.003
R10025 GND.n8859 GND.n8853 0.003
R10026 GND.n270 GND.n269 0.003
R10027 GND.n264 GND.n260 0.003
R10028 GND.n9044 GND.n9038 0.003
R10029 GND.n221 GND.n220 0.003
R10030 GND.n215 GND.n211 0.003
R10031 GND.n9229 GND.n9223 0.003
R10032 GND.n24 GND.n23 0.003
R10033 GND.n189 GND.n188 0.003
R10034 GND.n9254 GND.n9253 0.003
R10035 GND.n459 GND.n458 0.003
R10036 GND.n8069 GND.n8068 0.003
R10037 GND.n6370 GND.n6369 0.002
R10038 GND.n6583 GND.n6582 0.002
R10039 GND.n6577 GND.n6576 0.002
R10040 GND.n6571 GND.n6570 0.002
R10041 GND.n8104 GND.n8103 0.002
R10042 GND.n8116 GND.n8115 0.002
R10043 GND.n8292 GND.n8291 0.002
R10044 GND.n8134 GND.n8133 0.002
R10045 GND.n8103 GND.n8102 0.002
R10046 GND.n8293 GND.n8292 0.002
R10047 GND.n8115 GND.n8114 0.002
R10048 GND.n8135 GND.n8134 0.002
R10049 GND.n6369 GND.n6368 0.002
R10050 GND.n6572 GND.n6571 0.002
R10051 GND.n6584 GND.n6583 0.002
R10052 GND.n6578 GND.n6577 0.002
R10053 GND.n8079 GND.n8078 0.002
R10054 GND.n8082 GND.n8081 0.002
R10055 GND.n8087 GND.n8086 0.002
R10056 GND.n8085 GND.n8084 0.002
R10057 GND.n6591 GND.n6590 0.002
R10058 GND.n6594 GND.n6593 0.002
R10059 GND.n8031 GND.n7934 0.002
R10060 GND.n7804 GND.n7707 0.002
R10061 GND.n7577 GND.n7480 0.002
R10062 GND.n7350 GND.n7253 0.002
R10063 GND.n7123 GND.n7026 0.002
R10064 GND.n6896 GND.n6799 0.002
R10065 GND.n6564 GND.n6467 0.002
R10066 GND.n8304 GND.n8303 0.002
R10067 GND.n8305 GND.n8304 0.002
R10068 GND.n7873 GND.n7871 0.002
R10069 GND.n7972 GND.n7965 0.002
R10070 GND.n7907 GND.n7906 0.002
R10071 GND.n7876 GND.n7866 0.002
R10072 GND.n6600 GND.n6599 0.002
R10073 GND.n6601 GND.n6600 0.002
R10074 GND.n6604 GND.n6603 0.002
R10075 GND.n6607 GND.n6604 0.002
R10076 GND.n6607 GND.n6606 0.002
R10077 GND.n8051 GND.n8050 0.002
R10078 GND.n8049 GND.n8048 0.002
R10079 GND.n6596 GND.n6595 0.002
R10080 GND.n8044 GND.n8043 0.002
R10081 GND.n7646 GND.n7644 0.002
R10082 GND.n7745 GND.n7738 0.002
R10083 GND.n7680 GND.n7679 0.002
R10084 GND.n7649 GND.n7639 0.002
R10085 GND.n6617 GND.n6616 0.002
R10086 GND.n6618 GND.n6617 0.002
R10087 GND.n6621 GND.n6620 0.002
R10088 GND.n6624 GND.n6621 0.002
R10089 GND.n6624 GND.n6623 0.002
R10090 GND.n7824 GND.n7823 0.002
R10091 GND.n7822 GND.n7821 0.002
R10092 GND.n6613 GND.n6612 0.002
R10093 GND.n7817 GND.n7816 0.002
R10094 GND.n7419 GND.n7417 0.002
R10095 GND.n7518 GND.n7511 0.002
R10096 GND.n7453 GND.n7452 0.002
R10097 GND.n7422 GND.n7412 0.002
R10098 GND.n6634 GND.n6633 0.002
R10099 GND.n6635 GND.n6634 0.002
R10100 GND.n6638 GND.n6637 0.002
R10101 GND.n6641 GND.n6638 0.002
R10102 GND.n6641 GND.n6640 0.002
R10103 GND.n7597 GND.n7596 0.002
R10104 GND.n7595 GND.n7594 0.002
R10105 GND.n6630 GND.n6629 0.002
R10106 GND.n7590 GND.n7589 0.002
R10107 GND.n7192 GND.n7190 0.002
R10108 GND.n7291 GND.n7284 0.002
R10109 GND.n7226 GND.n7225 0.002
R10110 GND.n7195 GND.n7185 0.002
R10111 GND.n6651 GND.n6650 0.002
R10112 GND.n6652 GND.n6651 0.002
R10113 GND.n6655 GND.n6654 0.002
R10114 GND.n6658 GND.n6655 0.002
R10115 GND.n6658 GND.n6657 0.002
R10116 GND.n7370 GND.n7369 0.002
R10117 GND.n7368 GND.n7367 0.002
R10118 GND.n6647 GND.n6646 0.002
R10119 GND.n7363 GND.n7362 0.002
R10120 GND.n6965 GND.n6963 0.002
R10121 GND.n7064 GND.n7057 0.002
R10122 GND.n6999 GND.n6998 0.002
R10123 GND.n6968 GND.n6958 0.002
R10124 GND.n6668 GND.n6667 0.002
R10125 GND.n6669 GND.n6668 0.002
R10126 GND.n6672 GND.n6671 0.002
R10127 GND.n6675 GND.n6672 0.002
R10128 GND.n6675 GND.n6674 0.002
R10129 GND.n7143 GND.n7142 0.002
R10130 GND.n7141 GND.n7140 0.002
R10131 GND.n6664 GND.n6663 0.002
R10132 GND.n7136 GND.n7135 0.002
R10133 GND.n6738 GND.n6736 0.002
R10134 GND.n6837 GND.n6830 0.002
R10135 GND.n6772 GND.n6771 0.002
R10136 GND.n6741 GND.n6731 0.002
R10137 GND.n6685 GND.n6684 0.002
R10138 GND.n6686 GND.n6685 0.002
R10139 GND.n6689 GND.n6688 0.002
R10140 GND.n6692 GND.n6689 0.002
R10141 GND.n6692 GND.n6691 0.002
R10142 GND.n6916 GND.n6915 0.002
R10143 GND.n6914 GND.n6913 0.002
R10144 GND.n6681 GND.n6680 0.002
R10145 GND.n6909 GND.n6908 0.002
R10146 GND.n6419 GND.n6417 0.002
R10147 GND.n6505 GND.n6498 0.002
R10148 GND.n6451 GND.n6450 0.002
R10149 GND.n6421 GND.n6411 0.002
R10150 GND.n6365 GND.n6364 0.002
R10151 GND.n6367 GND.n6366 0.002
R10152 GND.n6368 GND.n6367 0.002
R10153 GND.n6372 GND.n6371 0.002
R10154 GND.n6586 GND.n6372 0.002
R10155 GND.n6586 GND.n6585 0.002
R10156 GND.n6569 GND.n6568 0.002
R10157 GND.n6567 GND.n6566 0.002
R10158 GND.n6566 GND.n6565 0.002
R10159 GND.n576 GND.n575 0.002
R10160 GND.n520 GND.n519 0.002
R10161 GND.n602 GND.n600 0.002
R10162 GND.n607 GND.n605 0.002
R10163 GND.n1696 GND.n1694 0.002
R10164 GND.n1686 GND.n1678 0.002
R10165 GND.n1378 GND.n1370 0.002
R10166 GND.n1388 GND.n1386 0.002
R10167 GND.n1191 GND.n1189 0.002
R10168 GND.n1181 GND.n1173 0.002
R10169 GND.n744 GND.n736 0.002
R10170 GND.n754 GND.n752 0.002
R10171 GND.n2806 GND.n2798 0.002
R10172 GND.n2816 GND.n2814 0.002
R10173 GND.n3119 GND.n3117 0.002
R10174 GND.n3109 GND.n3101 0.002
R10175 GND.n3709 GND.n3707 0.002
R10176 GND.n3699 GND.n3691 0.002
R10177 GND.n1007 GND.n1006 0.002
R10178 GND.n992 GND.n990 0.002
R10179 GND.n997 GND.n995 0.002
R10180 GND.n1077 GND.n1074 0.002
R10181 GND.n6046 GND.n6045 0.002
R10182 GND.n835 GND.n834 0.002
R10183 GND.n895 GND.n893 0.002
R10184 GND.n900 GND.n898 0.002
R10185 GND.n5989 GND.n5988 0.002
R10186 GND.n6072 GND.n6070 0.002
R10187 GND.n6077 GND.n6075 0.002
R10188 GND.n1277 GND.n1274 0.002
R10189 GND.n1265 GND.n1089 0.002
R10190 GND.n2629 GND.n2628 0.002
R10191 GND.n2614 GND.n2612 0.002
R10192 GND.n2619 GND.n2617 0.002
R10193 GND.n2699 GND.n2696 0.002
R10194 GND.n3874 GND.n3873 0.002
R10195 GND.n2457 GND.n2456 0.002
R10196 GND.n2517 GND.n2515 0.002
R10197 GND.n2522 GND.n2520 0.002
R10198 GND.n3817 GND.n3816 0.002
R10199 GND.n3900 GND.n3898 0.002
R10200 GND.n3905 GND.n3903 0.002
R10201 GND.n1922 GND.n1914 0.002
R10202 GND.n1932 GND.n1930 0.002
R10203 GND.n2102 GND.n2094 0.002
R10204 GND.n2112 GND.n2110 0.002
R10205 GND.n2205 GND.n2204 0.002
R10206 GND.n2206 GND.n2205 0.002
R10207 GND.n4350 GND.n2206 0.002
R10208 GND.n4351 GND.n4350 0.002
R10209 GND.n4354 GND.n4351 0.002
R10210 GND.n4354 GND.n4353 0.002
R10211 GND.n4368 GND.n4367 0.002
R10212 GND.n4383 GND.n4369 0.002
R10213 GND.n4383 GND.n4382 0.002
R10214 GND.n4382 GND.n4381 0.002
R10215 GND.n4381 GND.n4372 0.002
R10216 GND.n4372 GND.n4371 0.002
R10217 GND.n4371 GND.n4370 0.002
R10218 GND.n2197 GND.n2196 0.002
R10219 GND.n2200 GND.n2199 0.002
R10220 GND.n2201 GND.n2200 0.002
R10221 GND.n4355 GND.n2203 0.002
R10222 GND.n4356 GND.n4355 0.002
R10223 GND.n4387 GND.n4357 0.002
R10224 GND.n4387 GND.n4386 0.002
R10225 GND.n4385 GND.n4384 0.002
R10226 GND.n4384 GND.n4366 0.002
R10227 GND.n4364 GND.n4363 0.002
R10228 GND.n4363 GND.n4362 0.002
R10229 GND.n4360 GND.n4359 0.002
R10230 GND.n5232 GND.n5224 0.002
R10231 GND.n5242 GND.n5240 0.002
R10232 GND.n5412 GND.n5404 0.002
R10233 GND.n5422 GND.n5420 0.002
R10234 GND.n4482 GND.n4474 0.002
R10235 GND.n4492 GND.n4490 0.002
R10236 GND.n4664 GND.n4656 0.002
R10237 GND.n4675 GND.n4673 0.002
R10238 GND.n4853 GND.n4845 0.002
R10239 GND.n4863 GND.n4861 0.002
R10240 GND.n5033 GND.n5025 0.002
R10241 GND.n5043 GND.n5041 0.002
R10242 GND.n3500 GND.n3498 0.002
R10243 GND.n3490 GND.n3481 0.002
R10244 GND.n3316 GND.n3314 0.002
R10245 GND.n3306 GND.n3298 0.002
R10246 GND.n5798 GND.n5796 0.002
R10247 GND.n5788 GND.n5780 0.002
R10248 GND.n5618 GND.n5616 0.002
R10249 GND.n5608 GND.n5600 0.002
R10250 GND.n2218 GND.n2217 0.002
R10251 GND.n2223 GND.n2218 0.002
R10252 GND.n2240 GND.n2231 0.002
R10253 GND.n2241 GND.n2240 0.002
R10254 GND.n2243 GND.n2242 0.002
R10255 GND.n2244 GND.n2243 0.002
R10256 GND.n4317 GND.n2245 0.002
R10257 GND.n4318 GND.n4317 0.002
R10258 GND.n4338 GND.n4318 0.002
R10259 GND.n4338 GND.n4337 0.002
R10260 GND.n4337 GND.n4336 0.002
R10261 GND.n4336 GND.n4326 0.002
R10262 GND.n2222 GND.n2221 0.002
R10263 GND.n2239 GND.n2234 0.002
R10264 GND.n4310 GND.n2247 0.002
R10265 GND.n4311 GND.n4310 0.002
R10266 GND.n4316 GND.n4312 0.002
R10267 GND.n4325 GND.n4321 0.002
R10268 GND.n4325 GND.n4324 0.002
R10269 GND.n2342 GND.n2341 0.002
R10270 GND.n2286 GND.n2285 0.002
R10271 GND.n2368 GND.n2366 0.002
R10272 GND.n2373 GND.n2371 0.002
R10273 GND.n4006 GND.n4005 0.002
R10274 GND.n2966 GND.n2964 0.002
R10275 GND.n2962 GND.n2959 0.002
R10276 GND.n2910 GND.n2909 0.002
R10277 GND.n4077 GND.n4075 0.002
R10278 GND.n4073 GND.n4070 0.002
R10279 GND.n4021 GND.n4020 0.002
R10280 GND.n2896 GND.n2421 0.002
R10281 GND.n4304 GND.n4300 0.002
R10282 GND.n4211 GND.n4203 0.002
R10283 GND.n4221 GND.n4219 0.002
R10284 GND.n6302 GND.n6301 0.002
R10285 GND.n1545 GND.n1543 0.002
R10286 GND.n1541 GND.n1538 0.002
R10287 GND.n1483 GND.n1482 0.002
R10288 GND.n6213 GND.n6211 0.002
R10289 GND.n6218 GND.n6216 0.002
R10290 GND.n6278 GND.n6275 0.002
R10291 GND.n1469 GND.n655 0.002
R10292 GND.n6313 GND.n661 0.002
R10293 GND.n6345 GND.n6342 0.002
R10294 GND.n6346 GND.n6345 0.002
R10295 GND.n6351 GND.n6347 0.002
R10296 GND.n6352 GND.n6351 0.002
R10297 GND.n6358 GND.n6354 0.002
R10298 GND.n474 GND.n467 0.002
R10299 GND.n474 GND.n470 0.002
R10300 GND.n461 GND.n460 0.002
R10301 GND.n482 GND.n481 0.002
R10302 GND.n483 GND.n482 0.002
R10303 GND.n485 GND.n484 0.002
R10304 GND.n486 GND.n485 0.002
R10305 GND.n6359 GND.n486 0.002
R10306 GND.n6360 GND.n6359 0.002
R10307 GND.n475 GND.n464 0.002
R10308 GND.n462 GND.n452 0.002
R10309 GND.n8119 GND.n8118 0.002
R10310 GND.n8302 GND.n8121 0.002
R10311 GND.n8298 GND.n8297 0.002
R10312 GND.n8290 GND.n8143 0.002
R10313 GND.n8142 GND.n8141 0.002
R10314 GND.n409 GND.n408 0.002
R10315 GND.n8479 GND.n8478 0.002
R10316 GND.n421 GND.n411 0.002
R10317 GND.n420 GND.n419 0.002
R10318 GND.n8470 GND.n8469 0.002
R10319 GND.n8490 GND.n8489 0.002
R10320 GND.n426 GND.n425 0.002
R10321 GND.n8322 GND.n8321 0.002
R10322 GND.n360 GND.n359 0.002
R10323 GND.n8664 GND.n8663 0.002
R10324 GND.n372 GND.n362 0.002
R10325 GND.n371 GND.n370 0.002
R10326 GND.n8655 GND.n8654 0.002
R10327 GND.n8675 GND.n8674 0.002
R10328 GND.n377 GND.n376 0.002
R10329 GND.n8507 GND.n8506 0.002
R10330 GND.n311 GND.n310 0.002
R10331 GND.n8849 GND.n8848 0.002
R10332 GND.n323 GND.n313 0.002
R10333 GND.n322 GND.n321 0.002
R10334 GND.n8840 GND.n8839 0.002
R10335 GND.n8860 GND.n8859 0.002
R10336 GND.n328 GND.n327 0.002
R10337 GND.n8692 GND.n8691 0.002
R10338 GND.n262 GND.n261 0.002
R10339 GND.n9034 GND.n9033 0.002
R10340 GND.n274 GND.n264 0.002
R10341 GND.n273 GND.n272 0.002
R10342 GND.n9025 GND.n9024 0.002
R10343 GND.n9045 GND.n9044 0.002
R10344 GND.n279 GND.n278 0.002
R10345 GND.n8877 GND.n8876 0.002
R10346 GND.n213 GND.n212 0.002
R10347 GND.n9219 GND.n9218 0.002
R10348 GND.n225 GND.n215 0.002
R10349 GND.n224 GND.n223 0.002
R10350 GND.n9210 GND.n9209 0.002
R10351 GND.n9230 GND.n9229 0.002
R10352 GND.n230 GND.n229 0.002
R10353 GND.n9062 GND.n9061 0.002
R10354 GND.n7 GND.n6 0.002
R10355 GND.n13 GND.n12 0.002
R10356 GND.n17 GND.n16 0.002
R10357 GND.n19 GND.n18 0.002
R10358 GND.n9260 GND.n9259 0.002
R10359 GND.n190 GND.n189 0.002
R10360 GND.n192 GND.n191 0.002
R10361 GND.n196 GND.n195 0.002
R10362 GND.n9253 GND.n9252 0.002
R10363 GND.n198 GND.n197 0.002
R10364 GND.n9250 GND.n9249 0.002
R10365 GND.n8310 GND.n8309 0.002
R10366 GND.n8309 GND.n8308 0.002
R10367 GND.n8308 GND.n8307 0.002
R10368 GND.n8307 GND.n8077 0.002
R10369 GND.n8077 GND.n8076 0.002
R10370 GND.n8060 GND.n8059 0.002
R10371 GND.n8061 GND.n8060 0.002
R10372 GND.n8065 GND.n8061 0.002
R10373 GND.n8065 GND.n8064 0.002
R10374 GND.n8064 GND.n8063 0.002
R10375 GND.n8063 GND.n8062 0.002
R10376 GND.n2224 GND.n2208 0.002
R10377 GND.n2225 GND.n2224 0.002
R10378 GND.n2226 GND.n2225 0.002
R10379 GND.n2227 GND.n2226 0.002
R10380 GND.n2229 GND.n2228 0.002
R10381 GND.n2230 GND.n2229 0.002
R10382 GND.n4339 GND.n2230 0.002
R10383 GND.n4340 GND.n4339 0.002
R10384 GND.n4341 GND.n4340 0.002
R10385 GND.n4342 GND.n4341 0.002
R10386 GND.n4344 GND.n4343 0.002
R10387 GND.n4345 GND.n4344 0.002
R10388 GND.n4349 GND.n4345 0.002
R10389 GND.n4349 GND.n4348 0.002
R10390 GND.n4348 GND.n4347 0.002
R10391 GND.n4347 GND.n4346 0.002
R10392 GND.n4374 GND.n4373 0.002
R10393 GND.n4375 GND.n4374 0.002
R10394 GND.n4380 GND.n4375 0.002
R10395 GND.n4380 GND.n4379 0.002
R10396 GND.n4379 GND.n4378 0.002
R10397 GND.n4378 GND.n4377 0.002
R10398 GND.n477 GND.n476 0.002
R10399 GND.n8306 GND.n8305 0.002
R10400 GND.n6588 GND.n6587 0.002
R10401 GND.n8072 GND.n8071 0.002
R10402 GND.n2202 GND.n2201 0.002
R10403 GND.n4362 GND.n4361 0.002
R10404 GND.n4366 GND.n4365 0.002
R10405 GND.n2233 GND.n2232 0.002
R10406 GND.n2221 GND.n2220 0.002
R10407 GND.n4324 GND.n4323 0.002
R10408 GND.n4321 GND.n4320 0.002
R10409 GND.n6361 GND.n480 0.002
R10410 GND.n463 GND.n462 0.002
R10411 GND.n8068 GND.n8067 0.001
R10412 GND.n8067 GND.n8066 0.001
R10413 GND.n9247 GND.n9246 0.001
R10414 GND.n9248 GND.n9244 0.001
R10415 GND.n9242 GND.n9240 0.001
R10416 GND.n9238 GND.n9236 0.001
R10417 GND.n9234 GND.n9233 0.001
R10418 GND.n9232 GND.n9059 0.001
R10419 GND.n9058 GND.n9057 0.001
R10420 GND.n9056 GND.n9055 0.001
R10421 GND.n9054 GND.n9053 0.001
R10422 GND.n9052 GND.n9051 0.001
R10423 GND.n9049 GND.n9048 0.001
R10424 GND.n9047 GND.n8874 0.001
R10425 GND.n8873 GND.n8872 0.001
R10426 GND.n8871 GND.n8870 0.001
R10427 GND.n8869 GND.n8868 0.001
R10428 GND.n8867 GND.n8866 0.001
R10429 GND.n8864 GND.n8863 0.001
R10430 GND.n8862 GND.n8689 0.001
R10431 GND.n8688 GND.n8687 0.001
R10432 GND.n8686 GND.n8685 0.001
R10433 GND.n8684 GND.n8683 0.001
R10434 GND.n8682 GND.n8681 0.001
R10435 GND.n8679 GND.n8678 0.001
R10436 GND.n8677 GND.n8504 0.001
R10437 GND.n8503 GND.n8502 0.001
R10438 GND.n8501 GND.n8500 0.001
R10439 GND.n8499 GND.n8498 0.001
R10440 GND.n8497 GND.n8496 0.001
R10441 GND.n8494 GND.n8493 0.001
R10442 GND.n8492 GND.n8319 0.001
R10443 GND.n8318 GND.n8317 0.001
R10444 GND.n8316 GND.n8315 0.001
R10445 GND.n8314 GND.n8313 0.001
R10446 GND.n8312 GND.n8311 0.001
R10447 GND.n9248 GND.n9247 0.001
R10448 GND.n9242 GND.n9241 0.001
R10449 GND.n9238 GND.n9237 0.001
R10450 GND.n9246 GND.n9245 0.001
R10451 GND.n9240 GND.n9239 0.001
R10452 GND.n9244 GND.n9243 0.001
R10453 GND.n9233 GND.n9232 0.001
R10454 GND.n9057 GND.n9056 0.001
R10455 GND.n9053 GND.n9052 0.001
R10456 GND.n9235 GND.n9234 0.001
R10457 GND.n9055 GND.n9054 0.001
R10458 GND.n9059 GND.n9058 0.001
R10459 GND.n9048 GND.n9047 0.001
R10460 GND.n8872 GND.n8871 0.001
R10461 GND.n8868 GND.n8867 0.001
R10462 GND.n9050 GND.n9049 0.001
R10463 GND.n8870 GND.n8869 0.001
R10464 GND.n8874 GND.n8873 0.001
R10465 GND.n8863 GND.n8862 0.001
R10466 GND.n8687 GND.n8686 0.001
R10467 GND.n8683 GND.n8682 0.001
R10468 GND.n8865 GND.n8864 0.001
R10469 GND.n8685 GND.n8684 0.001
R10470 GND.n8689 GND.n8688 0.001
R10471 GND.n8678 GND.n8677 0.001
R10472 GND.n8502 GND.n8501 0.001
R10473 GND.n8498 GND.n8497 0.001
R10474 GND.n8680 GND.n8679 0.001
R10475 GND.n8500 GND.n8499 0.001
R10476 GND.n8504 GND.n8503 0.001
R10477 GND.n8493 GND.n8492 0.001
R10478 GND.n8317 GND.n8316 0.001
R10479 GND.n8313 GND.n8312 0.001
R10480 GND.n8495 GND.n8494 0.001
R10481 GND.n8315 GND.n8314 0.001
R10482 GND.n8319 GND.n8318 0.001
R10483 GND.n6699 GND.n6698 0.001
R10484 GND.n6701 GND.n6700 0.001
R10485 GND.n6899 GND.n6702 0.001
R10486 GND.n6901 GND.n6900 0.001
R10487 GND.n6903 GND.n6902 0.001
R10488 GND.n6923 GND.n6922 0.001
R10489 GND.n6926 GND.n6925 0.001
R10490 GND.n6928 GND.n6927 0.001
R10491 GND.n7126 GND.n6929 0.001
R10492 GND.n7128 GND.n7127 0.001
R10493 GND.n7130 GND.n7129 0.001
R10494 GND.n7150 GND.n7149 0.001
R10495 GND.n7153 GND.n7152 0.001
R10496 GND.n7155 GND.n7154 0.001
R10497 GND.n7353 GND.n7156 0.001
R10498 GND.n7355 GND.n7354 0.001
R10499 GND.n7357 GND.n7356 0.001
R10500 GND.n7377 GND.n7376 0.001
R10501 GND.n7380 GND.n7379 0.001
R10502 GND.n7382 GND.n7381 0.001
R10503 GND.n7580 GND.n7383 0.001
R10504 GND.n7582 GND.n7581 0.001
R10505 GND.n7584 GND.n7583 0.001
R10506 GND.n7604 GND.n7603 0.001
R10507 GND.n7607 GND.n7606 0.001
R10508 GND.n7609 GND.n7608 0.001
R10509 GND.n7807 GND.n7610 0.001
R10510 GND.n7809 GND.n7808 0.001
R10511 GND.n7811 GND.n7810 0.001
R10512 GND.n7831 GND.n7830 0.001
R10513 GND.n7834 GND.n7833 0.001
R10514 GND.n7836 GND.n7835 0.001
R10515 GND.n8034 GND.n7837 0.001
R10516 GND.n8036 GND.n8035 0.001
R10517 GND.n8038 GND.n8037 0.001
R10518 GND.n8058 GND.n8057 0.001
R10519 GND.n6700 GND.n6699 0.001
R10520 GND.n6900 GND.n6899 0.001
R10521 GND.n6922 GND.n6903 0.001
R10522 GND.n6698 GND.n6697 0.001
R10523 GND.n6902 GND.n6901 0.001
R10524 GND.n6702 GND.n6701 0.001
R10525 GND.n6927 GND.n6926 0.001
R10526 GND.n7127 GND.n7126 0.001
R10527 GND.n7149 GND.n7130 0.001
R10528 GND.n6925 GND.n6924 0.001
R10529 GND.n7129 GND.n7128 0.001
R10530 GND.n6929 GND.n6928 0.001
R10531 GND.n7154 GND.n7153 0.001
R10532 GND.n7354 GND.n7353 0.001
R10533 GND.n7376 GND.n7357 0.001
R10534 GND.n7152 GND.n7151 0.001
R10535 GND.n7356 GND.n7355 0.001
R10536 GND.n7156 GND.n7155 0.001
R10537 GND.n7381 GND.n7380 0.001
R10538 GND.n7581 GND.n7580 0.001
R10539 GND.n7603 GND.n7584 0.001
R10540 GND.n7379 GND.n7378 0.001
R10541 GND.n7583 GND.n7582 0.001
R10542 GND.n7383 GND.n7382 0.001
R10543 GND.n7608 GND.n7607 0.001
R10544 GND.n7808 GND.n7807 0.001
R10545 GND.n7830 GND.n7811 0.001
R10546 GND.n7606 GND.n7605 0.001
R10547 GND.n7810 GND.n7809 0.001
R10548 GND.n7610 GND.n7609 0.001
R10549 GND.n7835 GND.n7834 0.001
R10550 GND.n8035 GND.n8034 0.001
R10551 GND.n8057 GND.n8038 0.001
R10552 GND.n7833 GND.n7832 0.001
R10553 GND.n8037 GND.n8036 0.001
R10554 GND.n7837 GND.n7836 0.001
R10555 GND.n464 GND.n463 0.001
R10556 GND.n8070 GND.n8069 0.001
R10557 GND.n6354 GND.n6353 0.001
R10558 GND.n480 GND.n475 0.001
R10559 GND.n4361 GND.n4360 0.001
R10560 GND.n4365 GND.n4364 0.001
R10561 GND.n2203 GND.n2202 0.001
R10562 GND.n2220 GND.n2219 0.001
R10563 GND.n4320 GND.n4319 0.001
R10564 GND.n2234 GND.n2233 0.001
R10565 GND.n4323 GND.n4322 0.001
R10566 GND.n6589 GND.n6588 0.001
R10567 GND.n8071 GND.n8070 0.001
R10568 GND.n6580 GND.n6579 0.001
R10569 GND.n7974 GND.n7973 0.001
R10570 GND.n7992 GND.n7984 0.001
R10571 GND.n8004 GND.n7994 0.001
R10572 GND.n7886 GND.n7885 0.001
R10573 GND.n6599 GND.n6598 0.001
R10574 GND.n6603 GND.n6602 0.001
R10575 GND.n7839 GND.n7838 0.001
R10576 GND.n8055 GND.n8047 0.001
R10577 GND.n8054 GND.n8053 0.001
R10578 GND.n8050 GND.n8049 0.001
R10579 GND.n6610 GND.n6609 0.001
R10580 GND.n6609 GND.n6608 0.001
R10581 GND.n8040 GND.n8039 0.001
R10582 GND.n8041 GND.n8040 0.001
R10583 GND.n7747 GND.n7746 0.001
R10584 GND.n7765 GND.n7757 0.001
R10585 GND.n7777 GND.n7767 0.001
R10586 GND.n7659 GND.n7658 0.001
R10587 GND.n6616 GND.n6615 0.001
R10588 GND.n6620 GND.n6619 0.001
R10589 GND.n7612 GND.n7611 0.001
R10590 GND.n7828 GND.n7820 0.001
R10591 GND.n7827 GND.n7826 0.001
R10592 GND.n7823 GND.n7822 0.001
R10593 GND.n6627 GND.n6626 0.001
R10594 GND.n6626 GND.n6625 0.001
R10595 GND.n7813 GND.n7812 0.001
R10596 GND.n7814 GND.n7813 0.001
R10597 GND.n7520 GND.n7519 0.001
R10598 GND.n7538 GND.n7530 0.001
R10599 GND.n7550 GND.n7540 0.001
R10600 GND.n7432 GND.n7431 0.001
R10601 GND.n6633 GND.n6632 0.001
R10602 GND.n6637 GND.n6636 0.001
R10603 GND.n7385 GND.n7384 0.001
R10604 GND.n7601 GND.n7593 0.001
R10605 GND.n7600 GND.n7599 0.001
R10606 GND.n7596 GND.n7595 0.001
R10607 GND.n6644 GND.n6643 0.001
R10608 GND.n6643 GND.n6642 0.001
R10609 GND.n7586 GND.n7585 0.001
R10610 GND.n7587 GND.n7586 0.001
R10611 GND.n7293 GND.n7292 0.001
R10612 GND.n7311 GND.n7303 0.001
R10613 GND.n7323 GND.n7313 0.001
R10614 GND.n7205 GND.n7204 0.001
R10615 GND.n6650 GND.n6649 0.001
R10616 GND.n6654 GND.n6653 0.001
R10617 GND.n7158 GND.n7157 0.001
R10618 GND.n7374 GND.n7366 0.001
R10619 GND.n7373 GND.n7372 0.001
R10620 GND.n7369 GND.n7368 0.001
R10621 GND.n6661 GND.n6660 0.001
R10622 GND.n6660 GND.n6659 0.001
R10623 GND.n7359 GND.n7358 0.001
R10624 GND.n7360 GND.n7359 0.001
R10625 GND.n7066 GND.n7065 0.001
R10626 GND.n7084 GND.n7076 0.001
R10627 GND.n7096 GND.n7086 0.001
R10628 GND.n6978 GND.n6977 0.001
R10629 GND.n6667 GND.n6666 0.001
R10630 GND.n6671 GND.n6670 0.001
R10631 GND.n6931 GND.n6930 0.001
R10632 GND.n7147 GND.n7139 0.001
R10633 GND.n7146 GND.n7145 0.001
R10634 GND.n7142 GND.n7141 0.001
R10635 GND.n6678 GND.n6677 0.001
R10636 GND.n6677 GND.n6676 0.001
R10637 GND.n7132 GND.n7131 0.001
R10638 GND.n7133 GND.n7132 0.001
R10639 GND.n6839 GND.n6838 0.001
R10640 GND.n6857 GND.n6849 0.001
R10641 GND.n6869 GND.n6859 0.001
R10642 GND.n6751 GND.n6750 0.001
R10643 GND.n6684 GND.n6683 0.001
R10644 GND.n6688 GND.n6687 0.001
R10645 GND.n6704 GND.n6703 0.001
R10646 GND.n6920 GND.n6912 0.001
R10647 GND.n6919 GND.n6918 0.001
R10648 GND.n6915 GND.n6914 0.001
R10649 GND.n6695 GND.n6694 0.001
R10650 GND.n6694 GND.n6693 0.001
R10651 GND.n6905 GND.n6904 0.001
R10652 GND.n6906 GND.n6905 0.001
R10653 GND.n6507 GND.n6506 0.001
R10654 GND.n6525 GND.n6517 0.001
R10655 GND.n6537 GND.n6527 0.001
R10656 GND.n6431 GND.n6430 0.001
R10657 GND.n6366 GND.n6365 0.001
R10658 GND.n6371 GND.n6370 0.001
R10659 GND.n6582 GND.n6581 0.001
R10660 GND.n6575 GND.n6574 0.001
R10661 GND.n6573 GND.n6572 0.001
R10662 GND.n6568 GND.n6567 0.001
R10663 GND.n572 GND.n571 0.001
R10664 GND.n1003 GND.n1002 0.001
R10665 GND.n6042 GND.n6041 0.001
R10666 GND.n6122 GND.n1088 0.001
R10667 GND.n6139 GND.n6138 0.001
R10668 GND.n1283 GND.n1281 0.001
R10669 GND.n1271 GND.n1267 0.001
R10670 GND.n2625 GND.n2624 0.001
R10671 GND.n3870 GND.n3869 0.001
R10672 GND.n3950 GND.n2710 0.001
R10673 GND.n3967 GND.n3966 0.001
R10674 GND.n3783 GND.n3778 0.001
R10675 GND.n4353 GND.n4352 0.001
R10676 GND.n4369 GND.n4368 0.001
R10677 GND.n4357 GND.n4356 0.001
R10678 GND.n4386 GND.n4385 0.001
R10679 GND.n2242 GND.n2241 0.001
R10680 GND.n2245 GND.n2244 0.001
R10681 GND.n2247 GND.n2246 0.001
R10682 GND.n4312 GND.n4311 0.001
R10683 GND.n4308 GND.n4307 0.001
R10684 GND.n2338 GND.n2337 0.001
R10685 GND.n4011 GND.n4009 0.001
R10686 GND.n3012 GND.n3011 0.001
R10687 GND.n4123 GND.n4122 0.001
R10688 GND.n2897 GND.n2894 0.001
R10689 GND.n4298 GND.n4297 0.001
R10690 GND.n6307 GND.n6305 0.001
R10691 GND.n1591 GND.n1590 0.001
R10692 GND.n6165 GND.n6164 0.001
R10693 GND.n1470 GND.n1467 0.001
R10694 GND.n6315 GND.n6314 0.001
R10695 GND.n6342 GND.n6341 0.001
R10696 GND.n6347 GND.n6346 0.001
R10697 GND.n460 GND.n459 0.001
R10698 GND.n484 GND.n483 0.001
R10699 GND.n6361 GND.n6360 0.001
R10700 GND.n8093 GND.n8092 0.001
R10701 GND.n8111 GND.n8110 0.001
R10702 GND.n8123 GND.n8122 0.001
R10703 GND.n8090 GND.n8089 0.001
R10704 GND.n8101 GND.n8098 0.001
R10705 GND.n8112 GND.n8109 0.001
R10706 GND.n8114 GND.n8113 0.001
R10707 GND.n8302 GND.n8298 0.001
R10708 GND.n8297 GND.n8293 0.001
R10709 GND.n8291 GND.n8290 0.001
R10710 GND.n8143 GND.n8142 0.001
R10711 GND.n8133 GND.n8132 0.001
R10712 GND.n8131 GND.n8128 0.001
R10713 GND.n430 GND.n429 0.001
R10714 GND.n448 GND.n447 0.001
R10715 GND.n8473 GND.n8472 0.001
R10716 GND.n438 GND.n435 0.001
R10717 GND.n450 GND.n445 0.001
R10718 GND.n421 GND.n420 0.001
R10719 GND.n419 GND.n415 0.001
R10720 GND.n8469 GND.n8323 0.001
R10721 GND.n8490 GND.n8470 0.001
R10722 GND.n8482 GND.n8481 0.001
R10723 GND.n404 GND.n403 0.001
R10724 GND.n405 GND.n404 0.001
R10725 GND.n423 GND.n422 0.001
R10726 GND.n381 GND.n380 0.001
R10727 GND.n399 GND.n398 0.001
R10728 GND.n8658 GND.n8657 0.001
R10729 GND.n389 GND.n386 0.001
R10730 GND.n401 GND.n396 0.001
R10731 GND.n372 GND.n371 0.001
R10732 GND.n370 GND.n366 0.001
R10733 GND.n8654 GND.n8508 0.001
R10734 GND.n8675 GND.n8655 0.001
R10735 GND.n8667 GND.n8666 0.001
R10736 GND.n355 GND.n354 0.001
R10737 GND.n356 GND.n355 0.001
R10738 GND.n374 GND.n373 0.001
R10739 GND.n332 GND.n331 0.001
R10740 GND.n350 GND.n349 0.001
R10741 GND.n8843 GND.n8842 0.001
R10742 GND.n340 GND.n337 0.001
R10743 GND.n352 GND.n347 0.001
R10744 GND.n323 GND.n322 0.001
R10745 GND.n321 GND.n317 0.001
R10746 GND.n8839 GND.n8693 0.001
R10747 GND.n8860 GND.n8840 0.001
R10748 GND.n8852 GND.n8851 0.001
R10749 GND.n306 GND.n305 0.001
R10750 GND.n307 GND.n306 0.001
R10751 GND.n325 GND.n324 0.001
R10752 GND.n283 GND.n282 0.001
R10753 GND.n301 GND.n300 0.001
R10754 GND.n9028 GND.n9027 0.001
R10755 GND.n291 GND.n288 0.001
R10756 GND.n303 GND.n298 0.001
R10757 GND.n274 GND.n273 0.001
R10758 GND.n272 GND.n268 0.001
R10759 GND.n9024 GND.n8878 0.001
R10760 GND.n9045 GND.n9025 0.001
R10761 GND.n9037 GND.n9036 0.001
R10762 GND.n257 GND.n256 0.001
R10763 GND.n258 GND.n257 0.001
R10764 GND.n276 GND.n275 0.001
R10765 GND.n234 GND.n233 0.001
R10766 GND.n252 GND.n251 0.001
R10767 GND.n9213 GND.n9212 0.001
R10768 GND.n242 GND.n239 0.001
R10769 GND.n254 GND.n249 0.001
R10770 GND.n225 GND.n224 0.001
R10771 GND.n223 GND.n219 0.001
R10772 GND.n9209 GND.n9063 0.001
R10773 GND.n9230 GND.n9210 0.001
R10774 GND.n9222 GND.n9221 0.001
R10775 GND.n208 GND.n207 0.001
R10776 GND.n209 GND.n208 0.001
R10777 GND.n227 GND.n226 0.001
R10778 GND.n2 GND.n1 0.001
R10779 GND.n14 GND.n13 0.001
R10780 GND.n172 GND.n171 0.001
R10781 GND.n181 GND.n180 0.001
R10782 GND.n185 GND.n184 0.001
R10783 GND.n187 GND.n186 0.001
R10784 GND.n191 GND.n190 0.001
R10785 GND.n193 GND.n192 0.001
R10786 GND.n195 GND.n194 0.001
R10787 GND.n9252 GND.n196 0.001
R10788 GND.n9256 GND.n9255 0.001
R10789 GND.n201 GND.n200 0.001
R10790 GND.n202 GND.n201 0.001
R10791 GND.n205 GND.n204 0.001
R10792 GND.n206 GND.n205 0.001
R10793 GND.n479 GND.n477 0.001
R10794 GND.n2198 GND.n2197 0.001
R10795 GND.n2199 GND.n2198 0.001
R10796 GND.n467 GND.n466 0.001
R10797 GND.n469 GND.n468 0.001
R10798 GND.n466 GND.n465 0.001
R10799 GND.n470 GND.n469 0.001
R10800 GND.n2216 GND.n2215 0.001
R10801 GND.n4335 GND.n4334 0.001
R10802 GND.n8303 GND.n8088 0.001
R10803 GND.n8306 GND.n8085 0.001
R10804 GND.n8088 GND.n8087 0.001
R10805 GND.n8080 GND.n8079 0.001
R10806 GND.n8081 GND.n8080 0.001
R10807 GND.n6590 GND.n6589 0.001
R10808 GND.n8066 GND.n6594 0.001
R10809 GND.n6353 GND.n6352 0.001
R10810 GND.n8084 GND.n8083 0.001
R10811 GND.n8083 GND.n8082 0.001
R10812 GND.n6592 GND.n6591 0.001
R10813 GND.n6593 GND.n6592 0.001
R10814 OUT_N.n1173 OUT_N.t16 846.712
R10815 OUT_N.n1155 OUT_N.t23 846.712
R10816 OUT_N.n1100 OUT_N.t27 846.712
R10817 OUT_N.n1082 OUT_N.t25 846.712
R10818 OUT_N.n78 OUT_N.t18 846.712
R10819 OUT_N.n94 OUT_N.t19 846.712
R10820 OUT_N.n43 OUT_N.t14 846.712
R10821 OUT_N.n59 OUT_N.t15 846.712
R10822 OUT_N.n8 OUT_N.t21 846.712
R10823 OUT_N.n24 OUT_N.t17 846.712
R10824 OUT_N.n1252 OUT_N.t24 846.712
R10825 OUT_N.n1244 OUT_N.t20 846.712
R10826 OUT_N.n1312 OUT_N.t26 846.712
R10827 OUT_N.n1289 OUT_N.t22 846.712
R10828 OUT_N.n1174 OUT_N.n1173 24.127
R10829 OUT_N.n1156 OUT_N.n1155 24.127
R10830 OUT_N.n1000 OUT_N.n999 24.127
R10831 OUT_N.n1005 OUT_N.n1004 24.127
R10832 OUT_N.n1101 OUT_N.n1100 24.127
R10833 OUT_N.n1083 OUT_N.n1082 24.127
R10834 OUT_N.n974 OUT_N.n973 24.127
R10835 OUT_N.n979 OUT_N.n978 24.127
R10836 OUT_N.n95 OUT_N.n94 24.127
R10837 OUT_N.n79 OUT_N.n78 24.127
R10838 OUT_N.n228 OUT_N.n227 24.127
R10839 OUT_N.n232 OUT_N.n231 24.127
R10840 OUT_N.n60 OUT_N.n59 24.127
R10841 OUT_N.n44 OUT_N.n43 24.127
R10842 OUT_N.n191 OUT_N.n190 24.127
R10843 OUT_N.n195 OUT_N.n194 24.127
R10844 OUT_N.n25 OUT_N.n24 24.127
R10845 OUT_N.n9 OUT_N.n8 24.127
R10846 OUT_N.n154 OUT_N.n153 24.127
R10847 OUT_N.n158 OUT_N.n157 24.127
R10848 OUT_N.n1245 OUT_N.n1244 24.127
R10849 OUT_N.n1253 OUT_N.n1252 24.127
R10850 OUT_N.n122 OUT_N.n121 24.127
R10851 OUT_N.n126 OUT_N.n125 24.127
R10852 OUT_N.n1040 OUT_N.n1039 24.127
R10853 OUT_N.n1027 OUT_N.n1026 24.127
R10854 OUT_N.n1290 OUT_N.n1289 24.127
R10855 OUT_N.n1313 OUT_N.n1312 24.127
R10856 OUT_N.n603 OUT_N.n602 9.309
R10857 OUT_N.n702 OUT_N.n701 9.309
R10858 OUT_N.n801 OUT_N.n800 9.309
R10859 OUT_N.n900 OUT_N.n899 9.309
R10860 OUT_N.n261 OUT_N.n260 9.3
R10861 OUT_N.n264 OUT_N.n263 9.3
R10862 OUT_N.n320 OUT_N.n319 9.3
R10863 OUT_N.n318 OUT_N.n317 9.3
R10864 OUT_N.n326 OUT_N.n325 9.3
R10865 OUT_N.n314 OUT_N.n313 9.3
R10866 OUT_N.n304 OUT_N.n303 9.3
R10867 OUT_N.n307 OUT_N.n306 9.3
R10868 OUT_N.n309 OUT_N.n308 9.3
R10869 OUT_N.n288 OUT_N.n287 9.3
R10870 OUT_N.n274 OUT_N.n273 9.3
R10871 OUT_N.n279 OUT_N.n278 9.3
R10872 OUT_N.n283 OUT_N.n282 9.3
R10873 OUT_N.n269 OUT_N.n268 9.3
R10874 OUT_N.n360 OUT_N.n359 9.3
R10875 OUT_N.n363 OUT_N.n362 9.3
R10876 OUT_N.n419 OUT_N.n418 9.3
R10877 OUT_N.n417 OUT_N.n416 9.3
R10878 OUT_N.n425 OUT_N.n424 9.3
R10879 OUT_N.n413 OUT_N.n412 9.3
R10880 OUT_N.n403 OUT_N.n402 9.3
R10881 OUT_N.n406 OUT_N.n405 9.3
R10882 OUT_N.n408 OUT_N.n407 9.3
R10883 OUT_N.n387 OUT_N.n386 9.3
R10884 OUT_N.n373 OUT_N.n372 9.3
R10885 OUT_N.n378 OUT_N.n377 9.3
R10886 OUT_N.n382 OUT_N.n381 9.3
R10887 OUT_N.n368 OUT_N.n367 9.3
R10888 OUT_N.n459 OUT_N.n458 9.3
R10889 OUT_N.n462 OUT_N.n461 9.3
R10890 OUT_N.n518 OUT_N.n517 9.3
R10891 OUT_N.n516 OUT_N.n515 9.3
R10892 OUT_N.n524 OUT_N.n523 9.3
R10893 OUT_N.n512 OUT_N.n511 9.3
R10894 OUT_N.n502 OUT_N.n501 9.3
R10895 OUT_N.n505 OUT_N.n504 9.3
R10896 OUT_N.n507 OUT_N.n506 9.3
R10897 OUT_N.n486 OUT_N.n485 9.3
R10898 OUT_N.n472 OUT_N.n471 9.3
R10899 OUT_N.n477 OUT_N.n476 9.3
R10900 OUT_N.n481 OUT_N.n480 9.3
R10901 OUT_N.n467 OUT_N.n466 9.3
R10902 OUT_N.n1176 OUT_N.n1175 9.3
R10903 OUT_N.n1158 OUT_N.n1157 9.3
R10904 OUT_N.n1103 OUT_N.n1102 9.3
R10905 OUT_N.n1085 OUT_N.n1084 9.3
R10906 OUT_N.n598 OUT_N.n597 9.3
R10907 OUT_N.n641 OUT_N.n640 9.3
R10908 OUT_N.n636 OUT_N.n635 9.3
R10909 OUT_N.n594 OUT_N.n593 9.3
R10910 OUT_N.n588 OUT_N.n587 9.3
R10911 OUT_N.n583 OUT_N.n582 9.3
R10912 OUT_N.n634 OUT_N.n633 9.3
R10913 OUT_N.n647 OUT_N.n646 9.3
R10914 OUT_N.n645 OUT_N.n644 9.3
R10915 OUT_N.n652 OUT_N.n651 9.3
R10916 OUT_N.n658 OUT_N.n657 9.3
R10917 OUT_N.n656 OUT_N.n655 9.3
R10918 OUT_N.n629 OUT_N.n628 9.3
R10919 OUT_N.n764 OUT_N.n763 9.3
R10920 OUT_N.n697 OUT_N.n696 9.3
R10921 OUT_N.n745 OUT_N.n744 9.3
R10922 OUT_N.n730 OUT_N.n729 9.3
R10923 OUT_N.n725 OUT_N.n724 9.3
R10924 OUT_N.n693 OUT_N.n692 9.3
R10925 OUT_N.n687 OUT_N.n686 9.3
R10926 OUT_N.n682 OUT_N.n681 9.3
R10927 OUT_N.n723 OUT_N.n722 9.3
R10928 OUT_N.n736 OUT_N.n735 9.3
R10929 OUT_N.n734 OUT_N.n733 9.3
R10930 OUT_N.n741 OUT_N.n740 9.3
R10931 OUT_N.n747 OUT_N.n746 9.3
R10932 OUT_N.n863 OUT_N.n862 9.3
R10933 OUT_N.n796 OUT_N.n795 9.3
R10934 OUT_N.n844 OUT_N.n843 9.3
R10935 OUT_N.n829 OUT_N.n828 9.3
R10936 OUT_N.n824 OUT_N.n823 9.3
R10937 OUT_N.n792 OUT_N.n791 9.3
R10938 OUT_N.n786 OUT_N.n785 9.3
R10939 OUT_N.n781 OUT_N.n780 9.3
R10940 OUT_N.n822 OUT_N.n821 9.3
R10941 OUT_N.n835 OUT_N.n834 9.3
R10942 OUT_N.n833 OUT_N.n832 9.3
R10943 OUT_N.n840 OUT_N.n839 9.3
R10944 OUT_N.n846 OUT_N.n845 9.3
R10945 OUT_N.n962 OUT_N.n961 9.3
R10946 OUT_N.n895 OUT_N.n894 9.3
R10947 OUT_N.n943 OUT_N.n942 9.3
R10948 OUT_N.n928 OUT_N.n927 9.3
R10949 OUT_N.n923 OUT_N.n922 9.3
R10950 OUT_N.n891 OUT_N.n890 9.3
R10951 OUT_N.n885 OUT_N.n884 9.3
R10952 OUT_N.n880 OUT_N.n879 9.3
R10953 OUT_N.n921 OUT_N.n920 9.3
R10954 OUT_N.n934 OUT_N.n933 9.3
R10955 OUT_N.n932 OUT_N.n931 9.3
R10956 OUT_N.n939 OUT_N.n938 9.3
R10957 OUT_N.n945 OUT_N.n944 9.3
R10958 OUT_N.n81 OUT_N.n80 9.3
R10959 OUT_N.n46 OUT_N.n45 9.3
R10960 OUT_N.n11 OUT_N.n10 9.3
R10961 OUT_N.n1255 OUT_N.n1254 9.3
R10962 OUT_N.n1292 OUT_N.n1291 9.3
R10963 OUT_N.n1315 OUT_N.n1314 9.3
R10964 OUT_N.n327 OUT_N.n297 9
R10965 OUT_N.n305 OUT_N.n302 9
R10966 OUT_N.n321 OUT_N.n301 9
R10967 OUT_N.n316 OUT_N.n315 9
R10968 OUT_N.n276 OUT_N.n275 9
R10969 OUT_N.n286 OUT_N.n285 9
R10970 OUT_N.n266 OUT_N.n265 9
R10971 OUT_N.n426 OUT_N.n396 9
R10972 OUT_N.n404 OUT_N.n401 9
R10973 OUT_N.n420 OUT_N.n400 9
R10974 OUT_N.n415 OUT_N.n414 9
R10975 OUT_N.n375 OUT_N.n374 9
R10976 OUT_N.n385 OUT_N.n384 9
R10977 OUT_N.n365 OUT_N.n364 9
R10978 OUT_N.n525 OUT_N.n495 9
R10979 OUT_N.n503 OUT_N.n500 9
R10980 OUT_N.n519 OUT_N.n499 9
R10981 OUT_N.n514 OUT_N.n513 9
R10982 OUT_N.n474 OUT_N.n473 9
R10983 OUT_N.n484 OUT_N.n483 9
R10984 OUT_N.n464 OUT_N.n463 9
R10985 OUT_N.n660 OUT_N.n659 9
R10986 OUT_N.n654 OUT_N.n653 9
R10987 OUT_N.n643 OUT_N.n642 9
R10988 OUT_N.n590 OUT_N.n589 9
R10989 OUT_N.n632 OUT_N.n631 9
R10990 OUT_N.n601 OUT_N.n600 9
R10991 OUT_N.n626 OUT_N.n621 9
R10992 OUT_N.n732 OUT_N.n731 9
R10993 OUT_N.n689 OUT_N.n688 9
R10994 OUT_N.n721 OUT_N.n720 9
R10995 OUT_N.n749 OUT_N.n748 9
R10996 OUT_N.n743 OUT_N.n742 9
R10997 OUT_N.n700 OUT_N.n699 9
R10998 OUT_N.n761 OUT_N.n756 9
R10999 OUT_N.n831 OUT_N.n830 9
R11000 OUT_N.n788 OUT_N.n787 9
R11001 OUT_N.n820 OUT_N.n819 9
R11002 OUT_N.n848 OUT_N.n847 9
R11003 OUT_N.n842 OUT_N.n841 9
R11004 OUT_N.n799 OUT_N.n798 9
R11005 OUT_N.n860 OUT_N.n855 9
R11006 OUT_N.n930 OUT_N.n929 9
R11007 OUT_N.n887 OUT_N.n886 9
R11008 OUT_N.n919 OUT_N.n918 9
R11009 OUT_N.n947 OUT_N.n946 9
R11010 OUT_N.n941 OUT_N.n940 9
R11011 OUT_N.n898 OUT_N.n897 9
R11012 OUT_N.n959 OUT_N.n954 9
R11013 OUT_N.n1251 OUT_N.n1250 9
R11014 OUT_N.n1288 OUT_N.n2 9
R11015 OUT_N.n1317 OUT_N.n1316 9
R11016 OUT_N.n7 OUT_N.n6 9
R11017 OUT_N.n1178 OUT_N.n1177 9
R11018 OUT_N.n1154 OUT_N.n1153 9
R11019 OUT_N.n42 OUT_N.n41 9
R11020 OUT_N.n1105 OUT_N.n1104 9
R11021 OUT_N.n1081 OUT_N.n1080 9
R11022 OUT_N.n77 OUT_N.n76 9
R11023 OUT_N.n1165 OUT_N.n1164 8.764
R11024 OUT_N.n1002 OUT_N.n1001 8.764
R11025 OUT_N.n1092 OUT_N.n1091 8.764
R11026 OUT_N.n976 OUT_N.n975 8.764
R11027 OUT_N.n88 OUT_N.n87 8.764
R11028 OUT_N.n230 OUT_N.n229 8.764
R11029 OUT_N.n53 OUT_N.n52 8.764
R11030 OUT_N.n193 OUT_N.n192 8.764
R11031 OUT_N.n18 OUT_N.n17 8.764
R11032 OUT_N.n156 OUT_N.n155 8.764
R11033 OUT_N.n1262 OUT_N.n1261 8.764
R11034 OUT_N.n124 OUT_N.n123 8.764
R11035 OUT_N.n1035 OUT_N.n1034 8.764
R11036 OUT_N.n1300 OUT_N.n1299 8.764
R11037 OUT_N.n295 OUT_N.n294 8.043
R11038 OUT_N.n394 OUT_N.n393 8.043
R11039 OUT_N.n493 OUT_N.n492 8.043
R11040 OUT_N.n1007 OUT_N.n1006 6.364
R11041 OUT_N.n981 OUT_N.n980 6.364
R11042 OUT_N.n235 OUT_N.n233 6.364
R11043 OUT_N.n198 OUT_N.n196 6.364
R11044 OUT_N.n161 OUT_N.n159 6.364
R11045 OUT_N.n129 OUT_N.n127 6.364
R11046 OUT_N.n1029 OUT_N.n1028 6.364
R11047 OUT_N.n669 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN 6.312
R11048 OUT_N.n768 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/DRAIN 6.312
R11049 OUT_N.n867 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/DRAIN 6.312
R11050 OUT_N.n966 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/DRAIN 6.312
R11051 OUT_N.n323 OUT_N.n300 4.574
R11052 OUT_N.n422 OUT_N.n399 4.574
R11053 OUT_N.n521 OUT_N.n498 4.574
R11054 OUT_N.n1012 OUT_N.n1002 4.574
R11055 OUT_N.n986 OUT_N.n976 4.574
R11056 OUT_N.n666 OUT_N.n665 4.574
R11057 OUT_N.n755 OUT_N.n754 4.574
R11058 OUT_N.n854 OUT_N.n853 4.574
R11059 OUT_N.n953 OUT_N.n952 4.574
R11060 OUT_N.n241 OUT_N.n230 4.574
R11061 OUT_N.n204 OUT_N.n193 4.574
R11062 OUT_N.n167 OUT_N.n156 4.574
R11063 OUT_N.n1263 OUT_N.n1262 4.574
R11064 OUT_N.n135 OUT_N.n124 4.574
R11065 OUT_N.n1036 OUT_N.n1035 4.574
R11066 OUT_N.n1301 OUT_N.n1300 4.574
R11067 OUT_N.n19 OUT_N.n18 4.574
R11068 OUT_N.n1166 OUT_N.n1165 4.574
R11069 OUT_N.n54 OUT_N.n53 4.574
R11070 OUT_N.n1093 OUT_N.n1092 4.574
R11071 OUT_N.n89 OUT_N.n88 4.574
R11072 OUT_N.n1267 OUT_N.n1245 4.558
R11073 OUT_N.n26 OUT_N.n25 4.557
R11074 OUT_N.n61 OUT_N.n60 4.557
R11075 OUT_N.n96 OUT_N.n95 4.557
R11076 OUT_N.n244 OUT_N.n228 4.555
R11077 OUT_N.n207 OUT_N.n191 4.555
R11078 OUT_N.n170 OUT_N.n154 4.555
R11079 OUT_N.n138 OUT_N.n122 4.553
R11080 OUT_N.n1015 OUT_N.n1000 4.552
R11081 OUT_N.n989 OUT_N.n974 4.552
R11082 OUT_N.n1041 OUT_N.n1040 4.552
R11083 OUT_N.n73 OUT_N 4.125
R11084 OUT_N.n38 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/GATE 4.125
R11085 OUT_N.n3 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE 4.125
R11086 OUT_N.n1310 OUT_N.n1309 3.41
R11087 OUT_N.n300 OUT_N.n298 3.388
R11088 OUT_N.n399 OUT_N.n397 3.388
R11089 OUT_N.n498 OUT_N.n496 3.388
R11090 OUT_N.n665 OUT_N.n664 3.388
R11091 OUT_N.n754 OUT_N.n753 3.388
R11092 OUT_N.n853 OUT_N.n852 3.388
R11093 OUT_N.n952 OUT_N.n951 3.388
R11094 OUT_N.n295 OUT_N.t11 3.326
R11095 OUT_N.n295 OUT_N.t0 3.326
R11096 OUT_N.n394 OUT_N.t2 3.326
R11097 OUT_N.n394 OUT_N.t4 3.326
R11098 OUT_N.n493 OUT_N.t3 3.326
R11099 OUT_N.n493 OUT_N.t13 3.326
R11100 OUT_N.n622 OUT_N.t6 3.326
R11101 OUT_N.n622 OUT_N.t8 3.326
R11102 OUT_N.n757 OUT_N.t9 3.326
R11103 OUT_N.n757 OUT_N.t12 3.326
R11104 OUT_N.n856 OUT_N.t1 3.326
R11105 OUT_N.n856 OUT_N.t7 3.326
R11106 OUT_N.n955 OUT_N.t10 3.326
R11107 OUT_N.n955 OUT_N.t5 3.326
R11108 OUT_N.n1288 OUT_N.n1287 3
R11109 OUT_N.n1179 OUT_N.n1178 3
R11110 OUT_N.n1106 OUT_N.n1105 3
R11111 OUT_N.n604 OUT_N.n603 2.253
R11112 OUT_N.n703 OUT_N.n702 2.253
R11113 OUT_N.n802 OUT_N.n801 2.253
R11114 OUT_N.n901 OUT_N.n900 2.253
R11115 OUT_N.n769 OUT_N.n766 2.25
R11116 OUT_N.n868 OUT_N.n865 2.25
R11117 OUT_N.n967 OUT_N.n964 2.25
R11118 OUT_N.n670 OUT_N.n667 2.25
R11119 OUT_N.n491 OUT_N.n487 1.94
R11120 OUT_N.n392 OUT_N.n388 1.94
R11121 OUT_N.n293 OUT_N.n289 1.94
R11122 OUT_N.n1024 OUT_N.n1015 1.805
R11123 OUT_N.n998 OUT_N.n989 1.805
R11124 OUT_N.n1050 OUT_N.n1041 1.805
R11125 OUT_N.n329 OUT_N.n328 1.801
R11126 OUT_N.n428 OUT_N.n427 1.801
R11127 OUT_N.n527 OUT_N.n526 1.801
R11128 OUT_N.n972 OUT_N.n561 1.705
R11129 OUT_N.n873 OUT_N.n566 1.705
R11130 OUT_N.n774 OUT_N.n571 1.705
R11131 OUT_N.n675 OUT_N.n576 1.705
R11132 OUT_N.n675 OUT_N.n674 1.705
R11133 OUT_N.n774 OUT_N.n773 1.705
R11134 OUT_N.n873 OUT_N.n872 1.705
R11135 OUT_N.n972 OUT_N.n971 1.705
R11136 OUT_N.n1055 OUT_N.n998 1.705
R11137 OUT_N.n1053 OUT_N.n1024 1.705
R11138 OUT_N.n1051 OUT_N.n1050 1.705
R11139 OUT_N.n1212 OUT_N.n1211 1.705
R11140 OUT_N.n1139 OUT_N.n1138 1.705
R11141 OUT_N.n1066 OUT_N.n1065 1.705
R11142 OUT_N.n1056 OUT_N.n1055 1.474
R11143 OUT_N.n1149 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/GATE 1.375
R11144 OUT_N.n1076 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/GATE 1.375
R11145 OUT_N.n1246 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE 1.375
R11146 OUT_N.n1321 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/GATE 1.375
R11147 OUT_N.n254 OUT_N.n253 1.227
R11148 OUT_N.n27 OUT_N.n26 1.188
R11149 OUT_N.n62 OUT_N.n61 1.188
R11150 OUT_N.n97 OUT_N.n96 1.188
R11151 OUT_N.n1268 OUT_N.n1267 1.187
R11152 OUT_N.n139 OUT_N.n138 1.183
R11153 OUT_N.n245 OUT_N.n244 1.183
R11154 OUT_N.n208 OUT_N.n207 1.183
R11155 OUT_N.n171 OUT_N.n170 1.183
R11156 OUT_N.n296 OUT_N.n295 1.155
R11157 OUT_N.n395 OUT_N.n394 1.155
R11158 OUT_N.n494 OUT_N.n493 1.155
R11159 OUT_N.n623 OUT_N.n622 1.155
R11160 OUT_N.n758 OUT_N.n757 1.155
R11161 OUT_N.n857 OUT_N.n856 1.155
R11162 OUT_N.n956 OUT_N.n955 1.155
R11163 OUT_N.n1275 OUT_N.n1274 1.137
R11164 OUT_N.n1239 OUT_N.n1238 1.137
R11165 OUT_N.n252 OUT_N.n251 1.137
R11166 OUT_N.n224 OUT_N.n223 1.137
R11167 OUT_N.n215 OUT_N.n214 1.137
R11168 OUT_N.n187 OUT_N.n186 1.137
R11169 OUT_N.n178 OUT_N.n177 1.137
R11170 OUT_N.n150 OUT_N.n149 1.137
R11171 OUT_N.n141 OUT_N.n140 1.137
R11172 OUT_N.n1284 OUT_N.n1283 1.137
R11173 OUT_N.n1203 OUT_N.n1202 1.137
R11174 OUT_N.n1186 OUT_N.n1185 1.137
R11175 OUT_N.n1130 OUT_N.n1129 1.137
R11176 OUT_N.n1113 OUT_N.n1112 1.137
R11177 OUT_N.n550 OUT_N.n549 1.135
R11178 OUT_N.n451 OUT_N.n450 1.135
R11179 OUT_N.n352 OUT_N.n351 1.135
R11180 OUT_N.n328 OUT_N.n296 0.935
R11181 OUT_N.n427 OUT_N.n395 0.935
R11182 OUT_N.n526 OUT_N.n494 0.935
R11183 OUT_N.n624 OUT_N.n623 0.893
R11184 OUT_N.n759 OUT_N.n758 0.893
R11185 OUT_N.n858 OUT_N.n857 0.893
R11186 OUT_N.n957 OUT_N.n956 0.893
R11187 OUT_N.n119 OUT_N.n118 0.868
R11188 OUT_N.n1058 OUT_N.n1057 0.853
R11189 OUT_N.n256 OUT_N.n255 0.848
R11190 OUT_N.n1157 OUT_N.n1156 0.77
R11191 OUT_N.n1175 OUT_N.n1174 0.77
R11192 OUT_N.n1006 OUT_N.n1005 0.77
R11193 OUT_N.n1084 OUT_N.n1083 0.77
R11194 OUT_N.n1102 OUT_N.n1101 0.77
R11195 OUT_N.n980 OUT_N.n979 0.77
R11196 OUT_N.n80 OUT_N.n79 0.77
R11197 OUT_N.n233 OUT_N.n232 0.77
R11198 OUT_N.n45 OUT_N.n44 0.77
R11199 OUT_N.n196 OUT_N.n195 0.77
R11200 OUT_N.n10 OUT_N.n9 0.77
R11201 OUT_N.n159 OUT_N.n158 0.77
R11202 OUT_N.n1254 OUT_N.n1253 0.77
R11203 OUT_N.n127 OUT_N.n126 0.77
R11204 OUT_N.n1028 OUT_N.n1027 0.77
R11205 OUT_N.n1291 OUT_N.n1290 0.77
R11206 OUT_N.n1314 OUT_N.n1313 0.77
R11207 OUT_N.n1218 OUT_N.n1217 0.672
R11208 OUT_N.n1145 OUT_N.n1144 0.672
R11209 OUT_N.n1072 OUT_N.n1071 0.672
R11210 OUT_N.n1056 OUT_N.n972 0.648
R11211 OUT_N.n1059 OUT_N.n1058 0.595
R11212 OUT_N.n300 OUT_N.n299 0.506
R11213 OUT_N.n399 OUT_N.n398 0.506
R11214 OUT_N.n498 OUT_N.n497 0.506
R11215 OUT_N.n665 OUT_N.n663 0.506
R11216 OUT_N.n754 OUT_N.n752 0.506
R11217 OUT_N.n853 OUT_N.n851 0.506
R11218 OUT_N.n952 OUT_N.n950 0.506
R11219 OUT_N.n313 OUT_N.n312 0.476
R11220 OUT_N.n412 OUT_N.n411 0.476
R11221 OUT_N.n511 OUT_N.n510 0.476
R11222 OUT_N.n651 OUT_N.n650 0.476
R11223 OUT_N.n740 OUT_N.n739 0.476
R11224 OUT_N.n839 OUT_N.n838 0.476
R11225 OUT_N.n938 OUT_N.n937 0.476
R11226 OUT_N.n1054 OUT_N.n1053 0.456
R11227 OUT_N.n1052 OUT_N.n1051 0.456
R11228 OUT_N.n217 OUT_N.n216 0.45
R11229 OUT_N.n180 OUT_N.n179 0.45
R11230 OUT_N.n143 OUT_N.n142 0.45
R11231 OUT_N.n640 OUT_N.n639 0.445
R11232 OUT_N.n729 OUT_N.n728 0.445
R11233 OUT_N.n828 OUT_N.n827 0.445
R11234 OUT_N.n927 OUT_N.n926 0.445
R11235 OUT_N.n268 OUT_N.n267 0.414
R11236 OUT_N.n367 OUT_N.n366 0.414
R11237 OUT_N.n466 OUT_N.n465 0.414
R11238 OUT_N.n582 OUT_N.n581 0.414
R11239 OUT_N.n681 OUT_N.n680 0.414
R11240 OUT_N.n780 OUT_N.n779 0.414
R11241 OUT_N.n879 OUT_N.n878 0.414
R11242 OUT_N.n278 OUT_N.n277 0.382
R11243 OUT_N.n377 OUT_N.n376 0.382
R11244 OUT_N.n476 OUT_N.n475 0.382
R11245 OUT_N.n593 OUT_N.n592 0.382
R11246 OUT_N.n692 OUT_N.n691 0.382
R11247 OUT_N.n791 OUT_N.n790 0.382
R11248 OUT_N.n890 OUT_N.n889 0.382
R11249 OUT_N.n554 OUT_N.n553 0.324
R11250 OUT_N.n1277 OUT_N.n1276 0.293
R11251 OUT_N.n1205 OUT_N.n1204 0.292
R11252 OUT_N.n1132 OUT_N.n1131 0.292
R11253 OUT_N.n1057 OUT_N.n1056 0.186
R11254 OUT_N.n874 OUT_N.n873 0.163
R11255 OUT_N.n775 OUT_N.n774 0.163
R11256 OUT_N.n676 OUT_N.n675 0.163
R11257 OUT_N.n455 OUT_N.n454 0.163
R11258 OUT_N.n356 OUT_N.n355 0.163
R11259 OUT_N.n1055 OUT_N.n1054 0.088
R11260 OUT_N.n1053 OUT_N.n1052 0.088
R11261 OUT_N.n310 OUT_N.n309 0.06
R11262 OUT_N.n261 OUT_N.n259 0.06
R11263 OUT_N.n272 OUT_N.n271 0.06
R11264 OUT_N.n289 OUT_N.n281 0.06
R11265 OUT_N.n409 OUT_N.n408 0.06
R11266 OUT_N.n360 OUT_N.n358 0.06
R11267 OUT_N.n371 OUT_N.n370 0.06
R11268 OUT_N.n388 OUT_N.n380 0.06
R11269 OUT_N.n508 OUT_N.n507 0.06
R11270 OUT_N.n459 OUT_N.n457 0.06
R11271 OUT_N.n470 OUT_N.n469 0.06
R11272 OUT_N.n487 OUT_N.n479 0.06
R11273 OUT_N.n596 OUT_N.n595 0.06
R11274 OUT_N.n586 OUT_N.n585 0.06
R11275 OUT_N.n637 OUT_N.n636 0.06
R11276 OUT_N.n648 OUT_N.n647 0.06
R11277 OUT_N.n695 OUT_N.n694 0.06
R11278 OUT_N.n685 OUT_N.n684 0.06
R11279 OUT_N.n726 OUT_N.n725 0.06
R11280 OUT_N.n737 OUT_N.n736 0.06
R11281 OUT_N.n794 OUT_N.n793 0.06
R11282 OUT_N.n784 OUT_N.n783 0.06
R11283 OUT_N.n825 OUT_N.n824 0.06
R11284 OUT_N.n836 OUT_N.n835 0.06
R11285 OUT_N.n893 OUT_N.n892 0.06
R11286 OUT_N.n883 OUT_N.n882 0.06
R11287 OUT_N.n924 OUT_N.n923 0.06
R11288 OUT_N.n935 OUT_N.n934 0.06
R11289 OUT_N.n226 OUT_N.n225 0.055
R11290 OUT_N.n189 OUT_N.n188 0.055
R11291 OUT_N.n152 OUT_N.n151 0.055
R11292 OUT_N.n120 OUT_N.n119 0.055
R11293 OUT_N.n323 OUT_N.n322 0.053
R11294 OUT_N.n322 OUT_N.n321 0.053
R11295 OUT_N.n422 OUT_N.n421 0.053
R11296 OUT_N.n421 OUT_N.n420 0.053
R11297 OUT_N.n521 OUT_N.n520 0.053
R11298 OUT_N.n520 OUT_N.n519 0.053
R11299 OUT_N.n666 OUT_N.n662 0.052
R11300 OUT_N.n626 OUT_N.n625 0.052
R11301 OUT_N.n755 OUT_N.n751 0.052
R11302 OUT_N.n761 OUT_N.n760 0.052
R11303 OUT_N.n854 OUT_N.n850 0.052
R11304 OUT_N.n860 OUT_N.n859 0.052
R11305 OUT_N.n953 OUT_N.n949 0.052
R11306 OUT_N.n959 OUT_N.n958 0.052
R11307 OUT_N.n1038 OUT_N.n1037 0.051
R11308 OUT_N.n1033 OUT_N.n1032 0.051
R11309 OUT_N.n1014 OUT_N.n1013 0.051
R11310 OUT_N.n1011 OUT_N.n1010 0.051
R11311 OUT_N.n988 OUT_N.n987 0.051
R11312 OUT_N.n985 OUT_N.n984 0.051
R11313 OUT_N.n243 OUT_N.n242 0.051
R11314 OUT_N.n240 OUT_N.n239 0.051
R11315 OUT_N.n206 OUT_N.n205 0.051
R11316 OUT_N.n203 OUT_N.n202 0.051
R11317 OUT_N.n169 OUT_N.n168 0.051
R11318 OUT_N.n166 OUT_N.n165 0.051
R11319 OUT_N.n137 OUT_N.n136 0.051
R11320 OUT_N.n134 OUT_N.n133 0.051
R11321 OUT_N.n1171 OUT_N.n1170 0.048
R11322 OUT_N.n1162 OUT_N.n1161 0.048
R11323 OUT_N.n1098 OUT_N.n1097 0.048
R11324 OUT_N.n1089 OUT_N.n1088 0.048
R11325 OUT_N.n661 OUT_N.n660 0.048
R11326 OUT_N.n750 OUT_N.n749 0.048
R11327 OUT_N.n849 OUT_N.n848 0.048
R11328 OUT_N.n948 OUT_N.n947 0.048
R11329 OUT_N.n93 OUT_N.n92 0.048
R11330 OUT_N.n85 OUT_N.n84 0.048
R11331 OUT_N.n58 OUT_N.n57 0.048
R11332 OUT_N.n50 OUT_N.n49 0.048
R11333 OUT_N.n23 OUT_N.n22 0.048
R11334 OUT_N.n15 OUT_N.n14 0.048
R11335 OUT_N.n1266 OUT_N.n1265 0.048
R11336 OUT_N.n1259 OUT_N.n1258 0.048
R11337 OUT_N.n1295 OUT_N.n1294 0.048
R11338 OUT_N.n1304 OUT_N.n1303 0.048
R11339 OUT_N.n595 OUT_N.n594 0.043
R11340 OUT_N.n694 OUT_N.n693 0.043
R11341 OUT_N.n793 OUT_N.n792 0.043
R11342 OUT_N.n892 OUT_N.n891 0.043
R11343 OUT_N.n1015 OUT_N.n1014 0.041
R11344 OUT_N.n989 OUT_N.n988 0.041
R11345 OUT_N.n1041 OUT_N.n1038 0.041
R11346 OUT_N.n314 OUT_N.n311 0.04
R11347 OUT_N.n413 OUT_N.n410 0.04
R11348 OUT_N.n512 OUT_N.n509 0.04
R11349 OUT_N.n1036 OUT_N.n1033 0.04
R11350 OUT_N.n1012 OUT_N.n1011 0.04
R11351 OUT_N.n986 OUT_N.n985 0.04
R11352 OUT_N.n652 OUT_N.n649 0.04
R11353 OUT_N.n741 OUT_N.n738 0.04
R11354 OUT_N.n840 OUT_N.n837 0.04
R11355 OUT_N.n939 OUT_N.n936 0.04
R11356 OUT_N.n241 OUT_N.n240 0.04
R11357 OUT_N.n247 OUT_N.n246 0.04
R11358 OUT_N.n204 OUT_N.n203 0.04
R11359 OUT_N.n210 OUT_N.n209 0.04
R11360 OUT_N.n167 OUT_N.n166 0.04
R11361 OUT_N.n173 OUT_N.n172 0.04
R11362 OUT_N.n135 OUT_N.n134 0.04
R11363 OUT_N.n115 OUT_N.n114 0.04
R11364 OUT_N.n244 OUT_N.n243 0.04
R11365 OUT_N.n207 OUT_N.n206 0.04
R11366 OUT_N.n170 OUT_N.n169 0.04
R11367 OUT_N.n138 OUT_N.n137 0.039
R11368 OUT_N.n1037 OUT_N.n1036 0.038
R11369 OUT_N.n1013 OUT_N.n1012 0.038
R11370 OUT_N.n987 OUT_N.n986 0.038
R11371 OUT_N.n242 OUT_N.n241 0.038
R11372 OUT_N.n248 OUT_N.n247 0.038
R11373 OUT_N.n205 OUT_N.n204 0.038
R11374 OUT_N.n211 OUT_N.n210 0.038
R11375 OUT_N.n168 OUT_N.n167 0.038
R11376 OUT_N.n174 OUT_N.n173 0.038
R11377 OUT_N.n136 OUT_N.n135 0.038
R11378 OUT_N.n114 OUT_N.n113 0.038
R11379 OUT_N.n1032 OUT_N.n1031 0.036
R11380 OUT_N.n1010 OUT_N.n1009 0.036
R11381 OUT_N.n984 OUT_N.n983 0.036
R11382 OUT_N.n585 OUT_N.n584 0.036
R11383 OUT_N.n684 OUT_N.n683 0.036
R11384 OUT_N.n783 OUT_N.n782 0.036
R11385 OUT_N.n882 OUT_N.n881 0.036
R11386 OUT_N.n249 OUT_N.n248 0.034
R11387 OUT_N.n212 OUT_N.n211 0.034
R11388 OUT_N.n175 OUT_N.n174 0.034
R11389 OUT_N.n1272 OUT_N.n1271 0.034
R11390 OUT_N.n113 OUT_N.n112 0.034
R11391 OUT_N.n239 OUT_N.n238 0.033
R11392 OUT_N.n202 OUT_N.n201 0.033
R11393 OUT_N.n165 OUT_N.n164 0.033
R11394 OUT_N.n1265 OUT_N.n1264 0.033
R11395 OUT_N.n133 OUT_N.n132 0.033
R11396 OUT_N.n116 OUT_N.n115 0.033
R11397 OUT_N.n1169 OUT_N.n1168 0.032
R11398 OUT_N.n1096 OUT_N.n1095 0.032
R11399 OUT_N.n92 OUT_N.n91 0.032
R11400 OUT_N.n57 OUT_N.n56 0.032
R11401 OUT_N.n22 OUT_N.n21 0.032
R11402 OUT_N.n1297 OUT_N.n1296 0.032
R11403 OUT_N.n1227 OUT_N.n1226 0.032
R11404 OUT_N.n32 OUT_N.n31 0.032
R11405 OUT_N.n67 OUT_N.n66 0.032
R11406 OUT_N.n102 OUT_N.n101 0.032
R11407 OUT_N.n1267 OUT_N.n1266 0.032
R11408 OUT_N.n318 OUT_N.n316 0.031
R11409 OUT_N.n307 OUT_N.n305 0.031
R11410 OUT_N.n271 OUT_N.n270 0.031
R11411 OUT_N.n288 OUT_N.n286 0.031
R11412 OUT_N.n417 OUT_N.n415 0.031
R11413 OUT_N.n406 OUT_N.n404 0.031
R11414 OUT_N.n370 OUT_N.n369 0.031
R11415 OUT_N.n387 OUT_N.n385 0.031
R11416 OUT_N.n516 OUT_N.n514 0.031
R11417 OUT_N.n505 OUT_N.n503 0.031
R11418 OUT_N.n469 OUT_N.n468 0.031
R11419 OUT_N.n486 OUT_N.n484 0.031
R11420 OUT_N.n645 OUT_N.n643 0.031
R11421 OUT_N.n656 OUT_N.n654 0.031
R11422 OUT_N.n734 OUT_N.n732 0.031
R11423 OUT_N.n745 OUT_N.n743 0.031
R11424 OUT_N.n833 OUT_N.n831 0.031
R11425 OUT_N.n844 OUT_N.n842 0.031
R11426 OUT_N.n932 OUT_N.n930 0.031
R11427 OUT_N.n943 OUT_N.n941 0.031
R11428 OUT_N.n96 OUT_N.n93 0.031
R11429 OUT_N.n61 OUT_N.n58 0.031
R11430 OUT_N.n26 OUT_N.n23 0.031
R11431 OUT_N.n235 OUT_N.n234 0.029
R11432 OUT_N.n198 OUT_N.n197 0.029
R11433 OUT_N.n161 OUT_N.n160 0.029
R11434 OUT_N.n129 OUT_N.n128 0.029
R11435 OUT_N.n1029 OUT_N.n1025 0.028
R11436 OUT_N.n1007 OUT_N.n1003 0.028
R11437 OUT_N.n981 OUT_N.n977 0.028
R11438 OUT_N.n1166 OUT_N.n1163 0.028
R11439 OUT_N.n1093 OUT_N.n1090 0.028
R11440 OUT_N.n1302 OUT_N.n1301 0.028
R11441 OUT_N.n1224 OUT_N.n1223 0.028
R11442 OUT_N.n31 OUT_N.n30 0.028
R11443 OUT_N.n1194 OUT_N.n1193 0.028
R11444 OUT_N.n66 OUT_N.n65 0.028
R11445 OUT_N.n1121 OUT_N.n1120 0.028
R11446 OUT_N.n101 OUT_N.n100 0.028
R11447 OUT_N.n118 OUT_N.n117 0.027
R11448 OUT_N.n251 OUT_N.n250 0.027
R11449 OUT_N.n214 OUT_N.n213 0.027
R11450 OUT_N.n177 OUT_N.n176 0.027
R11451 OUT_N.n1273 OUT_N.n1272 0.027
R11452 OUT_N.n259 OUT_N.n258 0.026
R11453 OUT_N.n266 OUT_N.n264 0.026
R11454 OUT_N.n276 OUT_N.n274 0.026
R11455 OUT_N.n358 OUT_N.n357 0.026
R11456 OUT_N.n365 OUT_N.n363 0.026
R11457 OUT_N.n375 OUT_N.n373 0.026
R11458 OUT_N.n457 OUT_N.n456 0.026
R11459 OUT_N.n464 OUT_N.n462 0.026
R11460 OUT_N.n474 OUT_N.n472 0.026
R11461 OUT_N.n590 OUT_N.n588 0.026
R11462 OUT_N.n634 OUT_N.n632 0.026
R11463 OUT_N.n638 OUT_N.n637 0.026
R11464 OUT_N.n641 OUT_N.n638 0.026
R11465 OUT_N.n689 OUT_N.n687 0.026
R11466 OUT_N.n723 OUT_N.n721 0.026
R11467 OUT_N.n727 OUT_N.n726 0.026
R11468 OUT_N.n730 OUT_N.n727 0.026
R11469 OUT_N.n788 OUT_N.n786 0.026
R11470 OUT_N.n822 OUT_N.n820 0.026
R11471 OUT_N.n826 OUT_N.n825 0.026
R11472 OUT_N.n829 OUT_N.n826 0.026
R11473 OUT_N.n887 OUT_N.n885 0.026
R11474 OUT_N.n921 OUT_N.n919 0.026
R11475 OUT_N.n925 OUT_N.n924 0.026
R11476 OUT_N.n928 OUT_N.n925 0.026
R11477 OUT_N.n1263 OUT_N.n1260 0.026
R11478 OUT_N.n1281 OUT_N.n1280 0.026
R11479 OUT_N.n1242 OUT_N.n1241 0.026
R11480 OUT_N.n1229 OUT_N.n1228 0.026
R11481 OUT_N.n1209 OUT_N.n1208 0.026
R11482 OUT_N.n1189 OUT_N.n1188 0.026
R11483 OUT_N.n1184 OUT_N.n1183 0.026
R11484 OUT_N.n1136 OUT_N.n1135 0.026
R11485 OUT_N.n1116 OUT_N.n1115 0.026
R11486 OUT_N.n1111 OUT_N.n1110 0.026
R11487 OUT_N.n1063 OUT_N.n1062 0.026
R11488 OUT_N.n89 OUT_N.n86 0.025
R11489 OUT_N.n223 OUT_N.n219 0.025
R11490 OUT_N.n54 OUT_N.n51 0.025
R11491 OUT_N.n186 OUT_N.n182 0.025
R11492 OUT_N.n19 OUT_N.n16 0.025
R11493 OUT_N.n149 OUT_N.n145 0.025
R11494 OUT_N.n1287 OUT_N.n1286 0.025
R11495 OUT_N.n35 OUT_N.n34 0.025
R11496 OUT_N.n1180 OUT_N.n1179 0.025
R11497 OUT_N.n70 OUT_N.n69 0.025
R11498 OUT_N.n1107 OUT_N.n1106 0.025
R11499 OUT_N.n105 OUT_N.n104 0.025
R11500 OUT_N.n289 OUT_N.n288 0.024
R11501 OUT_N.n388 OUT_N.n387 0.024
R11502 OUT_N.n487 OUT_N.n486 0.024
R11503 OUT_N.n599 OUT_N.n598 0.024
R11504 OUT_N.n598 OUT_N.n596 0.024
R11505 OUT_N.n698 OUT_N.n697 0.024
R11506 OUT_N.n697 OUT_N.n695 0.024
R11507 OUT_N.n797 OUT_N.n796 0.024
R11508 OUT_N.n796 OUT_N.n794 0.024
R11509 OUT_N.n896 OUT_N.n895 0.024
R11510 OUT_N.n895 OUT_N.n893 0.024
R11511 OUT_N.n335 OUT_N.n334 0.023
R11512 OUT_N.n434 OUT_N.n433 0.023
R11513 OUT_N.n533 OUT_N.n532 0.023
R11514 OUT_N.n613 OUT_N.n612 0.023
R11515 OUT_N.n616 OUT_N.n615 0.023
R11516 OUT_N.n712 OUT_N.n711 0.023
R11517 OUT_N.n715 OUT_N.n714 0.023
R11518 OUT_N.n811 OUT_N.n810 0.023
R11519 OUT_N.n814 OUT_N.n813 0.023
R11520 OUT_N.n910 OUT_N.n909 0.023
R11521 OUT_N.n913 OUT_N.n912 0.023
R11522 OUT_N.n1257 OUT_N.n1256 0.023
R11523 OUT_N.n1236 OUT_N.n1235 0.023
R11524 OUT_N.n766 OUT_N.n765 0.022
R11525 OUT_N.n865 OUT_N.n864 0.022
R11526 OUT_N.n964 OUT_N.n963 0.022
R11527 OUT_N.n328 OUT_N.n327 0.022
R11528 OUT_N.n427 OUT_N.n426 0.022
R11529 OUT_N.n526 OUT_N.n525 0.022
R11530 OUT_N.n74 OUT_N.n73 0.021
R11531 OUT_N.n39 OUT_N.n38 0.021
R11532 OUT_N.n4 OUT_N.n3 0.021
R11533 OUT_N.n324 OUT_N.n323 0.021
R11534 OUT_N.n280 OUT_N.n279 0.021
R11535 OUT_N.n281 OUT_N.n280 0.021
R11536 OUT_N.n423 OUT_N.n422 0.021
R11537 OUT_N.n379 OUT_N.n378 0.021
R11538 OUT_N.n380 OUT_N.n379 0.021
R11539 OUT_N.n522 OUT_N.n521 0.021
R11540 OUT_N.n478 OUT_N.n477 0.021
R11541 OUT_N.n479 OUT_N.n478 0.021
R11542 OUT_N.n1178 OUT_N.n1148 0.021
R11543 OUT_N.n1176 OUT_N.n1172 0.021
R11544 OUT_N.n1160 OUT_N.n1159 0.021
R11545 OUT_N.n1105 OUT_N.n1075 0.021
R11546 OUT_N.n1103 OUT_N.n1099 0.021
R11547 OUT_N.n1087 OUT_N.n1086 0.021
R11548 OUT_N.n83 OUT_N.n82 0.021
R11549 OUT_N.n48 OUT_N.n47 0.021
R11550 OUT_N.n13 OUT_N.n12 0.021
R11551 OUT_N.n1288 OUT_N.n1 0.021
R11552 OUT_N.n1293 OUT_N.n1292 0.021
R11553 OUT_N.n1311 OUT_N.n1310 0.021
R11554 OUT_N.n1287 OUT_N.n1219 0.021
R11555 OUT_N.n1309 OUT_N.n1308 0.021
R11556 OUT_N.n1215 OUT_N.n1214 0.021
R11557 OUT_N.n1179 OUT_N.n1146 0.021
R11558 OUT_N.n1200 OUT_N.n1199 0.021
R11559 OUT_N.n1142 OUT_N.n1141 0.021
R11560 OUT_N.n1106 OUT_N.n1073 0.021
R11561 OUT_N.n1127 OUT_N.n1126 0.021
R11562 OUT_N.n1069 OUT_N.n1068 0.021
R11563 OUT_N.n667 OUT_N.n630 0.021
R11564 OUT_N.n75 OUT_N.n74 0.021
R11565 OUT_N.n40 OUT_N.n39 0.021
R11566 OUT_N.n5 OUT_N.n4 0.021
R11567 OUT_N.n875 OUT_N.n874 0.02
R11568 OUT_N.n776 OUT_N.n775 0.02
R11569 OUT_N.n677 OUT_N.n676 0.02
R11570 OUT_N.n578 OUT_N.n577 0.02
R11571 OUT_N.n1238 OUT_N.n1237 0.02
R11572 OUT_N.n1057 OUT_N.n556 0.02
R11573 OUT_N.n550 OUT_N.n455 0.02
R11574 OUT_N.n451 OUT_N.n356 0.02
R11575 OUT_N.n352 OUT_N.n257 0.02
R11576 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN OUT_N.n668 0.019
R11577 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/DRAIN OUT_N.n767 0.019
R11578 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/DRAIN OUT_N.n866 0.019
R11579 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/DRAIN OUT_N.n965 0.019
R11580 OUT_N.n326 OUT_N.n324 0.019
R11581 OUT_N.n321 OUT_N.n320 0.019
R11582 OUT_N.n274 OUT_N.n272 0.019
R11583 OUT_N.n425 OUT_N.n423 0.019
R11584 OUT_N.n420 OUT_N.n419 0.019
R11585 OUT_N.n373 OUT_N.n371 0.019
R11586 OUT_N.n524 OUT_N.n522 0.019
R11587 OUT_N.n519 OUT_N.n518 0.019
R11588 OUT_N.n472 OUT_N.n470 0.019
R11589 OUT_N.n588 OUT_N.n586 0.019
R11590 OUT_N.n660 OUT_N.n658 0.019
R11591 OUT_N.n630 OUT_N.n629 0.019
R11592 OUT_N.n687 OUT_N.n685 0.019
R11593 OUT_N.n749 OUT_N.n747 0.019
R11594 OUT_N.n765 OUT_N.n764 0.019
R11595 OUT_N.n786 OUT_N.n784 0.019
R11596 OUT_N.n848 OUT_N.n846 0.019
R11597 OUT_N.n864 OUT_N.n863 0.019
R11598 OUT_N.n885 OUT_N.n883 0.019
R11599 OUT_N.n947 OUT_N.n945 0.019
R11600 OUT_N.n963 OUT_N.n962 0.019
R11601 OUT_N.n219 OUT_N.n218 0.018
R11602 OUT_N.n182 OUT_N.n181 0.018
R11603 OUT_N.n145 OUT_N.n144 0.018
R11604 OUT_N.n1232 OUT_N.n1231 0.018
R11605 OUT_N.n117 OUT_N.n116 0.018
R11606 OUT_N.n1023 OUT_N.n1022 0.017
R11607 OUT_N.n1020 OUT_N.n1019 0.017
R11608 OUT_N.n997 OUT_N.n996 0.017
R11609 OUT_N.n994 OUT_N.n993 0.017
R11610 OUT_N.n1249 OUT_N.n1248 0.017
R11611 OUT_N.n1049 OUT_N.n1048 0.017
R11612 OUT_N.n1046 OUT_N.n1045 0.017
R11613 OUT_N.n1222 OUT_N.n1221 0.017
R11614 OUT_N.n1213 OUT_N.n1212 0.017
R11615 OUT_N.n1216 OUT_N.n1215 0.017
R11616 OUT_N.n1196 OUT_N.n1195 0.017
R11617 OUT_N.n1140 OUT_N.n1139 0.017
R11618 OUT_N.n1143 OUT_N.n1142 0.017
R11619 OUT_N.n1123 OUT_N.n1122 0.017
R11620 OUT_N.n1067 OUT_N.n1066 0.017
R11621 OUT_N.n1070 OUT_N.n1069 0.017
R11622 OUT_N.n311 OUT_N.n310 0.016
R11623 OUT_N.n270 OUT_N.n269 0.016
R11624 OUT_N.n410 OUT_N.n409 0.016
R11625 OUT_N.n369 OUT_N.n368 0.016
R11626 OUT_N.n509 OUT_N.n508 0.016
R11627 OUT_N.n468 OUT_N.n467 0.016
R11628 OUT_N.n1152 OUT_N.n1151 0.016
R11629 OUT_N.n1079 OUT_N.n1078 0.016
R11630 OUT_N.n649 OUT_N.n648 0.016
R11631 OUT_N.n738 OUT_N.n737 0.016
R11632 OUT_N.n837 OUT_N.n836 0.016
R11633 OUT_N.n936 OUT_N.n935 0.016
R11634 OUT_N.n250 OUT_N.n249 0.016
R11635 OUT_N.n213 OUT_N.n212 0.016
R11636 OUT_N.n176 OUT_N.n175 0.016
R11637 OUT_N.n1269 OUT_N.n1268 0.016
R11638 OUT_N.n112 OUT_N.n111 0.016
R11639 OUT_N.n252 OUT_N.n226 0.016
R11640 OUT_N.n225 OUT_N.n224 0.016
R11641 OUT_N.n215 OUT_N.n189 0.016
R11642 OUT_N.n188 OUT_N.n187 0.016
R11643 OUT_N.n178 OUT_N.n152 0.016
R11644 OUT_N.n151 OUT_N.n150 0.016
R11645 OUT_N.n141 OUT_N.n120 0.016
R11646 OUT_N.n1319 OUT_N.n1318 0.016
R11647 OUT_N.n1219 OUT_N.n1218 0.016
R11648 OUT_N.n28 OUT_N.n27 0.016
R11649 OUT_N.n37 OUT_N.n36 0.016
R11650 OUT_N.n1146 OUT_N.n1145 0.016
R11651 OUT_N.n1202 OUT_N.n1201 0.016
R11652 OUT_N.n63 OUT_N.n62 0.016
R11653 OUT_N.n72 OUT_N.n71 0.016
R11654 OUT_N.n1073 OUT_N.n1072 0.016
R11655 OUT_N.n1129 OUT_N.n1128 0.016
R11656 OUT_N.n98 OUT_N.n97 0.016
R11657 OUT_N.n107 OUT_N.n106 0.016
R11658 OUT_N.n338 OUT_N.n337 0.015
R11659 OUT_N.n437 OUT_N.n436 0.015
R11660 OUT_N.n536 OUT_N.n535 0.015
R11661 OUT_N.n327 OUT_N.n326 0.014
R11662 OUT_N.n269 OUT_N.n266 0.014
R11663 OUT_N.n279 OUT_N.n276 0.014
R11664 OUT_N.n426 OUT_N.n425 0.014
R11665 OUT_N.n368 OUT_N.n365 0.014
R11666 OUT_N.n378 OUT_N.n375 0.014
R11667 OUT_N.n525 OUT_N.n524 0.014
R11668 OUT_N.n467 OUT_N.n464 0.014
R11669 OUT_N.n477 OUT_N.n474 0.014
R11670 OUT_N.n1025 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/GATE 0.014
R11671 OUT_N.n1172 OUT_N.n1171 0.014
R11672 OUT_N.n1150 OUT_N.n1149 0.014
R11673 OUT_N.n1003 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/GATE 0.014
R11674 OUT_N.n1021 OUT_N.n1020 0.014
R11675 OUT_N.n1099 OUT_N.n1098 0.014
R11676 OUT_N.n1077 OUT_N.n1076 0.014
R11677 OUT_N.n977 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/GATE 0.014
R11678 OUT_N.n995 OUT_N.n994 0.014
R11679 OUT_N.n636 OUT_N.n634 0.014
R11680 OUT_N.n725 OUT_N.n723 0.014
R11681 OUT_N.n824 OUT_N.n822 0.014
R11682 OUT_N.n923 OUT_N.n921 0.014
R11683 OUT_N.n972 OUT_N.n877 0.014
R11684 OUT_N.n873 OUT_N.n778 0.014
R11685 OUT_N.n774 OUT_N.n679 0.014
R11686 OUT_N.n675 OUT_N.n580 0.014
R11687 OUT_N.n82 OUT_N.n81 0.014
R11688 OUT_N.n47 OUT_N.n46 0.014
R11689 OUT_N.n12 OUT_N.n11 0.014
R11690 OUT_N.n1247 OUT_N.n1246 0.014
R11691 OUT_N.n1235 OUT_N.n1234 0.014
R11692 OUT_N.n1047 OUT_N.n1046 0.014
R11693 OUT_N.n1294 OUT_N.n1293 0.014
R11694 OUT_N.n1321 OUT_N.n1320 0.014
R11695 OUT_N.n1286 OUT_N.n1285 0.014
R11696 OUT_N.n1285 OUT_N.n1284 0.014
R11697 OUT_N.n1221 OUT_N.n1220 0.014
R11698 OUT_N.n1308 OUT_N.n1307 0.014
R11699 OUT_N.n1212 OUT_N.n37 0.014
R11700 OUT_N.n1181 OUT_N.n1180 0.014
R11701 OUT_N.n1185 OUT_N.n1181 0.014
R11702 OUT_N.n1202 OUT_N.n1196 0.014
R11703 OUT_N.n1199 OUT_N.n1198 0.014
R11704 OUT_N.n1139 OUT_N.n72 0.014
R11705 OUT_N.n1108 OUT_N.n1107 0.014
R11706 OUT_N.n1112 OUT_N.n1108 0.014
R11707 OUT_N.n1129 OUT_N.n1123 0.014
R11708 OUT_N.n1126 OUT_N.n1125 0.014
R11709 OUT_N.n1066 OUT_N.n107 0.014
R11710 OUT_N.n553 OUT_N.n552 0.014
R11711 OUT_N.n454 OUT_N.n453 0.014
R11712 OUT_N.n355 OUT_N.n354 0.014
R11713 OUT_N.n1022 OUT_N.n1021 0.013
R11714 OUT_N.n996 OUT_N.n995 0.013
R11715 OUT_N.n606 OUT_N.n605 0.013
R11716 OUT_N.n610 OUT_N.n609 0.013
R11717 OUT_N.n705 OUT_N.n704 0.013
R11718 OUT_N.n709 OUT_N.n708 0.013
R11719 OUT_N.n804 OUT_N.n803 0.013
R11720 OUT_N.n808 OUT_N.n807 0.013
R11721 OUT_N.n903 OUT_N.n902 0.013
R11722 OUT_N.n907 OUT_N.n906 0.013
R11723 OUT_N.n234 OUT_N 0.013
R11724 OUT_N.n197 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/GATE 0.013
R11725 OUT_N.n160 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE 0.013
R11726 OUT_N.n128 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE 0.013
R11727 OUT_N.n1048 OUT_N.n1047 0.013
R11728 OUT_N.n330 OUT_N.n329 0.012
R11729 OUT_N.n331 OUT_N.n330 0.012
R11730 OUT_N.n332 OUT_N.n331 0.012
R11731 OUT_N.n293 OUT_N.n292 0.012
R11732 OUT_N.n429 OUT_N.n428 0.012
R11733 OUT_N.n430 OUT_N.n429 0.012
R11734 OUT_N.n431 OUT_N.n430 0.012
R11735 OUT_N.n392 OUT_N.n391 0.012
R11736 OUT_N.n528 OUT_N.n527 0.012
R11737 OUT_N.n529 OUT_N.n528 0.012
R11738 OUT_N.n530 OUT_N.n529 0.012
R11739 OUT_N.n491 OUT_N.n490 0.012
R11740 OUT_N.n591 OUT_N.n590 0.012
R11741 OUT_N.n584 OUT_N.n583 0.012
R11742 OUT_N.n671 OUT_N.n670 0.012
R11743 OUT_N.n574 OUT_N.n573 0.012
R11744 OUT_N.n690 OUT_N.n689 0.012
R11745 OUT_N.n683 OUT_N.n682 0.012
R11746 OUT_N.n770 OUT_N.n769 0.012
R11747 OUT_N.n569 OUT_N.n568 0.012
R11748 OUT_N.n789 OUT_N.n788 0.012
R11749 OUT_N.n782 OUT_N.n781 0.012
R11750 OUT_N.n869 OUT_N.n868 0.012
R11751 OUT_N.n564 OUT_N.n563 0.012
R11752 OUT_N.n888 OUT_N.n887 0.012
R11753 OUT_N.n881 OUT_N.n880 0.012
R11754 OUT_N.n968 OUT_N.n967 0.012
R11755 OUT_N.n559 OUT_N.n558 0.012
R11756 OUT_N.n29 OUT_N.n28 0.012
R11757 OUT_N.n64 OUT_N.n63 0.012
R11758 OUT_N.n99 OUT_N.n98 0.012
R11759 OUT_N.n1282 OUT_N.n1281 0.011
R11760 OUT_N.n1274 OUT_N.n1269 0.011
R11761 OUT_N.n1274 OUT_N.n1273 0.011
R11762 OUT_N.n1238 OUT_N.n1232 0.011
R11763 OUT_N.n1206 OUT_N.n1205 0.011
R11764 OUT_N.n1208 OUT_N.n1207 0.011
R11765 OUT_N.n1188 OUT_N.n1187 0.011
R11766 OUT_N.n1133 OUT_N.n1132 0.011
R11767 OUT_N.n1135 OUT_N.n1134 0.011
R11768 OUT_N.n1115 OUT_N.n1114 0.011
R11769 OUT_N.n1060 OUT_N.n1059 0.011
R11770 OUT_N.n1062 OUT_N.n1061 0.011
R11771 OUT_N.n255 OUT_N.n254 0.011
R11772 OUT_N.n1008 OUT_N.n1007 0.011
R11773 OUT_N.n982 OUT_N.n981 0.011
R11774 OUT_N.n236 OUT_N.n235 0.011
R11775 OUT_N.n199 OUT_N.n198 0.011
R11776 OUT_N.n162 OUT_N.n161 0.011
R11777 OUT_N.n130 OUT_N.n129 0.011
R11778 OUT_N.n1030 OUT_N.n1029 0.011
R11779 OUT_N.n333 OUT_N.n332 0.01
R11780 OUT_N.n432 OUT_N.n431 0.01
R11781 OUT_N.n531 OUT_N.n530 0.01
R11782 OUT_N.n1159 OUT_N.n1158 0.01
R11783 OUT_N.n1154 OUT_N.n1152 0.01
R11784 OUT_N.n1086 OUT_N.n1085 0.01
R11785 OUT_N.n1081 OUT_N.n1079 0.01
R11786 OUT_N.n605 OUT_N.n604 0.01
R11787 OUT_N.n607 OUT_N.n606 0.01
R11788 OUT_N.n609 OUT_N.n608 0.01
R11789 OUT_N.n618 OUT_N.n617 0.01
R11790 OUT_N.n704 OUT_N.n703 0.01
R11791 OUT_N.n706 OUT_N.n705 0.01
R11792 OUT_N.n708 OUT_N.n707 0.01
R11793 OUT_N.n717 OUT_N.n716 0.01
R11794 OUT_N.n803 OUT_N.n802 0.01
R11795 OUT_N.n805 OUT_N.n804 0.01
R11796 OUT_N.n807 OUT_N.n806 0.01
R11797 OUT_N.n816 OUT_N.n815 0.01
R11798 OUT_N.n902 OUT_N.n901 0.01
R11799 OUT_N.n904 OUT_N.n903 0.01
R11800 OUT_N.n906 OUT_N.n905 0.01
R11801 OUT_N.n915 OUT_N.n914 0.01
R11802 OUT_N.n1256 OUT_N.n1255 0.01
R11803 OUT_N.n1276 OUT_N.n1275 0.01
R11804 OUT_N.n1243 OUT_N.n1242 0.01
R11805 OUT_N.n1241 OUT_N.n1240 0.01
R11806 OUT_N.n1315 OUT_N.n1311 0.01
R11807 OUT_N.n1318 OUT_N.n1317 0.01
R11808 OUT_N.n1307 OUT_N.n1306 0.01
R11809 OUT_N.n1198 OUT_N.n1197 0.01
R11810 OUT_N.n1125 OUT_N.n1124 0.01
R11811 OUT_N.n555 OUT_N.n554 0.01
R11812 OUT_N.n309 OUT_N.n307 0.009
R11813 OUT_N.n305 OUT_N.n304 0.009
R11814 OUT_N.n262 OUT_N.n261 0.009
R11815 OUT_N.n291 OUT_N.n290 0.009
R11816 OUT_N.n408 OUT_N.n406 0.009
R11817 OUT_N.n404 OUT_N.n403 0.009
R11818 OUT_N.n361 OUT_N.n360 0.009
R11819 OUT_N.n390 OUT_N.n389 0.009
R11820 OUT_N.n507 OUT_N.n505 0.009
R11821 OUT_N.n503 OUT_N.n502 0.009
R11822 OUT_N.n460 OUT_N.n459 0.009
R11823 OUT_N.n489 OUT_N.n488 0.009
R11824 OUT_N.n1024 OUT_N.n1023 0.009
R11825 OUT_N.n998 OUT_N.n997 0.009
R11826 OUT_N.n643 OUT_N.n641 0.009
R11827 OUT_N.n647 OUT_N.n645 0.009
R11828 OUT_N.n627 OUT_N.n626 0.009
R11829 OUT_N.n625 OUT_N.n624 0.009
R11830 OUT_N.n732 OUT_N.n730 0.009
R11831 OUT_N.n736 OUT_N.n734 0.009
R11832 OUT_N.n762 OUT_N.n761 0.009
R11833 OUT_N.n760 OUT_N.n759 0.009
R11834 OUT_N.n831 OUT_N.n829 0.009
R11835 OUT_N.n835 OUT_N.n833 0.009
R11836 OUT_N.n861 OUT_N.n860 0.009
R11837 OUT_N.n859 OUT_N.n858 0.009
R11838 OUT_N.n930 OUT_N.n928 0.009
R11839 OUT_N.n934 OUT_N.n932 0.009
R11840 OUT_N.n960 OUT_N.n959 0.009
R11841 OUT_N.n958 OUT_N.n957 0.009
R11842 OUT_N.n1280 OUT_N.n1279 0.009
R11843 OUT_N.n1278 OUT_N.n1277 0.009
R11844 OUT_N.n1231 OUT_N.n1230 0.009
R11845 OUT_N.n1234 OUT_N.n1233 0.009
R11846 OUT_N.n1050 OUT_N.n1049 0.009
R11847 OUT_N.n1210 OUT_N.n1209 0.009
R11848 OUT_N.n1190 OUT_N.n1189 0.009
R11849 OUT_N.n1204 OUT_N.n1203 0.009
R11850 OUT_N.n1137 OUT_N.n1136 0.009
R11851 OUT_N.n1117 OUT_N.n1116 0.009
R11852 OUT_N.n1131 OUT_N.n1130 0.009
R11853 OUT_N.n1064 OUT_N.n1063 0.009
R11854 OUT_N.n555 OUT_N.n256 0.009
R11855 OUT_N.n1058 OUT_N.n555 0.009
R11856 OUT_N.n336 OUT_N.n335 0.008
R11857 OUT_N.n344 OUT_N.n343 0.008
R11858 OUT_N.n348 OUT_N.n347 0.008
R11859 OUT_N.n435 OUT_N.n434 0.008
R11860 OUT_N.n443 OUT_N.n442 0.008
R11861 OUT_N.n447 OUT_N.n446 0.008
R11862 OUT_N.n534 OUT_N.n533 0.008
R11863 OUT_N.n542 OUT_N.n541 0.008
R11864 OUT_N.n546 OUT_N.n545 0.008
R11865 OUT_N.n1161 OUT_N.n1160 0.008
R11866 OUT_N.n1019 OUT_N.n1018 0.008
R11867 OUT_N.n1088 OUT_N.n1087 0.008
R11868 OUT_N.n993 OUT_N.n992 0.008
R11869 OUT_N.n611 OUT_N.n610 0.008
R11870 OUT_N.n615 OUT_N.n614 0.008
R11871 OUT_N.n619 OUT_N.n618 0.008
R11872 OUT_N.n674 OUT_N.n620 0.008
R11873 OUT_N.n710 OUT_N.n709 0.008
R11874 OUT_N.n714 OUT_N.n713 0.008
R11875 OUT_N.n718 OUT_N.n717 0.008
R11876 OUT_N.n773 OUT_N.n719 0.008
R11877 OUT_N.n809 OUT_N.n808 0.008
R11878 OUT_N.n813 OUT_N.n812 0.008
R11879 OUT_N.n817 OUT_N.n816 0.008
R11880 OUT_N.n872 OUT_N.n818 0.008
R11881 OUT_N.n908 OUT_N.n907 0.008
R11882 OUT_N.n912 OUT_N.n911 0.008
R11883 OUT_N.n916 OUT_N.n915 0.008
R11884 OUT_N.n971 OUT_N.n917 0.008
R11885 OUT_N.n86 OUT_N.n85 0.008
R11886 OUT_N.n51 OUT_N.n50 0.008
R11887 OUT_N.n16 OUT_N.n15 0.008
R11888 OUT_N.n1260 OUT_N.n1259 0.008
R11889 OUT_N.n1251 OUT_N.n1249 0.008
R11890 OUT_N.n1045 OUT_N.n1044 0.008
R11891 OUT_N.n1310 OUT_N.n1304 0.008
R11892 OUT_N.n1309 OUT_N.n1305 0.008
R11893 OUT_N.n36 OUT_N.n35 0.008
R11894 OUT_N.n1201 OUT_N.n1200 0.008
R11895 OUT_N.n71 OUT_N.n70 0.008
R11896 OUT_N.n1128 OUT_N.n1127 0.008
R11897 OUT_N.n106 OUT_N.n105 0.008
R11898 OUT_N.n286 OUT_N.n284 0.007
R11899 OUT_N.n339 OUT_N.n338 0.007
R11900 OUT_N.n340 OUT_N.n339 0.007
R11901 OUT_N.n385 OUT_N.n383 0.007
R11902 OUT_N.n438 OUT_N.n437 0.007
R11903 OUT_N.n439 OUT_N.n438 0.007
R11904 OUT_N.n484 OUT_N.n482 0.007
R11905 OUT_N.n537 OUT_N.n536 0.007
R11906 OUT_N.n538 OUT_N.n537 0.007
R11907 OUT_N.n1163 OUT_N.n1162 0.007
R11908 OUT_N.n1090 OUT_N.n1089 0.007
R11909 OUT_N.n601 OUT_N.n599 0.007
R11910 OUT_N.n662 OUT_N.n661 0.007
R11911 OUT_N.n700 OUT_N.n698 0.007
R11912 OUT_N.n751 OUT_N.n750 0.007
R11913 OUT_N.n799 OUT_N.n797 0.007
R11914 OUT_N.n850 OUT_N.n849 0.007
R11915 OUT_N.n898 OUT_N.n896 0.007
R11916 OUT_N.n949 OUT_N.n948 0.007
R11917 OUT_N.n90 OUT_N.n89 0.007
R11918 OUT_N.n84 OUT_N.n83 0.007
R11919 OUT_N.n77 OUT_N.n75 0.007
R11920 OUT_N.n251 OUT_N.n245 0.007
R11921 OUT_N.n223 OUT_N.n222 0.007
R11922 OUT_N.n55 OUT_N.n54 0.007
R11923 OUT_N.n49 OUT_N.n48 0.007
R11924 OUT_N.n42 OUT_N.n40 0.007
R11925 OUT_N.n214 OUT_N.n208 0.007
R11926 OUT_N.n186 OUT_N.n185 0.007
R11927 OUT_N.n20 OUT_N.n19 0.007
R11928 OUT_N.n14 OUT_N.n13 0.007
R11929 OUT_N.n7 OUT_N.n5 0.007
R11930 OUT_N.n177 OUT_N.n171 0.007
R11931 OUT_N.n149 OUT_N.n148 0.007
R11932 OUT_N.n1264 OUT_N.n1263 0.007
R11933 OUT_N.n1258 OUT_N.n1257 0.007
R11934 OUT_N.n1271 OUT_N.n1270 0.007
R11935 OUT_N.n1237 OUT_N.n1236 0.007
R11936 OUT_N.n140 OUT_N.n139 0.007
R11937 OUT_N.n1303 OUT_N.n1302 0.007
R11938 OUT_N.n1284 OUT_N.n1229 0.007
R11939 OUT_N.n1223 OUT_N.n1222 0.007
R11940 OUT_N.n30 OUT_N.n29 0.007
R11941 OUT_N.n34 OUT_N.n33 0.007
R11942 OUT_N.n1214 OUT_N.n1213 0.007
R11943 OUT_N.n1217 OUT_N.n1216 0.007
R11944 OUT_N.n1185 OUT_N.n1184 0.007
R11945 OUT_N.n1195 OUT_N.n1194 0.007
R11946 OUT_N.n65 OUT_N.n64 0.007
R11947 OUT_N.n69 OUT_N.n68 0.007
R11948 OUT_N.n1141 OUT_N.n1140 0.007
R11949 OUT_N.n1144 OUT_N.n1143 0.007
R11950 OUT_N.n1112 OUT_N.n1111 0.007
R11951 OUT_N.n1122 OUT_N.n1121 0.007
R11952 OUT_N.n100 OUT_N.n99 0.007
R11953 OUT_N.n104 OUT_N.n103 0.007
R11954 OUT_N.n1068 OUT_N.n1067 0.007
R11955 OUT_N.n1071 OUT_N.n1070 0.007
R11956 OUT_N.n549 OUT_N.n548 0.006
R11957 OUT_N.n450 OUT_N.n449 0.006
R11958 OUT_N.n351 OUT_N.n350 0.006
R11959 OUT_N.n965 OUT_N.n561 0.006
R11960 OUT_N.n866 OUT_N.n566 0.006
R11961 OUT_N.n767 OUT_N.n571 0.006
R11962 OUT_N.n668 OUT_N.n576 0.006
R11963 OUT_N.n351 OUT_N.n293 0.006
R11964 OUT_N.n450 OUT_N.n392 0.006
R11965 OUT_N.n549 OUT_N.n491 0.006
R11966 OUT_N.n337 OUT_N.n336 0.006
R11967 OUT_N.n347 OUT_N.n346 0.006
R11968 OUT_N.n436 OUT_N.n435 0.006
R11969 OUT_N.n446 OUT_N.n445 0.006
R11970 OUT_N.n535 OUT_N.n534 0.006
R11971 OUT_N.n545 OUT_N.n544 0.006
R11972 OUT_N.n612 OUT_N.n611 0.006
R11973 OUT_N.n614 OUT_N.n613 0.006
R11974 OUT_N.n711 OUT_N.n710 0.006
R11975 OUT_N.n713 OUT_N.n712 0.006
R11976 OUT_N.n810 OUT_N.n809 0.006
R11977 OUT_N.n812 OUT_N.n811 0.006
R11978 OUT_N.n909 OUT_N.n908 0.006
R11979 OUT_N.n911 OUT_N.n910 0.006
R11980 OUT_N.n256 OUT_N 0.006
R11981 OUT_N.n118 OUT_N.n110 0.006
R11982 OUT_N.n345 OUT_N.n344 0.005
R11983 OUT_N.n444 OUT_N.n443 0.005
R11984 OUT_N.n543 OUT_N.n542 0.005
R11985 OUT_N.n1148 OUT_N.n1147 0.005
R11986 OUT_N.n1151 OUT_N.n1150 0.005
R11987 OUT_N.n1149 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/GATE 0.005
R11988 OUT_N.n1075 OUT_N.n1074 0.005
R11989 OUT_N.n1078 OUT_N.n1077 0.005
R11990 OUT_N.n1076 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/GATE 0.005
R11991 OUT_N.n1248 OUT_N.n1247 0.005
R11992 OUT_N.n1246 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE 0.005
R11993 OUT_N.n1279 OUT_N.n1278 0.005
R11994 OUT_N.n1 OUT_N.n0 0.005
R11995 OUT_N.n1320 OUT_N.n1319 0.005
R11996 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/GATE OUT_N.n1321 0.005
R11997 OUT_N.n1211 OUT_N.n1210 0.005
R11998 OUT_N.n1203 OUT_N.n1190 0.005
R11999 OUT_N.n1138 OUT_N.n1137 0.005
R12000 OUT_N.n1130 OUT_N.n1117 0.005
R12001 OUT_N.n1065 OUT_N.n1064 0.005
R12002 OUT_N.n320 OUT_N.n318 0.004
R12003 OUT_N.n316 OUT_N.n314 0.004
R12004 OUT_N.n264 OUT_N.n262 0.004
R12005 OUT_N.n343 OUT_N.n342 0.004
R12006 OUT_N.n346 OUT_N.n345 0.004
R12007 OUT_N.n349 OUT_N.n348 0.004
R12008 OUT_N.n290 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/DRAIN 0.004
R12009 OUT_N.n419 OUT_N.n417 0.004
R12010 OUT_N.n415 OUT_N.n413 0.004
R12011 OUT_N.n363 OUT_N.n361 0.004
R12012 OUT_N.n442 OUT_N.n441 0.004
R12013 OUT_N.n445 OUT_N.n444 0.004
R12014 OUT_N.n448 OUT_N.n447 0.004
R12015 OUT_N.n389 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/DRAIN 0.004
R12016 OUT_N.n518 OUT_N.n516 0.004
R12017 OUT_N.n514 OUT_N.n512 0.004
R12018 OUT_N.n462 OUT_N.n460 0.004
R12019 OUT_N.n541 OUT_N.n540 0.004
R12020 OUT_N.n544 OUT_N.n543 0.004
R12021 OUT_N.n547 OUT_N.n546 0.004
R12022 OUT_N.n488 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/DRAIN 0.004
R12023 OUT_N.n654 OUT_N.n652 0.004
R12024 OUT_N.n658 OUT_N.n656 0.004
R12025 OUT_N.n629 OUT_N.n627 0.004
R12026 OUT_N.n620 OUT_N.n619 0.004
R12027 OUT_N.n670 OUT_N.n669 0.004
R12028 OUT_N.n743 OUT_N.n741 0.004
R12029 OUT_N.n747 OUT_N.n745 0.004
R12030 OUT_N.n764 OUT_N.n762 0.004
R12031 OUT_N.n719 OUT_N.n718 0.004
R12032 OUT_N.n769 OUT_N.n768 0.004
R12033 OUT_N.n842 OUT_N.n840 0.004
R12034 OUT_N.n846 OUT_N.n844 0.004
R12035 OUT_N.n863 OUT_N.n861 0.004
R12036 OUT_N.n818 OUT_N.n817 0.004
R12037 OUT_N.n868 OUT_N.n867 0.004
R12038 OUT_N.n941 OUT_N.n939 0.004
R12039 OUT_N.n945 OUT_N.n943 0.004
R12040 OUT_N.n962 OUT_N.n960 0.004
R12041 OUT_N.n917 OUT_N.n916 0.004
R12042 OUT_N.n967 OUT_N.n966 0.004
R12043 OUT_N.n1275 OUT_N.n1243 0.004
R12044 OUT_N.n1240 OUT_N.n1239 0.004
R12045 OUT_N.n877 OUT_N.n876 0.003
R12046 OUT_N.n778 OUT_N.n777 0.003
R12047 OUT_N.n679 OUT_N.n678 0.003
R12048 OUT_N.n580 OUT_N.n579 0.003
R12049 OUT_N.n579 OUT_N.n578 0.003
R12050 OUT_N.n876 OUT_N.n875 0.003
R12051 OUT_N.n777 OUT_N.n776 0.003
R12052 OUT_N.n678 OUT_N.n677 0.003
R12053 OUT_N.n552 OUT_N.n551 0.003
R12054 OUT_N.n453 OUT_N.n452 0.003
R12055 OUT_N.n354 OUT_N.n353 0.003
R12056 OUT_N.n551 OUT_N.n550 0.003
R12057 OUT_N.n452 OUT_N.n451 0.003
R12058 OUT_N.n353 OUT_N.n352 0.003
R12059 OUT_N.n603 OUT_N.n601 0.003
R12060 OUT_N.n702 OUT_N.n700 0.003
R12061 OUT_N.n801 OUT_N.n799 0.003
R12062 OUT_N.n900 OUT_N.n898 0.003
R12063 OUT_N.n334 OUT_N.n333 0.003
R12064 OUT_N.n433 OUT_N.n432 0.003
R12065 OUT_N.n532 OUT_N.n531 0.003
R12066 OUT_N.n1031 OUT_N.n1030 0.003
R12067 OUT_N.n1178 OUT_N.n1176 0.003
R12068 OUT_N.n1168 OUT_N.n1167 0.003
R12069 OUT_N.n1167 OUT_N.n1166 0.003
R12070 OUT_N.n1158 OUT_N.n1154 0.003
R12071 OUT_N.n1009 OUT_N.n1008 0.003
R12072 OUT_N.n1018 OUT_N.n1017 0.003
R12073 OUT_N.n1105 OUT_N.n1103 0.003
R12074 OUT_N.n1095 OUT_N.n1094 0.003
R12075 OUT_N.n1094 OUT_N.n1093 0.003
R12076 OUT_N.n1085 OUT_N.n1081 0.003
R12077 OUT_N.n983 OUT_N.n982 0.003
R12078 OUT_N.n992 OUT_N.n991 0.003
R12079 OUT_N.n617 OUT_N.n616 0.003
R12080 OUT_N.n716 OUT_N.n715 0.003
R12081 OUT_N.n815 OUT_N.n814 0.003
R12082 OUT_N.n914 OUT_N.n913 0.003
R12083 OUT_N.n91 OUT_N.n90 0.003
R12084 OUT_N.n81 OUT_N.n77 0.003
R12085 OUT_N.n238 OUT_N.n237 0.003
R12086 OUT_N.n237 OUT_N.n236 0.003
R12087 OUT_N.n222 OUT_N.n221 0.003
R12088 OUT_N.n221 OUT_N.n220 0.003
R12089 OUT_N.n56 OUT_N.n55 0.003
R12090 OUT_N.n46 OUT_N.n42 0.003
R12091 OUT_N.n201 OUT_N.n200 0.003
R12092 OUT_N.n200 OUT_N.n199 0.003
R12093 OUT_N.n185 OUT_N.n184 0.003
R12094 OUT_N.n184 OUT_N.n183 0.003
R12095 OUT_N.n21 OUT_N.n20 0.003
R12096 OUT_N.n11 OUT_N.n7 0.003
R12097 OUT_N.n164 OUT_N.n163 0.003
R12098 OUT_N.n163 OUT_N.n162 0.003
R12099 OUT_N.n148 OUT_N.n147 0.003
R12100 OUT_N.n147 OUT_N.n146 0.003
R12101 OUT_N.n1255 OUT_N.n1251 0.003
R12102 OUT_N.n132 OUT_N.n131 0.003
R12103 OUT_N.n131 OUT_N.n130 0.003
R12104 OUT_N.n110 OUT_N.n109 0.003
R12105 OUT_N.n109 OUT_N.n108 0.003
R12106 OUT_N.n1044 OUT_N.n1043 0.003
R12107 OUT_N.n1292 OUT_N.n1288 0.003
R12108 OUT_N.n1298 OUT_N.n1297 0.003
R12109 OUT_N.n1301 OUT_N.n1298 0.003
R12110 OUT_N.n1317 OUT_N.n1315 0.003
R12111 OUT_N.n1226 OUT_N.n1225 0.003
R12112 OUT_N.n1225 OUT_N.n1224 0.003
R12113 OUT_N.n33 OUT_N.n32 0.003
R12114 OUT_N.n1192 OUT_N.n1191 0.003
R12115 OUT_N.n1193 OUT_N.n1192 0.003
R12116 OUT_N.n68 OUT_N.n67 0.003
R12117 OUT_N.n1119 OUT_N.n1118 0.003
R12118 OUT_N.n1120 OUT_N.n1119 0.003
R12119 OUT_N.n103 OUT_N.n102 0.003
R12120 OUT_N.n284 OUT_N.n283 0.002
R12121 OUT_N.n383 OUT_N.n382 0.002
R12122 OUT_N.n482 OUT_N.n481 0.002
R12123 OUT_N.n594 OUT_N.n591 0.002
R12124 OUT_N.n608 OUT_N.n607 0.002
R12125 OUT_N.n573 OUT_N.n572 0.002
R12126 OUT_N.n575 OUT_N.n574 0.002
R12127 OUT_N.n693 OUT_N.n690 0.002
R12128 OUT_N.n707 OUT_N.n706 0.002
R12129 OUT_N.n568 OUT_N.n567 0.002
R12130 OUT_N.n570 OUT_N.n569 0.002
R12131 OUT_N.n792 OUT_N.n789 0.002
R12132 OUT_N.n806 OUT_N.n805 0.002
R12133 OUT_N.n563 OUT_N.n562 0.002
R12134 OUT_N.n565 OUT_N.n564 0.002
R12135 OUT_N.n891 OUT_N.n888 0.002
R12136 OUT_N.n905 OUT_N.n904 0.002
R12137 OUT_N.n558 OUT_N.n557 0.002
R12138 OUT_N.n560 OUT_N.n559 0.002
R12139 OUT_N.n1283 OUT_N.n1282 0.002
R12140 OUT_N.n253 OUT_N.n252 0.002
R12141 OUT_N.n224 OUT_N.n217 0.002
R12142 OUT_N.n216 OUT_N.n215 0.002
R12143 OUT_N.n187 OUT_N.n180 0.002
R12144 OUT_N.n179 OUT_N.n178 0.002
R12145 OUT_N.n150 OUT_N.n143 0.002
R12146 OUT_N.n142 OUT_N.n141 0.002
R12147 OUT_N.n1207 OUT_N.n1206 0.002
R12148 OUT_N.n1187 OUT_N.n1186 0.002
R12149 OUT_N.n1134 OUT_N.n1133 0.002
R12150 OUT_N.n1114 OUT_N.n1113 0.002
R12151 OUT_N.n1061 OUT_N.n1060 0.002
R12152 OUT_N.n766 OUT_N.n755 0.002
R12153 OUT_N.n865 OUT_N.n854 0.002
R12154 OUT_N.n964 OUT_N.n953 0.002
R12155 OUT_N.n341 OUT_N.n340 0.001
R12156 OUT_N.n440 OUT_N.n439 0.001
R12157 OUT_N.n539 OUT_N.n538 0.001
R12158 OUT_N.n673 OUT_N.n672 0.001
R12159 OUT_N.n772 OUT_N.n771 0.001
R12160 OUT_N.n871 OUT_N.n870 0.001
R12161 OUT_N.n970 OUT_N.n969 0.001
R12162 OUT_N.n971 OUT_N.n970 0.001
R12163 OUT_N.n872 OUT_N.n871 0.001
R12164 OUT_N.n773 OUT_N.n772 0.001
R12165 OUT_N.n674 OUT_N.n673 0.001
R12166 OUT_N.n540 OUT_N.n539 0.001
R12167 OUT_N.n441 OUT_N.n440 0.001
R12168 OUT_N.n342 OUT_N.n341 0.001
R12169 OUT_N.n350 OUT_N.n349 0.001
R12170 OUT_N.n292 OUT_N.n291 0.001
R12171 OUT_N.n449 OUT_N.n448 0.001
R12172 OUT_N.n391 OUT_N.n390 0.001
R12173 OUT_N.n548 OUT_N.n547 0.001
R12174 OUT_N.n490 OUT_N.n489 0.001
R12175 OUT_N.n1170 OUT_N.n1169 0.001
R12176 OUT_N.n1017 OUT_N.n1016 0.001
R12177 OUT_N.n1097 OUT_N.n1096 0.001
R12178 OUT_N.n991 OUT_N.n990 0.001
R12179 OUT_N.n672 OUT_N.n671 0.001
R12180 OUT_N.n576 OUT_N.n575 0.001
R12181 OUT_N.n771 OUT_N.n770 0.001
R12182 OUT_N.n571 OUT_N.n570 0.001
R12183 OUT_N.n870 OUT_N.n869 0.001
R12184 OUT_N.n566 OUT_N.n565 0.001
R12185 OUT_N.n969 OUT_N.n968 0.001
R12186 OUT_N.n561 OUT_N.n560 0.001
R12187 OUT_N.n73 OUT_N 0.001
R12188 OUT_N.n38 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/GATE 0.001
R12189 OUT_N.n3 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE 0.001
R12190 OUT_N.n1043 OUT_N.n1042 0.001
R12191 OUT_N.n1296 OUT_N.n1295 0.001
R12192 OUT_N.n1228 OUT_N.n1227 0.001
R12193 OUT_N.n1183 OUT_N.n1182 0.001
R12194 OUT_N.n1110 OUT_N.n1109 0.001
R12195 OUT_N.n667 OUT_N.n666 0.001
C0 OUT_N OUT_P 36.49fF
C1 OUT_P GND 51.63fF
C2 OUT_N GND 52.72fF
C3 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/GATE GND 0.00fF $ **FLOATING
C4 OUT_N.n0 GND 0.03fF $ **FLOATING
C5 OUT_N.n1 GND 0.01fF $ **FLOATING
C6 OUT_N.n2 GND 0.01fF $ **FLOATING
C7 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/GATE GND 0.00fF $ **FLOATING
C8 OUT_N.n3 GND 0.01fF $ **FLOATING
C9 OUT_N.n4 GND 0.02fF $ **FLOATING
C10 OUT_N.n5 GND 0.01fF $ **FLOATING
C11 OUT_N.n6 GND 0.01fF $ **FLOATING
C12 OUT_N.n7 GND 0.00fF $ **FLOATING
C13 OUT_N.t21 GND 0.25fF
C14 OUT_N.n8 GND 0.18fF $ **FLOATING
C15 OUT_N.n9 GND 0.03fF $ **FLOATING
C16 OUT_N.n10 GND 0.03fF $ **FLOATING
C17 OUT_N.n11 GND 0.01fF $ **FLOATING
C18 OUT_N.n12 GND 0.01fF $ **FLOATING
C19 OUT_N.n13 GND 0.01fF $ **FLOATING
C20 OUT_N.n14 GND 0.02fF $ **FLOATING
C21 OUT_N.n15 GND 0.02fF $ **FLOATING
C22 OUT_N.n16 GND 0.01fF $ **FLOATING
C23 OUT_N.n17 GND 0.05fF $ **FLOATING
C24 OUT_N.n18 GND 0.04fF $ **FLOATING
C25 OUT_N.n19 GND 0.01fF $ **FLOATING
C26 OUT_N.n20 GND 0.00fF $ **FLOATING
C27 OUT_N.n21 GND 0.01fF $ **FLOATING
C28 OUT_N.n22 GND 0.03fF $ **FLOATING
C29 OUT_N.n23 GND 0.03fF $ **FLOATING
C30 OUT_N.t17 GND 0.25fF
C31 OUT_N.n24 GND 0.18fF $ **FLOATING
C32 OUT_N.n25 GND 0.06fF $ **FLOATING
C33 OUT_N.n26 GND 0.07fF $ **FLOATING
C34 OUT_N.n27 GND 0.06fF $ **FLOATING
C35 OUT_N.n28 GND 0.01fF $ **FLOATING
C36 OUT_N.n29 GND 0.01fF $ **FLOATING
C37 OUT_N.n30 GND 0.01fF $ **FLOATING
C38 OUT_N.n31 GND 0.02fF $ **FLOATING
C39 OUT_N.n32 GND 0.01fF $ **FLOATING
C40 OUT_N.n33 GND 0.00fF $ **FLOATING
C41 OUT_N.n34 GND 0.01fF $ **FLOATING
C42 OUT_N.n35 GND 0.01fF $ **FLOATING
C43 OUT_N.n36 GND 0.01fF $ **FLOATING
C44 OUT_N.n37 GND 0.01fF $ **FLOATING
C45 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/GATE GND 0.00fF $ **FLOATING
C46 OUT_N.n38 GND 0.01fF $ **FLOATING
C47 OUT_N.n39 GND 0.02fF $ **FLOATING
C48 OUT_N.n40 GND 0.01fF $ **FLOATING
C49 OUT_N.n41 GND 0.01fF $ **FLOATING
C50 OUT_N.n42 GND 0.00fF $ **FLOATING
C51 OUT_N.t14 GND 0.25fF
C52 OUT_N.n43 GND 0.18fF $ **FLOATING
C53 OUT_N.n44 GND 0.03fF $ **FLOATING
C54 OUT_N.n45 GND 0.03fF $ **FLOATING
C55 OUT_N.n46 GND 0.01fF $ **FLOATING
C56 OUT_N.n47 GND 0.01fF $ **FLOATING
C57 OUT_N.n48 GND 0.01fF $ **FLOATING
C58 OUT_N.n49 GND 0.02fF $ **FLOATING
C59 OUT_N.n50 GND 0.02fF $ **FLOATING
C60 OUT_N.n51 GND 0.01fF $ **FLOATING
C61 OUT_N.n52 GND 0.05fF $ **FLOATING
C62 OUT_N.n53 GND 0.04fF $ **FLOATING
C63 OUT_N.n54 GND 0.01fF $ **FLOATING
C64 OUT_N.n55 GND 0.00fF $ **FLOATING
C65 OUT_N.n56 GND 0.01fF $ **FLOATING
C66 OUT_N.n57 GND 0.03fF $ **FLOATING
C67 OUT_N.n58 GND 0.03fF $ **FLOATING
C68 OUT_N.t15 GND 0.25fF
C69 OUT_N.n59 GND 0.18fF $ **FLOATING
C70 OUT_N.n60 GND 0.06fF $ **FLOATING
C71 OUT_N.n61 GND 0.07fF $ **FLOATING
C72 OUT_N.n62 GND 0.06fF $ **FLOATING
C73 OUT_N.n63 GND 0.01fF $ **FLOATING
C74 OUT_N.n64 GND 0.01fF $ **FLOATING
C75 OUT_N.n65 GND 0.01fF $ **FLOATING
C76 OUT_N.n66 GND 0.02fF $ **FLOATING
C77 OUT_N.n67 GND 0.01fF $ **FLOATING
C78 OUT_N.n68 GND 0.00fF $ **FLOATING
C79 OUT_N.n69 GND 0.01fF $ **FLOATING
C80 OUT_N.n70 GND 0.01fF $ **FLOATING
C81 OUT_N.n71 GND 0.01fF $ **FLOATING
C82 OUT_N.n72 GND 0.01fF $ **FLOATING
C83 OUT_N.n73 GND 0.01fF $ **FLOATING
C84 OUT_N.n74 GND 0.02fF $ **FLOATING
C85 OUT_N.n75 GND 0.01fF $ **FLOATING
C86 OUT_N.n76 GND 0.01fF $ **FLOATING
C87 OUT_N.n77 GND 0.00fF $ **FLOATING
C88 OUT_N.t18 GND 0.25fF
C89 OUT_N.n78 GND 0.18fF $ **FLOATING
C90 OUT_N.n79 GND 0.03fF $ **FLOATING
C91 OUT_N.n80 GND 0.03fF $ **FLOATING
C92 OUT_N.n81 GND 0.01fF $ **FLOATING
C93 OUT_N.n82 GND 0.01fF $ **FLOATING
C94 OUT_N.n83 GND 0.01fF $ **FLOATING
C95 OUT_N.n84 GND 0.02fF $ **FLOATING
C96 OUT_N.n85 GND 0.02fF $ **FLOATING
C97 OUT_N.n86 GND 0.01fF $ **FLOATING
C98 OUT_N.n87 GND 0.05fF $ **FLOATING
C99 OUT_N.n88 GND 0.04fF $ **FLOATING
C100 OUT_N.n89 GND 0.01fF $ **FLOATING
C101 OUT_N.n90 GND 0.00fF $ **FLOATING
C102 OUT_N.n91 GND 0.01fF $ **FLOATING
C103 OUT_N.n92 GND 0.03fF $ **FLOATING
C104 OUT_N.n93 GND 0.03fF $ **FLOATING
C105 OUT_N.t19 GND 0.25fF
C106 OUT_N.n94 GND 0.18fF $ **FLOATING
C107 OUT_N.n95 GND 0.06fF $ **FLOATING
C108 OUT_N.n96 GND 0.07fF $ **FLOATING
C109 OUT_N.n97 GND 0.06fF $ **FLOATING
C110 OUT_N.n98 GND 0.01fF $ **FLOATING
C111 OUT_N.n99 GND 0.01fF $ **FLOATING
C112 OUT_N.n100 GND 0.01fF $ **FLOATING
C113 OUT_N.n101 GND 0.02fF $ **FLOATING
C114 OUT_N.n102 GND 0.01fF $ **FLOATING
C115 OUT_N.n103 GND 0.00fF $ **FLOATING
C116 OUT_N.n104 GND 0.01fF $ **FLOATING
C117 OUT_N.n105 GND 0.01fF $ **FLOATING
C118 OUT_N.n106 GND 0.01fF $ **FLOATING
C119 OUT_N.n107 GND 0.01fF $ **FLOATING
C120 OUT_N.n108 GND 0.03fF $ **FLOATING
C121 OUT_N.n109 GND 0.00fF $ **FLOATING
C122 OUT_N.n110 GND 0.00fF $ **FLOATING
C123 OUT_N.n111 GND 0.01fF $ **FLOATING
C124 OUT_N.n112 GND 0.02fF $ **FLOATING
C125 OUT_N.n113 GND 0.02fF $ **FLOATING
C126 OUT_N.n114 GND 0.02fF $ **FLOATING
C127 OUT_N.n115 GND 0.02fF $ **FLOATING
C128 OUT_N.n116 GND 0.02fF $ **FLOATING
C129 OUT_N.n117 GND 0.01fF $ **FLOATING
C130 OUT_N.n118 GND 0.01fF $ **FLOATING
C131 OUT_N.n119 GND 0.11fF $ **FLOATING
C132 OUT_N.n120 GND 0.06fF $ **FLOATING
C133 OUT_N.n121 GND 0.18fF $ **FLOATING
C134 OUT_N.n122 GND 0.06fF $ **FLOATING
C135 OUT_N.n123 GND 0.05fF $ **FLOATING
C136 OUT_N.n124 GND 0.04fF $ **FLOATING
C137 OUT_N.n125 GND 0.18fF $ **FLOATING
C138 OUT_N.n126 GND 0.03fF $ **FLOATING
C139 OUT_N.n127 GND 0.04fF $ **FLOATING
C140 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/GATE GND 0.00fF $ **FLOATING
C141 OUT_N.n128 GND 0.02fF $ **FLOATING
C142 OUT_N.n129 GND 0.01fF $ **FLOATING
C143 OUT_N.n130 GND 0.01fF $ **FLOATING
C144 OUT_N.n131 GND 0.00fF $ **FLOATING
C145 OUT_N.n132 GND 0.01fF $ **FLOATING
C146 OUT_N.n133 GND 0.03fF $ **FLOATING
C147 OUT_N.n134 GND 0.03fF $ **FLOATING
C148 OUT_N.n135 GND 0.02fF $ **FLOATING
C149 OUT_N.n136 GND 0.03fF $ **FLOATING
C150 OUT_N.n137 GND 0.03fF $ **FLOATING
C151 OUT_N.n138 GND 0.06fF $ **FLOATING
C152 OUT_N.n139 GND 0.04fF $ **FLOATING
C153 OUT_N.n140 GND 0.01fF $ **FLOATING
C154 OUT_N.n141 GND 0.02fF $ **FLOATING
C155 OUT_N.n142 GND 0.36fF $ **FLOATING
C156 OUT_N.n143 GND 0.36fF $ **FLOATING
C157 OUT_N.n144 GND 0.02fF $ **FLOATING
C158 OUT_N.n145 GND 0.01fF $ **FLOATING
C159 OUT_N.n146 GND 0.03fF $ **FLOATING
C160 OUT_N.n147 GND 0.00fF $ **FLOATING
C161 OUT_N.n148 GND 0.00fF $ **FLOATING
C162 OUT_N.n149 GND 0.01fF $ **FLOATING
C163 OUT_N.n150 GND 0.02fF $ **FLOATING
C164 OUT_N.n151 GND 0.06fF $ **FLOATING
C165 OUT_N.n152 GND 0.06fF $ **FLOATING
C166 OUT_N.n153 GND 0.18fF $ **FLOATING
C167 OUT_N.n154 GND 0.06fF $ **FLOATING
C168 OUT_N.n155 GND 0.05fF $ **FLOATING
C169 OUT_N.n156 GND 0.04fF $ **FLOATING
C170 OUT_N.n157 GND 0.18fF $ **FLOATING
C171 OUT_N.n158 GND 0.03fF $ **FLOATING
C172 OUT_N.n159 GND 0.04fF $ **FLOATING
C173 OUT_N.n160 GND 0.02fF $ **FLOATING
C174 OUT_N.n161 GND 0.01fF $ **FLOATING
C175 OUT_N.n162 GND 0.01fF $ **FLOATING
C176 OUT_N.n163 GND 0.00fF $ **FLOATING
C177 OUT_N.n164 GND 0.01fF $ **FLOATING
C178 OUT_N.n165 GND 0.03fF $ **FLOATING
C179 OUT_N.n166 GND 0.03fF $ **FLOATING
C180 OUT_N.n167 GND 0.02fF $ **FLOATING
C181 OUT_N.n168 GND 0.03fF $ **FLOATING
C182 OUT_N.n169 GND 0.03fF $ **FLOATING
C183 OUT_N.n170 GND 0.06fF $ **FLOATING
C184 OUT_N.n171 GND 0.04fF $ **FLOATING
C185 OUT_N.n172 GND 0.02fF $ **FLOATING
C186 OUT_N.n173 GND 0.02fF $ **FLOATING
C187 OUT_N.n174 GND 0.02fF $ **FLOATING
C188 OUT_N.n175 GND 0.02fF $ **FLOATING
C189 OUT_N.n176 GND 0.01fF $ **FLOATING
C190 OUT_N.n177 GND 0.01fF $ **FLOATING
C191 OUT_N.n178 GND 0.02fF $ **FLOATING
C192 OUT_N.n179 GND 0.36fF $ **FLOATING
C193 OUT_N.n180 GND 0.36fF $ **FLOATING
C194 OUT_N.n181 GND 0.02fF $ **FLOATING
C195 OUT_N.n182 GND 0.01fF $ **FLOATING
C196 OUT_N.n183 GND 0.03fF $ **FLOATING
C197 OUT_N.n184 GND 0.00fF $ **FLOATING
C198 OUT_N.n185 GND 0.00fF $ **FLOATING
C199 OUT_N.n186 GND 0.01fF $ **FLOATING
C200 OUT_N.n187 GND 0.02fF $ **FLOATING
C201 OUT_N.n188 GND 0.06fF $ **FLOATING
C202 OUT_N.n189 GND 0.06fF $ **FLOATING
C203 OUT_N.n190 GND 0.18fF $ **FLOATING
C204 OUT_N.n191 GND 0.06fF $ **FLOATING
C205 OUT_N.n192 GND 0.05fF $ **FLOATING
C206 OUT_N.n193 GND 0.04fF $ **FLOATING
C207 OUT_N.n194 GND 0.18fF $ **FLOATING
C208 OUT_N.n195 GND 0.03fF $ **FLOATING
C209 OUT_N.n196 GND 0.04fF $ **FLOATING
C210 OUT_N.n197 GND 0.02fF $ **FLOATING
C211 OUT_N.n198 GND 0.01fF $ **FLOATING
C212 OUT_N.n199 GND 0.01fF $ **FLOATING
C213 OUT_N.n200 GND 0.00fF $ **FLOATING
C214 OUT_N.n201 GND 0.01fF $ **FLOATING
C215 OUT_N.n202 GND 0.03fF $ **FLOATING
C216 OUT_N.n203 GND 0.03fF $ **FLOATING
C217 OUT_N.n204 GND 0.02fF $ **FLOATING
C218 OUT_N.n205 GND 0.03fF $ **FLOATING
C219 OUT_N.n206 GND 0.03fF $ **FLOATING
C220 OUT_N.n207 GND 0.06fF $ **FLOATING
C221 OUT_N.n208 GND 0.04fF $ **FLOATING
C222 OUT_N.n209 GND 0.02fF $ **FLOATING
C223 OUT_N.n210 GND 0.02fF $ **FLOATING
C224 OUT_N.n211 GND 0.02fF $ **FLOATING
C225 OUT_N.n212 GND 0.02fF $ **FLOATING
C226 OUT_N.n213 GND 0.01fF $ **FLOATING
C227 OUT_N.n214 GND 0.01fF $ **FLOATING
C228 OUT_N.n215 GND 0.02fF $ **FLOATING
C229 OUT_N.n216 GND 0.36fF $ **FLOATING
C230 OUT_N.n217 GND 0.36fF $ **FLOATING
C231 OUT_N.n218 GND 0.02fF $ **FLOATING
C232 OUT_N.n219 GND 0.01fF $ **FLOATING
C233 OUT_N.n220 GND 0.03fF $ **FLOATING
C234 OUT_N.n221 GND 0.00fF $ **FLOATING
C235 OUT_N.n222 GND 0.00fF $ **FLOATING
C236 OUT_N.n223 GND 0.01fF $ **FLOATING
C237 OUT_N.n224 GND 0.02fF $ **FLOATING
C238 OUT_N.n225 GND 0.06fF $ **FLOATING
C239 OUT_N.n226 GND 0.06fF $ **FLOATING
C240 OUT_N.n227 GND 0.18fF $ **FLOATING
C241 OUT_N.n228 GND 0.06fF $ **FLOATING
C242 OUT_N.n229 GND 0.05fF $ **FLOATING
C243 OUT_N.n230 GND 0.04fF $ **FLOATING
C244 OUT_N.n231 GND 0.18fF $ **FLOATING
C245 OUT_N.n232 GND 0.03fF $ **FLOATING
C246 OUT_N.n233 GND 0.04fF $ **FLOATING
C247 OUT_N.n234 GND 0.02fF $ **FLOATING
C248 OUT_N.n235 GND 0.01fF $ **FLOATING
C249 OUT_N.n236 GND 0.01fF $ **FLOATING
C250 OUT_N.n237 GND 0.00fF $ **FLOATING
C251 OUT_N.n238 GND 0.01fF $ **FLOATING
C252 OUT_N.n239 GND 0.03fF $ **FLOATING
C253 OUT_N.n240 GND 0.03fF $ **FLOATING
C254 OUT_N.n241 GND 0.02fF $ **FLOATING
C255 OUT_N.n242 GND 0.03fF $ **FLOATING
C256 OUT_N.n243 GND 0.03fF $ **FLOATING
C257 OUT_N.n244 GND 0.06fF $ **FLOATING
C258 OUT_N.n245 GND 0.04fF $ **FLOATING
C259 OUT_N.n246 GND 0.02fF $ **FLOATING
C260 OUT_N.n247 GND 0.02fF $ **FLOATING
C261 OUT_N.n248 GND 0.02fF $ **FLOATING
C262 OUT_N.n249 GND 0.02fF $ **FLOATING
C263 OUT_N.n250 GND 0.01fF $ **FLOATING
C264 OUT_N.n251 GND 0.01fF $ **FLOATING
C265 OUT_N.n252 GND 0.02fF $ **FLOATING
C266 OUT_N.n253 GND 1.23fF $ **FLOATING
C267 OUT_N.n254 GND 3.01fF $ **FLOATING
C268 OUT_N.n256 GND 0.09fF $ **FLOATING
C269 OUT_N.n257 GND 1.35fF $ **FLOATING
C270 OUT_N.n258 GND 0.01fF $ **FLOATING
C271 OUT_N.n259 GND 0.02fF $ **FLOATING
C272 OUT_N.n260 GND 0.01fF $ **FLOATING
C273 OUT_N.n261 GND 0.01fF $ **FLOATING
C274 OUT_N.n262 GND 0.00fF $ **FLOATING
C275 OUT_N.n263 GND 0.00fF $ **FLOATING
C276 OUT_N.n264 GND 0.01fF $ **FLOATING
C277 OUT_N.n265 GND 0.00fF $ **FLOATING
C278 OUT_N.n266 GND 0.01fF $ **FLOATING
C279 OUT_N.n267 GND 0.01fF $ **FLOATING
C280 OUT_N.n268 GND 0.01fF $ **FLOATING
C281 OUT_N.n269 GND 0.01fF $ **FLOATING
C282 OUT_N.n270 GND 0.01fF $ **FLOATING
C283 OUT_N.n271 GND 0.02fF $ **FLOATING
C284 OUT_N.n272 GND 0.01fF $ **FLOATING
C285 OUT_N.n273 GND 0.02fF $ **FLOATING
C286 OUT_N.n274 GND 0.01fF $ **FLOATING
C287 OUT_N.n275 GND 0.00fF $ **FLOATING
C288 OUT_N.n276 GND 0.01fF $ **FLOATING
C289 OUT_N.n277 GND 0.01fF $ **FLOATING
C290 OUT_N.n278 GND 0.01fF $ **FLOATING
C291 OUT_N.n279 GND 0.01fF $ **FLOATING
C292 OUT_N.n280 GND 0.01fF $ **FLOATING
C293 OUT_N.n281 GND 0.01fF $ **FLOATING
C294 OUT_N.n282 GND 0.02fF $ **FLOATING
C295 OUT_N.n283 GND 0.02fF $ **FLOATING
C296 OUT_N.n284 GND 0.00fF $ **FLOATING
C297 OUT_N.n285 GND 0.00fF $ **FLOATING
C298 OUT_N.n286 GND 0.01fF $ **FLOATING
C299 OUT_N.n287 GND 0.02fF $ **FLOATING
C300 OUT_N.n288 GND 0.01fF $ **FLOATING
C301 OUT_N.n289 GND 0.01fF $ **FLOATING
C302 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/DRAIN GND 0.02fF $ **FLOATING
C303 OUT_N.n290 GND 0.05fF $ **FLOATING
C304 OUT_N.n291 GND 0.04fF $ **FLOATING
C305 OUT_N.n292 GND 0.05fF $ **FLOATING
C306 OUT_N.n293 GND 0.08fF $ **FLOATING
C307 OUT_N.t11 GND 0.23fF
C308 OUT_N.n294 GND 0.01fF $ **FLOATING
C309 OUT_N.t0 GND 0.23fF
C310 OUT_N.n295 GND 0.66fF $ **FLOATING
C311 OUT_N.n296 GND 0.09fF $ **FLOATING
C312 OUT_N.n297 GND 0.02fF $ **FLOATING
C313 OUT_N.n298 GND 0.00fF $ **FLOATING
C314 OUT_N.n299 GND 0.01fF $ **FLOATING
C315 OUT_N.n300 GND 0.01fF $ **FLOATING
C316 OUT_N.n301 GND 0.01fF $ **FLOATING
C317 OUT_N.n302 GND 0.00fF $ **FLOATING
C318 OUT_N.n303 GND 0.01fF $ **FLOATING
C319 OUT_N.n304 GND 0.01fF $ **FLOATING
C320 OUT_N.n305 GND 0.01fF $ **FLOATING
C321 OUT_N.n306 GND 0.00fF $ **FLOATING
C322 OUT_N.n307 GND 0.01fF $ **FLOATING
C323 OUT_N.n308 GND 0.01fF $ **FLOATING
C324 OUT_N.n309 GND 0.01fF $ **FLOATING
C325 OUT_N.n310 GND 0.01fF $ **FLOATING
C326 OUT_N.n311 GND 0.01fF $ **FLOATING
C327 OUT_N.n312 GND 0.01fF $ **FLOATING
C328 OUT_N.n313 GND 0.00fF $ **FLOATING
C329 OUT_N.n314 GND 0.01fF $ **FLOATING
C330 OUT_N.n315 GND 0.00fF $ **FLOATING
C331 OUT_N.n316 GND 0.01fF $ **FLOATING
C332 OUT_N.n317 GND 0.00fF $ **FLOATING
C333 OUT_N.n318 GND 0.01fF $ **FLOATING
C334 OUT_N.n319 GND 0.00fF $ **FLOATING
C335 OUT_N.n320 GND 0.00fF $ **FLOATING
C336 OUT_N.n321 GND 0.01fF $ **FLOATING
C337 OUT_N.n322 GND 0.02fF $ **FLOATING
C338 OUT_N.n323 GND 0.01fF $ **FLOATING
C339 OUT_N.n324 GND 0.01fF $ **FLOATING
C340 OUT_N.n325 GND 0.00fF $ **FLOATING
C341 OUT_N.n326 GND 0.01fF $ **FLOATING
C342 OUT_N.n327 GND 0.01fF $ **FLOATING
C343 OUT_N.n328 GND 0.51fF $ **FLOATING
C344 OUT_N.n329 GND 0.39fF $ **FLOATING
C345 OUT_N.n330 GND 0.08fF $ **FLOATING
C346 OUT_N.n331 GND 0.08fF $ **FLOATING
C347 OUT_N.n332 GND 0.08fF $ **FLOATING
C348 OUT_N.n333 GND 0.05fF $ **FLOATING
C349 OUT_N.n334 GND 0.09fF $ **FLOATING
C350 OUT_N.n335 GND 0.10fF $ **FLOATING
C351 OUT_N.n336 GND 0.05fF $ **FLOATING
C352 OUT_N.n337 GND 0.07fF $ **FLOATING
C353 OUT_N.n338 GND 0.08fF $ **FLOATING
C354 OUT_N.n339 GND 0.05fF $ **FLOATING
C355 OUT_N.n340 GND 0.03fF $ **FLOATING
C356 OUT_N.n342 GND 0.02fF $ **FLOATING
C357 OUT_N.n343 GND 0.04fF $ **FLOATING
C358 OUT_N.n344 GND 0.05fF $ **FLOATING
C359 OUT_N.n345 GND 0.03fF $ **FLOATING
C360 OUT_N.n346 GND 0.03fF $ **FLOATING
C361 OUT_N.n347 GND 0.05fF $ **FLOATING
C362 OUT_N.n348 GND 0.04fF $ **FLOATING
C363 OUT_N.n349 GND 0.02fF $ **FLOATING
C364 OUT_N.n350 GND 0.04fF $ **FLOATING
C365 OUT_N.n351 GND 0.01fF $ **FLOATING
C366 OUT_N.n352 GND 0.16fF $ **FLOATING
C367 OUT_N.n354 GND 0.12fF $ **FLOATING
C368 OUT_N.n355 GND 0.99fF $ **FLOATING
C369 OUT_N.n356 GND 1.02fF $ **FLOATING
C370 OUT_N.n357 GND 0.01fF $ **FLOATING
C371 OUT_N.n358 GND 0.02fF $ **FLOATING
C372 OUT_N.n359 GND 0.01fF $ **FLOATING
C373 OUT_N.n360 GND 0.01fF $ **FLOATING
C374 OUT_N.n361 GND 0.00fF $ **FLOATING
C375 OUT_N.n362 GND 0.00fF $ **FLOATING
C376 OUT_N.n363 GND 0.01fF $ **FLOATING
C377 OUT_N.n364 GND 0.00fF $ **FLOATING
C378 OUT_N.n365 GND 0.01fF $ **FLOATING
C379 OUT_N.n366 GND 0.01fF $ **FLOATING
C380 OUT_N.n367 GND 0.01fF $ **FLOATING
C381 OUT_N.n368 GND 0.01fF $ **FLOATING
C382 OUT_N.n369 GND 0.01fF $ **FLOATING
C383 OUT_N.n370 GND 0.02fF $ **FLOATING
C384 OUT_N.n371 GND 0.01fF $ **FLOATING
C385 OUT_N.n372 GND 0.02fF $ **FLOATING
C386 OUT_N.n373 GND 0.01fF $ **FLOATING
C387 OUT_N.n374 GND 0.00fF $ **FLOATING
C388 OUT_N.n375 GND 0.01fF $ **FLOATING
C389 OUT_N.n376 GND 0.01fF $ **FLOATING
C390 OUT_N.n377 GND 0.01fF $ **FLOATING
C391 OUT_N.n378 GND 0.01fF $ **FLOATING
C392 OUT_N.n379 GND 0.01fF $ **FLOATING
C393 OUT_N.n380 GND 0.01fF $ **FLOATING
C394 OUT_N.n381 GND 0.02fF $ **FLOATING
C395 OUT_N.n382 GND 0.02fF $ **FLOATING
C396 OUT_N.n383 GND 0.00fF $ **FLOATING
C397 OUT_N.n384 GND 0.00fF $ **FLOATING
C398 OUT_N.n385 GND 0.01fF $ **FLOATING
C399 OUT_N.n386 GND 0.02fF $ **FLOATING
C400 OUT_N.n387 GND 0.01fF $ **FLOATING
C401 OUT_N.n388 GND 0.01fF $ **FLOATING
C402 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/DRAIN GND 0.02fF $ **FLOATING
C403 OUT_N.n389 GND 0.05fF $ **FLOATING
C404 OUT_N.n390 GND 0.04fF $ **FLOATING
C405 OUT_N.n391 GND 0.05fF $ **FLOATING
C406 OUT_N.n392 GND 0.08fF $ **FLOATING
C407 OUT_N.t2 GND 0.23fF
C408 OUT_N.n393 GND 0.01fF $ **FLOATING
C409 OUT_N.t4 GND 0.23fF
C410 OUT_N.n394 GND 0.66fF $ **FLOATING
C411 OUT_N.n395 GND 0.09fF $ **FLOATING
C412 OUT_N.n396 GND 0.02fF $ **FLOATING
C413 OUT_N.n397 GND 0.00fF $ **FLOATING
C414 OUT_N.n398 GND 0.01fF $ **FLOATING
C415 OUT_N.n399 GND 0.01fF $ **FLOATING
C416 OUT_N.n400 GND 0.01fF $ **FLOATING
C417 OUT_N.n401 GND 0.00fF $ **FLOATING
C418 OUT_N.n402 GND 0.01fF $ **FLOATING
C419 OUT_N.n403 GND 0.01fF $ **FLOATING
C420 OUT_N.n404 GND 0.01fF $ **FLOATING
C421 OUT_N.n405 GND 0.00fF $ **FLOATING
C422 OUT_N.n406 GND 0.01fF $ **FLOATING
C423 OUT_N.n407 GND 0.01fF $ **FLOATING
C424 OUT_N.n408 GND 0.01fF $ **FLOATING
C425 OUT_N.n409 GND 0.01fF $ **FLOATING
C426 OUT_N.n410 GND 0.01fF $ **FLOATING
C427 OUT_N.n411 GND 0.01fF $ **FLOATING
C428 OUT_N.n412 GND 0.00fF $ **FLOATING
C429 OUT_N.n413 GND 0.01fF $ **FLOATING
C430 OUT_N.n414 GND 0.00fF $ **FLOATING
C431 OUT_N.n415 GND 0.01fF $ **FLOATING
C432 OUT_N.n416 GND 0.00fF $ **FLOATING
C433 OUT_N.n417 GND 0.01fF $ **FLOATING
C434 OUT_N.n418 GND 0.00fF $ **FLOATING
C435 OUT_N.n419 GND 0.00fF $ **FLOATING
C436 OUT_N.n420 GND 0.01fF $ **FLOATING
C437 OUT_N.n421 GND 0.02fF $ **FLOATING
C438 OUT_N.n422 GND 0.01fF $ **FLOATING
C439 OUT_N.n423 GND 0.01fF $ **FLOATING
C440 OUT_N.n424 GND 0.00fF $ **FLOATING
C441 OUT_N.n425 GND 0.01fF $ **FLOATING
C442 OUT_N.n426 GND 0.01fF $ **FLOATING
C443 OUT_N.n427 GND 0.51fF $ **FLOATING
C444 OUT_N.n428 GND 0.39fF $ **FLOATING
C445 OUT_N.n429 GND 0.08fF $ **FLOATING
C446 OUT_N.n430 GND 0.08fF $ **FLOATING
C447 OUT_N.n431 GND 0.08fF $ **FLOATING
C448 OUT_N.n432 GND 0.05fF $ **FLOATING
C449 OUT_N.n433 GND 0.09fF $ **FLOATING
C450 OUT_N.n434 GND 0.10fF $ **FLOATING
C451 OUT_N.n435 GND 0.05fF $ **FLOATING
C452 OUT_N.n436 GND 0.07fF $ **FLOATING
C453 OUT_N.n437 GND 0.08fF $ **FLOATING
C454 OUT_N.n438 GND 0.05fF $ **FLOATING
C455 OUT_N.n439 GND 0.03fF $ **FLOATING
C456 OUT_N.n441 GND 0.02fF $ **FLOATING
C457 OUT_N.n442 GND 0.04fF $ **FLOATING
C458 OUT_N.n443 GND 0.05fF $ **FLOATING
C459 OUT_N.n444 GND 0.03fF $ **FLOATING
C460 OUT_N.n445 GND 0.03fF $ **FLOATING
C461 OUT_N.n446 GND 0.05fF $ **FLOATING
C462 OUT_N.n447 GND 0.04fF $ **FLOATING
C463 OUT_N.n448 GND 0.02fF $ **FLOATING
C464 OUT_N.n449 GND 0.04fF $ **FLOATING
C465 OUT_N.n450 GND 0.01fF $ **FLOATING
C466 OUT_N.n451 GND 0.16fF $ **FLOATING
C467 OUT_N.n453 GND 0.12fF $ **FLOATING
C468 OUT_N.n454 GND 0.99fF $ **FLOATING
C469 OUT_N.n455 GND 1.02fF $ **FLOATING
C470 OUT_N.n456 GND 0.01fF $ **FLOATING
C471 OUT_N.n457 GND 0.02fF $ **FLOATING
C472 OUT_N.n458 GND 0.01fF $ **FLOATING
C473 OUT_N.n459 GND 0.01fF $ **FLOATING
C474 OUT_N.n460 GND 0.00fF $ **FLOATING
C475 OUT_N.n461 GND 0.00fF $ **FLOATING
C476 OUT_N.n462 GND 0.01fF $ **FLOATING
C477 OUT_N.n463 GND 0.00fF $ **FLOATING
C478 OUT_N.n464 GND 0.01fF $ **FLOATING
C479 OUT_N.n465 GND 0.01fF $ **FLOATING
C480 OUT_N.n466 GND 0.01fF $ **FLOATING
C481 OUT_N.n467 GND 0.01fF $ **FLOATING
C482 OUT_N.n468 GND 0.01fF $ **FLOATING
C483 OUT_N.n469 GND 0.02fF $ **FLOATING
C484 OUT_N.n470 GND 0.01fF $ **FLOATING
C485 OUT_N.n471 GND 0.02fF $ **FLOATING
C486 OUT_N.n472 GND 0.01fF $ **FLOATING
C487 OUT_N.n473 GND 0.00fF $ **FLOATING
C488 OUT_N.n474 GND 0.01fF $ **FLOATING
C489 OUT_N.n475 GND 0.01fF $ **FLOATING
C490 OUT_N.n476 GND 0.01fF $ **FLOATING
C491 OUT_N.n477 GND 0.01fF $ **FLOATING
C492 OUT_N.n478 GND 0.01fF $ **FLOATING
C493 OUT_N.n479 GND 0.01fF $ **FLOATING
C494 OUT_N.n480 GND 0.02fF $ **FLOATING
C495 OUT_N.n481 GND 0.02fF $ **FLOATING
C496 OUT_N.n482 GND 0.00fF $ **FLOATING
C497 OUT_N.n483 GND 0.00fF $ **FLOATING
C498 OUT_N.n484 GND 0.01fF $ **FLOATING
C499 OUT_N.n485 GND 0.02fF $ **FLOATING
C500 OUT_N.n486 GND 0.01fF $ **FLOATING
C501 OUT_N.n487 GND 0.01fF $ **FLOATING
C502 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/DRAIN GND 0.02fF $ **FLOATING
C503 OUT_N.n488 GND 0.05fF $ **FLOATING
C504 OUT_N.n489 GND 0.04fF $ **FLOATING
C505 OUT_N.n490 GND 0.05fF $ **FLOATING
C506 OUT_N.n491 GND 0.08fF $ **FLOATING
C507 OUT_N.t3 GND 0.23fF
C508 OUT_N.n492 GND 0.01fF $ **FLOATING
C509 OUT_N.t13 GND 0.23fF
C510 OUT_N.n493 GND 0.66fF $ **FLOATING
C511 OUT_N.n494 GND 0.09fF $ **FLOATING
C512 OUT_N.n495 GND 0.02fF $ **FLOATING
C513 OUT_N.n496 GND 0.00fF $ **FLOATING
C514 OUT_N.n497 GND 0.01fF $ **FLOATING
C515 OUT_N.n498 GND 0.01fF $ **FLOATING
C516 OUT_N.n499 GND 0.01fF $ **FLOATING
C517 OUT_N.n500 GND 0.00fF $ **FLOATING
C518 OUT_N.n501 GND 0.01fF $ **FLOATING
C519 OUT_N.n502 GND 0.01fF $ **FLOATING
C520 OUT_N.n503 GND 0.01fF $ **FLOATING
C521 OUT_N.n504 GND 0.00fF $ **FLOATING
C522 OUT_N.n505 GND 0.01fF $ **FLOATING
C523 OUT_N.n506 GND 0.01fF $ **FLOATING
C524 OUT_N.n507 GND 0.01fF $ **FLOATING
C525 OUT_N.n508 GND 0.01fF $ **FLOATING
C526 OUT_N.n509 GND 0.01fF $ **FLOATING
C527 OUT_N.n510 GND 0.01fF $ **FLOATING
C528 OUT_N.n511 GND 0.00fF $ **FLOATING
C529 OUT_N.n512 GND 0.01fF $ **FLOATING
C530 OUT_N.n513 GND 0.00fF $ **FLOATING
C531 OUT_N.n514 GND 0.01fF $ **FLOATING
C532 OUT_N.n515 GND 0.00fF $ **FLOATING
C533 OUT_N.n516 GND 0.01fF $ **FLOATING
C534 OUT_N.n517 GND 0.00fF $ **FLOATING
C535 OUT_N.n518 GND 0.00fF $ **FLOATING
C536 OUT_N.n519 GND 0.01fF $ **FLOATING
C537 OUT_N.n520 GND 0.02fF $ **FLOATING
C538 OUT_N.n521 GND 0.01fF $ **FLOATING
C539 OUT_N.n522 GND 0.01fF $ **FLOATING
C540 OUT_N.n523 GND 0.00fF $ **FLOATING
C541 OUT_N.n524 GND 0.01fF $ **FLOATING
C542 OUT_N.n525 GND 0.01fF $ **FLOATING
C543 OUT_N.n526 GND 0.51fF $ **FLOATING
C544 OUT_N.n527 GND 0.39fF $ **FLOATING
C545 OUT_N.n528 GND 0.08fF $ **FLOATING
C546 OUT_N.n529 GND 0.08fF $ **FLOATING
C547 OUT_N.n530 GND 0.08fF $ **FLOATING
C548 OUT_N.n531 GND 0.05fF $ **FLOATING
C549 OUT_N.n532 GND 0.09fF $ **FLOATING
C550 OUT_N.n533 GND 0.10fF $ **FLOATING
C551 OUT_N.n534 GND 0.05fF $ **FLOATING
C552 OUT_N.n535 GND 0.07fF $ **FLOATING
C553 OUT_N.n536 GND 0.08fF $ **FLOATING
C554 OUT_N.n537 GND 0.05fF $ **FLOATING
C555 OUT_N.n538 GND 0.03fF $ **FLOATING
C556 OUT_N.n540 GND 0.02fF $ **FLOATING
C557 OUT_N.n541 GND 0.04fF $ **FLOATING
C558 OUT_N.n542 GND 0.05fF $ **FLOATING
C559 OUT_N.n543 GND 0.03fF $ **FLOATING
C560 OUT_N.n544 GND 0.03fF $ **FLOATING
C561 OUT_N.n545 GND 0.05fF $ **FLOATING
C562 OUT_N.n546 GND 0.04fF $ **FLOATING
C563 OUT_N.n547 GND 0.02fF $ **FLOATING
C564 OUT_N.n548 GND 0.04fF $ **FLOATING
C565 OUT_N.n549 GND 0.01fF $ **FLOATING
C566 OUT_N.n550 GND 0.16fF $ **FLOATING
C567 OUT_N.n552 GND 0.12fF $ **FLOATING
C568 OUT_N.n553 GND 1.88fF $ **FLOATING
C569 OUT_N.n554 GND 1.86fF $ **FLOATING
C570 OUT_N.n555 GND 0.34fF $ **FLOATING
C571 OUT_N.n556 GND 0.23fF $ **FLOATING
C572 OUT_N.n557 GND 0.03fF $ **FLOATING
C573 OUT_N.n558 GND 0.05fF $ **FLOATING
C574 OUT_N.n559 GND 0.05fF $ **FLOATING
C575 OUT_N.n560 GND 0.01fF $ **FLOATING
C576 OUT_N.n561 GND 0.04fF $ **FLOATING
C577 OUT_N.n562 GND 0.03fF $ **FLOATING
C578 OUT_N.n563 GND 0.05fF $ **FLOATING
C579 OUT_N.n564 GND 0.05fF $ **FLOATING
C580 OUT_N.n565 GND 0.01fF $ **FLOATING
C581 OUT_N.n566 GND 0.04fF $ **FLOATING
C582 OUT_N.n567 GND 0.03fF $ **FLOATING
C583 OUT_N.n568 GND 0.05fF $ **FLOATING
C584 OUT_N.n569 GND 0.05fF $ **FLOATING
C585 OUT_N.n570 GND 0.01fF $ **FLOATING
C586 OUT_N.n571 GND 0.04fF $ **FLOATING
C587 OUT_N.n572 GND 0.03fF $ **FLOATING
C588 OUT_N.n573 GND 0.05fF $ **FLOATING
C589 OUT_N.n574 GND 0.05fF $ **FLOATING
C590 OUT_N.n575 GND 0.01fF $ **FLOATING
C591 OUT_N.n576 GND 0.04fF $ **FLOATING
C592 OUT_N.n577 GND 0.21fF $ **FLOATING
C593 OUT_N.n578 GND 0.16fF $ **FLOATING
C594 OUT_N.n580 GND 0.12fF $ **FLOATING
C595 OUT_N.n581 GND 0.01fF $ **FLOATING
C596 OUT_N.n582 GND 0.01fF $ **FLOATING
C597 OUT_N.n583 GND 0.00fF $ **FLOATING
C598 OUT_N.n584 GND 0.01fF $ **FLOATING
C599 OUT_N.n585 GND 0.02fF $ **FLOATING
C600 OUT_N.n586 GND 0.01fF $ **FLOATING
C601 OUT_N.n587 GND 0.02fF $ **FLOATING
C602 OUT_N.n588 GND 0.01fF $ **FLOATING
C603 OUT_N.n589 GND 0.00fF $ **FLOATING
C604 OUT_N.n590 GND 0.01fF $ **FLOATING
C605 OUT_N.n591 GND 0.00fF $ **FLOATING
C606 OUT_N.n592 GND 0.01fF $ **FLOATING
C607 OUT_N.n593 GND 0.01fF $ **FLOATING
C608 OUT_N.n594 GND 0.01fF $ **FLOATING
C609 OUT_N.n595 GND 0.02fF $ **FLOATING
C610 OUT_N.n596 GND 0.01fF $ **FLOATING
C611 OUT_N.n597 GND 0.02fF $ **FLOATING
C612 OUT_N.n598 GND 0.01fF $ **FLOATING
C613 OUT_N.n599 GND 0.01fF $ **FLOATING
C614 OUT_N.n600 GND 0.00fF $ **FLOATING
C615 OUT_N.n601 GND 0.00fF $ **FLOATING
C616 OUT_N.n602 GND 0.02fF $ **FLOATING
C617 OUT_N.n603 GND 0.02fF $ **FLOATING
C618 OUT_N.n604 GND 0.15fF $ **FLOATING
C619 OUT_N.n605 GND 0.08fF $ **FLOATING
C620 OUT_N.n606 GND 0.08fF $ **FLOATING
C621 OUT_N.n607 GND 0.04fF $ **FLOATING
C622 OUT_N.n608 GND 0.04fF $ **FLOATING
C623 OUT_N.n609 GND 0.08fF $ **FLOATING
C624 OUT_N.n610 GND 0.07fF $ **FLOATING
C625 OUT_N.n611 GND 0.05fF $ **FLOATING
C626 OUT_N.n612 GND 0.10fF $ **FLOATING
C627 OUT_N.n613 GND 0.10fF $ **FLOATING
C628 OUT_N.n614 GND 0.05fF $ **FLOATING
C629 OUT_N.n615 GND 0.10fF $ **FLOATING
C630 OUT_N.n616 GND 0.09fF $ **FLOATING
C631 OUT_N.n617 GND 0.05fF $ **FLOATING
C632 OUT_N.n618 GND 0.06fF $ **FLOATING
C633 OUT_N.n619 GND 0.04fF $ **FLOATING
C634 OUT_N.n620 GND 0.04fF $ **FLOATING
C635 OUT_N.n621 GND 0.02fF $ **FLOATING
C636 OUT_N.t6 GND 0.23fF
C637 OUT_N.t8 GND 0.23fF
C638 OUT_N.n622 GND 0.66fF $ **FLOATING
C639 OUT_N.n623 GND 0.07fF $ **FLOATING
C640 OUT_N.n624 GND 0.52fF $ **FLOATING
C641 OUT_N.n625 GND 0.01fF $ **FLOATING
C642 OUT_N.n626 GND 0.01fF $ **FLOATING
C643 OUT_N.n627 GND 0.00fF $ **FLOATING
C644 OUT_N.n628 GND 0.00fF $ **FLOATING
C645 OUT_N.n629 GND 0.00fF $ **FLOATING
C646 OUT_N.n630 GND 0.01fF $ **FLOATING
C647 OUT_N.n631 GND 0.00fF $ **FLOATING
C648 OUT_N.n632 GND 0.01fF $ **FLOATING
C649 OUT_N.n633 GND 0.00fF $ **FLOATING
C650 OUT_N.n634 GND 0.01fF $ **FLOATING
C651 OUT_N.n635 GND 0.01fF $ **FLOATING
C652 OUT_N.n636 GND 0.01fF $ **FLOATING
C653 OUT_N.n637 GND 0.02fF $ **FLOATING
C654 OUT_N.n638 GND 0.01fF $ **FLOATING
C655 OUT_N.n639 GND 0.01fF $ **FLOATING
C656 OUT_N.n640 GND 0.01fF $ **FLOATING
C657 OUT_N.n641 GND 0.01fF $ **FLOATING
C658 OUT_N.n642 GND 0.00fF $ **FLOATING
C659 OUT_N.n643 GND 0.01fF $ **FLOATING
C660 OUT_N.n644 GND 0.00fF $ **FLOATING
C661 OUT_N.n645 GND 0.01fF $ **FLOATING
C662 OUT_N.n646 GND 0.01fF $ **FLOATING
C663 OUT_N.n647 GND 0.01fF $ **FLOATING
C664 OUT_N.n648 GND 0.01fF $ **FLOATING
C665 OUT_N.n649 GND 0.01fF $ **FLOATING
C666 OUT_N.n650 GND 0.01fF $ **FLOATING
C667 OUT_N.n651 GND 0.00fF $ **FLOATING
C668 OUT_N.n652 GND 0.01fF $ **FLOATING
C669 OUT_N.n653 GND 0.00fF $ **FLOATING
C670 OUT_N.n654 GND 0.01fF $ **FLOATING
C671 OUT_N.n655 GND 0.00fF $ **FLOATING
C672 OUT_N.n656 GND 0.01fF $ **FLOATING
C673 OUT_N.n657 GND 0.00fF $ **FLOATING
C674 OUT_N.n658 GND 0.00fF $ **FLOATING
C675 OUT_N.n659 GND 0.01fF $ **FLOATING
C676 OUT_N.n660 GND 0.01fF $ **FLOATING
C677 OUT_N.n661 GND 0.01fF $ **FLOATING
C678 OUT_N.n662 GND 0.01fF $ **FLOATING
C679 OUT_N.n663 GND 0.01fF $ **FLOATING
C680 OUT_N.n664 GND 0.00fF $ **FLOATING
C681 OUT_N.n665 GND 0.01fF $ **FLOATING
C682 OUT_N.n666 GND 0.01fF $ **FLOATING
C683 OUT_N.n667 GND 0.00fF $ **FLOATING
C684 OUT_N.n668 GND 0.06fF $ **FLOATING
C685 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN GND 0.09fF $ **FLOATING
C686 OUT_N.n669 GND 0.05fF $ **FLOATING
C687 OUT_N.n670 GND 0.06fF $ **FLOATING
C688 OUT_N.n671 GND 0.05fF $ **FLOATING
C689 OUT_N.n672 GND 0.01fF $ **FLOATING
C690 OUT_N.n674 GND 0.04fF $ **FLOATING
C691 OUT_N.n675 GND 0.99fF $ **FLOATING
C692 OUT_N.n676 GND 1.02fF $ **FLOATING
C693 OUT_N.n677 GND 0.16fF $ **FLOATING
C694 OUT_N.n679 GND 0.12fF $ **FLOATING
C695 OUT_N.n680 GND 0.01fF $ **FLOATING
C696 OUT_N.n681 GND 0.01fF $ **FLOATING
C697 OUT_N.n682 GND 0.00fF $ **FLOATING
C698 OUT_N.n683 GND 0.01fF $ **FLOATING
C699 OUT_N.n684 GND 0.02fF $ **FLOATING
C700 OUT_N.n685 GND 0.01fF $ **FLOATING
C701 OUT_N.n686 GND 0.02fF $ **FLOATING
C702 OUT_N.n687 GND 0.01fF $ **FLOATING
C703 OUT_N.n688 GND 0.00fF $ **FLOATING
C704 OUT_N.n689 GND 0.01fF $ **FLOATING
C705 OUT_N.n690 GND 0.00fF $ **FLOATING
C706 OUT_N.n691 GND 0.01fF $ **FLOATING
C707 OUT_N.n692 GND 0.01fF $ **FLOATING
C708 OUT_N.n693 GND 0.01fF $ **FLOATING
C709 OUT_N.n694 GND 0.02fF $ **FLOATING
C710 OUT_N.n695 GND 0.01fF $ **FLOATING
C711 OUT_N.n696 GND 0.02fF $ **FLOATING
C712 OUT_N.n697 GND 0.01fF $ **FLOATING
C713 OUT_N.n698 GND 0.01fF $ **FLOATING
C714 OUT_N.n699 GND 0.00fF $ **FLOATING
C715 OUT_N.n700 GND 0.00fF $ **FLOATING
C716 OUT_N.n701 GND 0.02fF $ **FLOATING
C717 OUT_N.n702 GND 0.02fF $ **FLOATING
C718 OUT_N.n703 GND 0.15fF $ **FLOATING
C719 OUT_N.n704 GND 0.08fF $ **FLOATING
C720 OUT_N.n705 GND 0.08fF $ **FLOATING
C721 OUT_N.n706 GND 0.04fF $ **FLOATING
C722 OUT_N.n707 GND 0.04fF $ **FLOATING
C723 OUT_N.n708 GND 0.08fF $ **FLOATING
C724 OUT_N.n709 GND 0.07fF $ **FLOATING
C725 OUT_N.n710 GND 0.05fF $ **FLOATING
C726 OUT_N.n711 GND 0.10fF $ **FLOATING
C727 OUT_N.n712 GND 0.10fF $ **FLOATING
C728 OUT_N.n713 GND 0.05fF $ **FLOATING
C729 OUT_N.n714 GND 0.10fF $ **FLOATING
C730 OUT_N.n715 GND 0.09fF $ **FLOATING
C731 OUT_N.n716 GND 0.05fF $ **FLOATING
C732 OUT_N.n717 GND 0.06fF $ **FLOATING
C733 OUT_N.n718 GND 0.04fF $ **FLOATING
C734 OUT_N.n719 GND 0.04fF $ **FLOATING
C735 OUT_N.n720 GND 0.00fF $ **FLOATING
C736 OUT_N.n721 GND 0.01fF $ **FLOATING
C737 OUT_N.n722 GND 0.00fF $ **FLOATING
C738 OUT_N.n723 GND 0.01fF $ **FLOATING
C739 OUT_N.n724 GND 0.01fF $ **FLOATING
C740 OUT_N.n725 GND 0.01fF $ **FLOATING
C741 OUT_N.n726 GND 0.02fF $ **FLOATING
C742 OUT_N.n727 GND 0.01fF $ **FLOATING
C743 OUT_N.n728 GND 0.01fF $ **FLOATING
C744 OUT_N.n729 GND 0.01fF $ **FLOATING
C745 OUT_N.n730 GND 0.01fF $ **FLOATING
C746 OUT_N.n731 GND 0.00fF $ **FLOATING
C747 OUT_N.n732 GND 0.01fF $ **FLOATING
C748 OUT_N.n733 GND 0.00fF $ **FLOATING
C749 OUT_N.n734 GND 0.01fF $ **FLOATING
C750 OUT_N.n735 GND 0.01fF $ **FLOATING
C751 OUT_N.n736 GND 0.01fF $ **FLOATING
C752 OUT_N.n737 GND 0.01fF $ **FLOATING
C753 OUT_N.n738 GND 0.01fF $ **FLOATING
C754 OUT_N.n739 GND 0.01fF $ **FLOATING
C755 OUT_N.n740 GND 0.00fF $ **FLOATING
C756 OUT_N.n741 GND 0.01fF $ **FLOATING
C757 OUT_N.n742 GND 0.00fF $ **FLOATING
C758 OUT_N.n743 GND 0.01fF $ **FLOATING
C759 OUT_N.n744 GND 0.00fF $ **FLOATING
C760 OUT_N.n745 GND 0.01fF $ **FLOATING
C761 OUT_N.n746 GND 0.00fF $ **FLOATING
C762 OUT_N.n747 GND 0.00fF $ **FLOATING
C763 OUT_N.n748 GND 0.01fF $ **FLOATING
C764 OUT_N.n749 GND 0.01fF $ **FLOATING
C765 OUT_N.n750 GND 0.01fF $ **FLOATING
C766 OUT_N.n751 GND 0.01fF $ **FLOATING
C767 OUT_N.n752 GND 0.01fF $ **FLOATING
C768 OUT_N.n753 GND 0.00fF $ **FLOATING
C769 OUT_N.n754 GND 0.01fF $ **FLOATING
C770 OUT_N.n755 GND 0.01fF $ **FLOATING
C771 OUT_N.n756 GND 0.02fF $ **FLOATING
C772 OUT_N.t9 GND 0.23fF
C773 OUT_N.t12 GND 0.23fF
C774 OUT_N.n757 GND 0.66fF $ **FLOATING
C775 OUT_N.n758 GND 0.07fF $ **FLOATING
C776 OUT_N.n759 GND 0.52fF $ **FLOATING
C777 OUT_N.n760 GND 0.01fF $ **FLOATING
C778 OUT_N.n761 GND 0.01fF $ **FLOATING
C779 OUT_N.n762 GND 0.00fF $ **FLOATING
C780 OUT_N.n763 GND 0.00fF $ **FLOATING
C781 OUT_N.n764 GND 0.00fF $ **FLOATING
C782 OUT_N.n765 GND 0.01fF $ **FLOATING
C783 OUT_N.n766 GND 0.00fF $ **FLOATING
C784 OUT_N.n767 GND 0.06fF $ **FLOATING
C785 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/DRAIN GND 0.09fF $ **FLOATING
C786 OUT_N.n768 GND 0.05fF $ **FLOATING
C787 OUT_N.n769 GND 0.06fF $ **FLOATING
C788 OUT_N.n770 GND 0.05fF $ **FLOATING
C789 OUT_N.n771 GND 0.01fF $ **FLOATING
C790 OUT_N.n773 GND 0.04fF $ **FLOATING
C791 OUT_N.n774 GND 0.99fF $ **FLOATING
C792 OUT_N.n775 GND 1.02fF $ **FLOATING
C793 OUT_N.n776 GND 0.16fF $ **FLOATING
C794 OUT_N.n778 GND 0.12fF $ **FLOATING
C795 OUT_N.n779 GND 0.01fF $ **FLOATING
C796 OUT_N.n780 GND 0.01fF $ **FLOATING
C797 OUT_N.n781 GND 0.00fF $ **FLOATING
C798 OUT_N.n782 GND 0.01fF $ **FLOATING
C799 OUT_N.n783 GND 0.02fF $ **FLOATING
C800 OUT_N.n784 GND 0.01fF $ **FLOATING
C801 OUT_N.n785 GND 0.02fF $ **FLOATING
C802 OUT_N.n786 GND 0.01fF $ **FLOATING
C803 OUT_N.n787 GND 0.00fF $ **FLOATING
C804 OUT_N.n788 GND 0.01fF $ **FLOATING
C805 OUT_N.n789 GND 0.00fF $ **FLOATING
C806 OUT_N.n790 GND 0.01fF $ **FLOATING
C807 OUT_N.n791 GND 0.01fF $ **FLOATING
C808 OUT_N.n792 GND 0.01fF $ **FLOATING
C809 OUT_N.n793 GND 0.02fF $ **FLOATING
C810 OUT_N.n794 GND 0.01fF $ **FLOATING
C811 OUT_N.n795 GND 0.02fF $ **FLOATING
C812 OUT_N.n796 GND 0.01fF $ **FLOATING
C813 OUT_N.n797 GND 0.01fF $ **FLOATING
C814 OUT_N.n798 GND 0.00fF $ **FLOATING
C815 OUT_N.n799 GND 0.00fF $ **FLOATING
C816 OUT_N.n800 GND 0.02fF $ **FLOATING
C817 OUT_N.n801 GND 0.02fF $ **FLOATING
C818 OUT_N.n802 GND 0.15fF $ **FLOATING
C819 OUT_N.n803 GND 0.08fF $ **FLOATING
C820 OUT_N.n804 GND 0.08fF $ **FLOATING
C821 OUT_N.n805 GND 0.04fF $ **FLOATING
C822 OUT_N.n806 GND 0.04fF $ **FLOATING
C823 OUT_N.n807 GND 0.08fF $ **FLOATING
C824 OUT_N.n808 GND 0.07fF $ **FLOATING
C825 OUT_N.n809 GND 0.05fF $ **FLOATING
C826 OUT_N.n810 GND 0.10fF $ **FLOATING
C827 OUT_N.n811 GND 0.10fF $ **FLOATING
C828 OUT_N.n812 GND 0.05fF $ **FLOATING
C829 OUT_N.n813 GND 0.10fF $ **FLOATING
C830 OUT_N.n814 GND 0.09fF $ **FLOATING
C831 OUT_N.n815 GND 0.05fF $ **FLOATING
C832 OUT_N.n816 GND 0.06fF $ **FLOATING
C833 OUT_N.n817 GND 0.04fF $ **FLOATING
C834 OUT_N.n818 GND 0.04fF $ **FLOATING
C835 OUT_N.n819 GND 0.00fF $ **FLOATING
C836 OUT_N.n820 GND 0.01fF $ **FLOATING
C837 OUT_N.n821 GND 0.00fF $ **FLOATING
C838 OUT_N.n822 GND 0.01fF $ **FLOATING
C839 OUT_N.n823 GND 0.01fF $ **FLOATING
C840 OUT_N.n824 GND 0.01fF $ **FLOATING
C841 OUT_N.n825 GND 0.02fF $ **FLOATING
C842 OUT_N.n826 GND 0.01fF $ **FLOATING
C843 OUT_N.n827 GND 0.01fF $ **FLOATING
C844 OUT_N.n828 GND 0.01fF $ **FLOATING
C845 OUT_N.n829 GND 0.01fF $ **FLOATING
C846 OUT_N.n830 GND 0.00fF $ **FLOATING
C847 OUT_N.n831 GND 0.01fF $ **FLOATING
C848 OUT_N.n832 GND 0.00fF $ **FLOATING
C849 OUT_N.n833 GND 0.01fF $ **FLOATING
C850 OUT_N.n834 GND 0.01fF $ **FLOATING
C851 OUT_N.n835 GND 0.01fF $ **FLOATING
C852 OUT_N.n836 GND 0.01fF $ **FLOATING
C853 OUT_N.n837 GND 0.01fF $ **FLOATING
C854 OUT_N.n838 GND 0.01fF $ **FLOATING
C855 OUT_N.n839 GND 0.00fF $ **FLOATING
C856 OUT_N.n840 GND 0.01fF $ **FLOATING
C857 OUT_N.n841 GND 0.00fF $ **FLOATING
C858 OUT_N.n842 GND 0.01fF $ **FLOATING
C859 OUT_N.n843 GND 0.00fF $ **FLOATING
C860 OUT_N.n844 GND 0.01fF $ **FLOATING
C861 OUT_N.n845 GND 0.00fF $ **FLOATING
C862 OUT_N.n846 GND 0.00fF $ **FLOATING
C863 OUT_N.n847 GND 0.01fF $ **FLOATING
C864 OUT_N.n848 GND 0.01fF $ **FLOATING
C865 OUT_N.n849 GND 0.01fF $ **FLOATING
C866 OUT_N.n850 GND 0.01fF $ **FLOATING
C867 OUT_N.n851 GND 0.01fF $ **FLOATING
C868 OUT_N.n852 GND 0.00fF $ **FLOATING
C869 OUT_N.n853 GND 0.01fF $ **FLOATING
C870 OUT_N.n854 GND 0.01fF $ **FLOATING
C871 OUT_N.n855 GND 0.02fF $ **FLOATING
C872 OUT_N.t1 GND 0.23fF
C873 OUT_N.t7 GND 0.23fF
C874 OUT_N.n856 GND 0.66fF $ **FLOATING
C875 OUT_N.n857 GND 0.07fF $ **FLOATING
C876 OUT_N.n858 GND 0.52fF $ **FLOATING
C877 OUT_N.n859 GND 0.01fF $ **FLOATING
C878 OUT_N.n860 GND 0.01fF $ **FLOATING
C879 OUT_N.n861 GND 0.00fF $ **FLOATING
C880 OUT_N.n862 GND 0.00fF $ **FLOATING
C881 OUT_N.n863 GND 0.00fF $ **FLOATING
C882 OUT_N.n864 GND 0.01fF $ **FLOATING
C883 OUT_N.n865 GND 0.00fF $ **FLOATING
C884 OUT_N.n866 GND 0.06fF $ **FLOATING
C885 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/DRAIN GND 0.09fF $ **FLOATING
C886 OUT_N.n867 GND 0.05fF $ **FLOATING
C887 OUT_N.n868 GND 0.06fF $ **FLOATING
C888 OUT_N.n869 GND 0.05fF $ **FLOATING
C889 OUT_N.n870 GND 0.01fF $ **FLOATING
C890 OUT_N.n872 GND 0.04fF $ **FLOATING
C891 OUT_N.n873 GND 0.99fF $ **FLOATING
C892 OUT_N.n874 GND 1.02fF $ **FLOATING
C893 OUT_N.n875 GND 0.16fF $ **FLOATING
C894 OUT_N.n877 GND 0.12fF $ **FLOATING
C895 OUT_N.n878 GND 0.01fF $ **FLOATING
C896 OUT_N.n879 GND 0.01fF $ **FLOATING
C897 OUT_N.n880 GND 0.00fF $ **FLOATING
C898 OUT_N.n881 GND 0.01fF $ **FLOATING
C899 OUT_N.n882 GND 0.02fF $ **FLOATING
C900 OUT_N.n883 GND 0.01fF $ **FLOATING
C901 OUT_N.n884 GND 0.02fF $ **FLOATING
C902 OUT_N.n885 GND 0.01fF $ **FLOATING
C903 OUT_N.n886 GND 0.00fF $ **FLOATING
C904 OUT_N.n887 GND 0.01fF $ **FLOATING
C905 OUT_N.n888 GND 0.00fF $ **FLOATING
C906 OUT_N.n889 GND 0.01fF $ **FLOATING
C907 OUT_N.n890 GND 0.01fF $ **FLOATING
C908 OUT_N.n891 GND 0.01fF $ **FLOATING
C909 OUT_N.n892 GND 0.02fF $ **FLOATING
C910 OUT_N.n893 GND 0.01fF $ **FLOATING
C911 OUT_N.n894 GND 0.02fF $ **FLOATING
C912 OUT_N.n895 GND 0.01fF $ **FLOATING
C913 OUT_N.n896 GND 0.01fF $ **FLOATING
C914 OUT_N.n897 GND 0.00fF $ **FLOATING
C915 OUT_N.n898 GND 0.00fF $ **FLOATING
C916 OUT_N.n899 GND 0.02fF $ **FLOATING
C917 OUT_N.n900 GND 0.02fF $ **FLOATING
C918 OUT_N.n901 GND 0.15fF $ **FLOATING
C919 OUT_N.n902 GND 0.08fF $ **FLOATING
C920 OUT_N.n903 GND 0.08fF $ **FLOATING
C921 OUT_N.n904 GND 0.04fF $ **FLOATING
C922 OUT_N.n905 GND 0.04fF $ **FLOATING
C923 OUT_N.n906 GND 0.08fF $ **FLOATING
C924 OUT_N.n907 GND 0.07fF $ **FLOATING
C925 OUT_N.n908 GND 0.05fF $ **FLOATING
C926 OUT_N.n909 GND 0.10fF $ **FLOATING
C927 OUT_N.n910 GND 0.10fF $ **FLOATING
C928 OUT_N.n911 GND 0.05fF $ **FLOATING
C929 OUT_N.n912 GND 0.10fF $ **FLOATING
C930 OUT_N.n913 GND 0.09fF $ **FLOATING
C931 OUT_N.n914 GND 0.05fF $ **FLOATING
C932 OUT_N.n915 GND 0.06fF $ **FLOATING
C933 OUT_N.n916 GND 0.04fF $ **FLOATING
C934 OUT_N.n917 GND 0.04fF $ **FLOATING
C935 OUT_N.n918 GND 0.00fF $ **FLOATING
C936 OUT_N.n919 GND 0.01fF $ **FLOATING
C937 OUT_N.n920 GND 0.00fF $ **FLOATING
C938 OUT_N.n921 GND 0.01fF $ **FLOATING
C939 OUT_N.n922 GND 0.01fF $ **FLOATING
C940 OUT_N.n923 GND 0.01fF $ **FLOATING
C941 OUT_N.n924 GND 0.02fF $ **FLOATING
C942 OUT_N.n925 GND 0.01fF $ **FLOATING
C943 OUT_N.n926 GND 0.01fF $ **FLOATING
C944 OUT_N.n927 GND 0.01fF $ **FLOATING
C945 OUT_N.n928 GND 0.01fF $ **FLOATING
C946 OUT_N.n929 GND 0.00fF $ **FLOATING
C947 OUT_N.n930 GND 0.01fF $ **FLOATING
C948 OUT_N.n931 GND 0.00fF $ **FLOATING
C949 OUT_N.n932 GND 0.01fF $ **FLOATING
C950 OUT_N.n933 GND 0.01fF $ **FLOATING
C951 OUT_N.n934 GND 0.01fF $ **FLOATING
C952 OUT_N.n935 GND 0.01fF $ **FLOATING
C953 OUT_N.n936 GND 0.01fF $ **FLOATING
C954 OUT_N.n937 GND 0.01fF $ **FLOATING
C955 OUT_N.n938 GND 0.00fF $ **FLOATING
C956 OUT_N.n939 GND 0.01fF $ **FLOATING
C957 OUT_N.n940 GND 0.00fF $ **FLOATING
C958 OUT_N.n941 GND 0.01fF $ **FLOATING
C959 OUT_N.n942 GND 0.00fF $ **FLOATING
C960 OUT_N.n943 GND 0.01fF $ **FLOATING
C961 OUT_N.n944 GND 0.00fF $ **FLOATING
C962 OUT_N.n945 GND 0.00fF $ **FLOATING
C963 OUT_N.n946 GND 0.01fF $ **FLOATING
C964 OUT_N.n947 GND 0.01fF $ **FLOATING
C965 OUT_N.n948 GND 0.01fF $ **FLOATING
C966 OUT_N.n949 GND 0.01fF $ **FLOATING
C967 OUT_N.n950 GND 0.01fF $ **FLOATING
C968 OUT_N.n951 GND 0.00fF $ **FLOATING
C969 OUT_N.n952 GND 0.01fF $ **FLOATING
C970 OUT_N.n953 GND 0.01fF $ **FLOATING
C971 OUT_N.n954 GND 0.02fF $ **FLOATING
C972 OUT_N.t10 GND 0.23fF
C973 OUT_N.t5 GND 0.23fF
C974 OUT_N.n955 GND 0.66fF $ **FLOATING
C975 OUT_N.n956 GND 0.07fF $ **FLOATING
C976 OUT_N.n957 GND 0.52fF $ **FLOATING
C977 OUT_N.n958 GND 0.01fF $ **FLOATING
C978 OUT_N.n959 GND 0.01fF $ **FLOATING
C979 OUT_N.n960 GND 0.00fF $ **FLOATING
C980 OUT_N.n961 GND 0.00fF $ **FLOATING
C981 OUT_N.n962 GND 0.00fF $ **FLOATING
C982 OUT_N.n963 GND 0.01fF $ **FLOATING
C983 OUT_N.n964 GND 0.00fF $ **FLOATING
C984 OUT_N.n965 GND 0.06fF $ **FLOATING
C985 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/DRAIN GND 0.09fF $ **FLOATING
C986 OUT_N.n966 GND 0.05fF $ **FLOATING
C987 OUT_N.n967 GND 0.06fF $ **FLOATING
C988 OUT_N.n968 GND 0.05fF $ **FLOATING
C989 OUT_N.n969 GND 0.01fF $ **FLOATING
C990 OUT_N.n971 GND 0.04fF $ **FLOATING
C991 OUT_N.n972 GND 2.37fF $ **FLOATING
C992 OUT_N.n973 GND 0.18fF $ **FLOATING
C993 OUT_N.n974 GND 0.06fF $ **FLOATING
C994 OUT_N.n975 GND 0.05fF $ **FLOATING
C995 OUT_N.n976 GND 0.04fF $ **FLOATING
C996 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/GATE GND 0.00fF $ **FLOATING
C997 OUT_N.n977 GND 0.02fF $ **FLOATING
C998 OUT_N.n978 GND 0.18fF $ **FLOATING
C999 OUT_N.n979 GND 0.03fF $ **FLOATING
C1000 OUT_N.n980 GND 0.04fF $ **FLOATING
C1001 OUT_N.n981 GND 0.01fF $ **FLOATING
C1002 OUT_N.n982 GND 0.01fF $ **FLOATING
C1003 OUT_N.n983 GND 0.01fF $ **FLOATING
C1004 OUT_N.n984 GND 0.03fF $ **FLOATING
C1005 OUT_N.n985 GND 0.03fF $ **FLOATING
C1006 OUT_N.n986 GND 0.02fF $ **FLOATING
C1007 OUT_N.n987 GND 0.03fF $ **FLOATING
C1008 OUT_N.n988 GND 0.03fF $ **FLOATING
C1009 OUT_N.n989 GND 0.06fF $ **FLOATING
C1010 OUT_N.n990 GND 0.10fF $ **FLOATING
C1011 OUT_N.n991 GND 0.01fF $ **FLOATING
C1012 OUT_N.n992 GND 0.03fF $ **FLOATING
C1013 OUT_N.n993 GND 0.07fF $ **FLOATING
C1014 OUT_N.n994 GND 0.08fF $ **FLOATING
C1015 OUT_N.n995 GND 0.07fF $ **FLOATING
C1016 OUT_N.n996 GND 0.08fF $ **FLOATING
C1017 OUT_N.n997 GND 0.07fF $ **FLOATING
C1018 OUT_N.n998 GND 0.14fF $ **FLOATING
C1019 OUT_N.n999 GND 0.18fF $ **FLOATING
C1020 OUT_N.n1000 GND 0.06fF $ **FLOATING
C1021 OUT_N.n1001 GND 0.05fF $ **FLOATING
C1022 OUT_N.n1002 GND 0.04fF $ **FLOATING
C1023 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/GATE GND 0.00fF $ **FLOATING
C1024 OUT_N.n1003 GND 0.02fF $ **FLOATING
C1025 OUT_N.n1004 GND 0.18fF $ **FLOATING
C1026 OUT_N.n1005 GND 0.03fF $ **FLOATING
C1027 OUT_N.n1006 GND 0.04fF $ **FLOATING
C1028 OUT_N.n1007 GND 0.01fF $ **FLOATING
C1029 OUT_N.n1008 GND 0.01fF $ **FLOATING
C1030 OUT_N.n1009 GND 0.01fF $ **FLOATING
C1031 OUT_N.n1010 GND 0.03fF $ **FLOATING
C1032 OUT_N.n1011 GND 0.03fF $ **FLOATING
C1033 OUT_N.n1012 GND 0.02fF $ **FLOATING
C1034 OUT_N.n1013 GND 0.03fF $ **FLOATING
C1035 OUT_N.n1014 GND 0.03fF $ **FLOATING
C1036 OUT_N.n1015 GND 0.06fF $ **FLOATING
C1037 OUT_N.n1016 GND 0.10fF $ **FLOATING
C1038 OUT_N.n1017 GND 0.01fF $ **FLOATING
C1039 OUT_N.n1018 GND 0.03fF $ **FLOATING
C1040 OUT_N.n1019 GND 0.07fF $ **FLOATING
C1041 OUT_N.n1020 GND 0.08fF $ **FLOATING
C1042 OUT_N.n1021 GND 0.07fF $ **FLOATING
C1043 OUT_N.n1022 GND 0.08fF $ **FLOATING
C1044 OUT_N.n1023 GND 0.07fF $ **FLOATING
C1045 OUT_N.n1024 GND 0.14fF $ **FLOATING
C1046 OUT_N.n1025 GND 0.02fF $ **FLOATING
C1047 OUT_N.n1026 GND 0.18fF $ **FLOATING
C1048 OUT_N.n1027 GND 0.03fF $ **FLOATING
C1049 OUT_N.n1028 GND 0.04fF $ **FLOATING
C1050 OUT_N.n1029 GND 0.01fF $ **FLOATING
C1051 OUT_N.n1030 GND 0.01fF $ **FLOATING
C1052 OUT_N.n1031 GND 0.01fF $ **FLOATING
C1053 OUT_N.n1032 GND 0.03fF $ **FLOATING
C1054 OUT_N.n1033 GND 0.03fF $ **FLOATING
C1055 OUT_N.n1034 GND 0.05fF $ **FLOATING
C1056 OUT_N.n1035 GND 0.04fF $ **FLOATING
C1057 OUT_N.n1036 GND 0.02fF $ **FLOATING
C1058 OUT_N.n1037 GND 0.03fF $ **FLOATING
C1059 OUT_N.n1038 GND 0.03fF $ **FLOATING
C1060 OUT_N.n1039 GND 0.18fF $ **FLOATING
C1061 OUT_N.n1040 GND 0.06fF $ **FLOATING
C1062 OUT_N.n1041 GND 0.06fF $ **FLOATING
C1063 OUT_N.n1042 GND 0.10fF $ **FLOATING
C1064 OUT_N.n1043 GND 0.01fF $ **FLOATING
C1065 OUT_N.n1044 GND 0.04fF $ **FLOATING
C1066 OUT_N.n1045 GND 0.07fF $ **FLOATING
C1067 OUT_N.n1046 GND 0.08fF $ **FLOATING
C1068 OUT_N.n1047 GND 0.07fF $ **FLOATING
C1069 OUT_N.n1048 GND 0.08fF $ **FLOATING
C1070 OUT_N.n1049 GND 0.07fF $ **FLOATING
C1071 OUT_N.n1050 GND 0.14fF $ **FLOATING
C1072 OUT_N.n1051 GND 0.54fF $ **FLOATING
C1073 OUT_N.n1052 GND 0.43fF $ **FLOATING
C1074 OUT_N.n1053 GND 0.43fF $ **FLOATING
C1075 OUT_N.n1054 GND 0.43fF $ **FLOATING
C1076 OUT_N.n1055 GND 1.44fF $ **FLOATING
C1077 OUT_N.n1056 GND 4.52fF $ **FLOATING
C1078 OUT_N.n1057 GND 1.16fF $ **FLOATING
C1079 OUT_N.n1058 GND 0.57fF $ **FLOATING
C1080 OUT_N.n1059 GND 0.48fF $ **FLOATING
C1081 OUT_N.n1060 GND 0.01fF $ **FLOATING
C1082 OUT_N.n1061 GND 0.01fF $ **FLOATING
C1083 OUT_N.n1062 GND 0.03fF $ **FLOATING
C1084 OUT_N.n1063 GND 0.03fF $ **FLOATING
C1085 OUT_N.n1064 GND 0.01fF $ **FLOATING
C1086 OUT_N.n1065 GND 0.07fF $ **FLOATING
C1087 OUT_N.n1066 GND 0.01fF $ **FLOATING
C1088 OUT_N.n1067 GND 0.01fF $ **FLOATING
C1089 OUT_N.n1068 GND 0.01fF $ **FLOATING
C1090 OUT_N.n1069 GND 0.01fF $ **FLOATING
C1091 OUT_N.n1070 GND 0.01fF $ **FLOATING
C1092 OUT_N.n1071 GND 0.22fF $ **FLOATING
C1093 OUT_N.n1072 GND 0.23fF $ **FLOATING
C1094 OUT_N.n1073 GND 0.01fF $ **FLOATING
C1095 OUT_N.n1074 GND 0.03fF $ **FLOATING
C1096 OUT_N.n1075 GND 0.01fF $ **FLOATING
C1097 OUT_N.n1076 GND 0.01fF $ **FLOATING
C1098 OUT_N.n1077 GND 0.01fF $ **FLOATING
C1099 OUT_N.n1078 GND 0.01fF $ **FLOATING
C1100 OUT_N.n1079 GND 0.01fF $ **FLOATING
C1101 OUT_N.n1080 GND 0.01fF $ **FLOATING
C1102 OUT_N.n1081 GND 0.00fF $ **FLOATING
C1103 OUT_N.t25 GND 0.25fF
C1104 OUT_N.n1082 GND 0.18fF $ **FLOATING
C1105 OUT_N.n1083 GND 0.03fF $ **FLOATING
C1106 OUT_N.n1084 GND 0.03fF $ **FLOATING
C1107 OUT_N.n1085 GND 0.00fF $ **FLOATING
C1108 OUT_N.n1086 GND 0.01fF $ **FLOATING
C1109 OUT_N.n1087 GND 0.01fF $ **FLOATING
C1110 OUT_N.n1088 GND 0.02fF $ **FLOATING
C1111 OUT_N.n1089 GND 0.02fF $ **FLOATING
C1112 OUT_N.n1090 GND 0.01fF $ **FLOATING
C1113 OUT_N.n1091 GND 0.05fF $ **FLOATING
C1114 OUT_N.n1092 GND 0.04fF $ **FLOATING
C1115 OUT_N.n1093 GND 0.01fF $ **FLOATING
C1116 OUT_N.n1094 GND 0.00fF $ **FLOATING
C1117 OUT_N.n1095 GND 0.01fF $ **FLOATING
C1118 OUT_N.n1096 GND 0.01fF $ **FLOATING
C1119 OUT_N.n1097 GND 0.02fF $ **FLOATING
C1120 OUT_N.n1098 GND 0.02fF $ **FLOATING
C1121 OUT_N.n1099 GND 0.01fF $ **FLOATING
C1122 OUT_N.t27 GND 0.25fF
C1123 OUT_N.n1100 GND 0.18fF $ **FLOATING
C1124 OUT_N.n1101 GND 0.03fF $ **FLOATING
C1125 OUT_N.n1102 GND 0.03fF $ **FLOATING
C1126 OUT_N.n1103 GND 0.01fF $ **FLOATING
C1127 OUT_N.n1104 GND 0.01fF $ **FLOATING
C1128 OUT_N.n1105 GND 0.01fF $ **FLOATING
C1129 OUT_N.n1106 GND 0.01fF $ **FLOATING
C1130 OUT_N.n1107 GND 0.01fF $ **FLOATING
C1131 OUT_N.n1108 GND 0.01fF $ **FLOATING
C1132 OUT_N.n1109 GND 0.01fF $ **FLOATING
C1133 OUT_N.n1110 GND 0.01fF $ **FLOATING
C1134 OUT_N.n1111 GND 0.01fF $ **FLOATING
C1135 OUT_N.n1112 GND 0.01fF $ **FLOATING
C1136 OUT_N.n1113 GND 0.07fF $ **FLOATING
C1137 OUT_N.n1114 GND 0.01fF $ **FLOATING
C1138 OUT_N.n1115 GND 0.03fF $ **FLOATING
C1139 OUT_N.n1116 GND 0.03fF $ **FLOATING
C1140 OUT_N.n1117 GND 0.01fF $ **FLOATING
C1141 OUT_N.n1118 GND 0.01fF $ **FLOATING
C1142 OUT_N.n1119 GND 0.00fF $ **FLOATING
C1143 OUT_N.n1120 GND 0.01fF $ **FLOATING
C1144 OUT_N.n1121 GND 0.01fF $ **FLOATING
C1145 OUT_N.n1122 GND 0.01fF $ **FLOATING
C1146 OUT_N.n1123 GND 0.01fF $ **FLOATING
C1147 OUT_N.n1124 GND 0.03fF $ **FLOATING
C1148 OUT_N.n1125 GND 0.01fF $ **FLOATING
C1149 OUT_N.n1126 GND 0.01fF $ **FLOATING
C1150 OUT_N.n1127 GND 0.01fF $ **FLOATING
C1151 OUT_N.n1128 GND 0.01fF $ **FLOATING
C1152 OUT_N.n1129 GND 0.01fF $ **FLOATING
C1153 OUT_N.n1130 GND 0.01fF $ **FLOATING
C1154 OUT_N.n1131 GND 0.26fF $ **FLOATING
C1155 OUT_N.n1132 GND 0.26fF $ **FLOATING
C1156 OUT_N.n1133 GND 0.01fF $ **FLOATING
C1157 OUT_N.n1134 GND 0.01fF $ **FLOATING
C1158 OUT_N.n1135 GND 0.03fF $ **FLOATING
C1159 OUT_N.n1136 GND 0.03fF $ **FLOATING
C1160 OUT_N.n1137 GND 0.01fF $ **FLOATING
C1161 OUT_N.n1138 GND 0.07fF $ **FLOATING
C1162 OUT_N.n1139 GND 0.01fF $ **FLOATING
C1163 OUT_N.n1140 GND 0.01fF $ **FLOATING
C1164 OUT_N.n1141 GND 0.01fF $ **FLOATING
C1165 OUT_N.n1142 GND 0.01fF $ **FLOATING
C1166 OUT_N.n1143 GND 0.01fF $ **FLOATING
C1167 OUT_N.n1144 GND 0.22fF $ **FLOATING
C1168 OUT_N.n1145 GND 0.23fF $ **FLOATING
C1169 OUT_N.n1146 GND 0.01fF $ **FLOATING
C1170 OUT_N.n1147 GND 0.03fF $ **FLOATING
C1171 OUT_N.n1148 GND 0.01fF $ **FLOATING
C1172 OUT_N.n1149 GND 0.01fF $ **FLOATING
C1173 OUT_N.n1150 GND 0.01fF $ **FLOATING
C1174 OUT_N.n1151 GND 0.01fF $ **FLOATING
C1175 OUT_N.n1152 GND 0.01fF $ **FLOATING
C1176 OUT_N.n1153 GND 0.01fF $ **FLOATING
C1177 OUT_N.n1154 GND 0.00fF $ **FLOATING
C1178 OUT_N.t23 GND 0.25fF
C1179 OUT_N.n1155 GND 0.18fF $ **FLOATING
C1180 OUT_N.n1156 GND 0.03fF $ **FLOATING
C1181 OUT_N.n1157 GND 0.03fF $ **FLOATING
C1182 OUT_N.n1158 GND 0.00fF $ **FLOATING
C1183 OUT_N.n1159 GND 0.01fF $ **FLOATING
C1184 OUT_N.n1160 GND 0.01fF $ **FLOATING
C1185 OUT_N.n1161 GND 0.02fF $ **FLOATING
C1186 OUT_N.n1162 GND 0.02fF $ **FLOATING
C1187 OUT_N.n1163 GND 0.01fF $ **FLOATING
C1188 OUT_N.n1164 GND 0.05fF $ **FLOATING
C1189 OUT_N.n1165 GND 0.04fF $ **FLOATING
C1190 OUT_N.n1166 GND 0.01fF $ **FLOATING
C1191 OUT_N.n1167 GND 0.00fF $ **FLOATING
C1192 OUT_N.n1168 GND 0.01fF $ **FLOATING
C1193 OUT_N.n1169 GND 0.01fF $ **FLOATING
C1194 OUT_N.n1170 GND 0.02fF $ **FLOATING
C1195 OUT_N.n1171 GND 0.02fF $ **FLOATING
C1196 OUT_N.n1172 GND 0.01fF $ **FLOATING
C1197 OUT_N.t16 GND 0.25fF
C1198 OUT_N.n1173 GND 0.18fF $ **FLOATING
C1199 OUT_N.n1174 GND 0.03fF $ **FLOATING
C1200 OUT_N.n1175 GND 0.03fF $ **FLOATING
C1201 OUT_N.n1176 GND 0.01fF $ **FLOATING
C1202 OUT_N.n1177 GND 0.01fF $ **FLOATING
C1203 OUT_N.n1178 GND 0.01fF $ **FLOATING
C1204 OUT_N.n1179 GND 0.01fF $ **FLOATING
C1205 OUT_N.n1180 GND 0.01fF $ **FLOATING
C1206 OUT_N.n1181 GND 0.01fF $ **FLOATING
C1207 OUT_N.n1182 GND 0.01fF $ **FLOATING
C1208 OUT_N.n1183 GND 0.01fF $ **FLOATING
C1209 OUT_N.n1184 GND 0.01fF $ **FLOATING
C1210 OUT_N.n1185 GND 0.01fF $ **FLOATING
C1211 OUT_N.n1186 GND 0.07fF $ **FLOATING
C1212 OUT_N.n1187 GND 0.01fF $ **FLOATING
C1213 OUT_N.n1188 GND 0.03fF $ **FLOATING
C1214 OUT_N.n1189 GND 0.03fF $ **FLOATING
C1215 OUT_N.n1190 GND 0.01fF $ **FLOATING
C1216 OUT_N.n1191 GND 0.01fF $ **FLOATING
C1217 OUT_N.n1192 GND 0.00fF $ **FLOATING
C1218 OUT_N.n1193 GND 0.01fF $ **FLOATING
C1219 OUT_N.n1194 GND 0.01fF $ **FLOATING
C1220 OUT_N.n1195 GND 0.01fF $ **FLOATING
C1221 OUT_N.n1196 GND 0.01fF $ **FLOATING
C1222 OUT_N.n1197 GND 0.03fF $ **FLOATING
C1223 OUT_N.n1198 GND 0.01fF $ **FLOATING
C1224 OUT_N.n1199 GND 0.01fF $ **FLOATING
C1225 OUT_N.n1200 GND 0.01fF $ **FLOATING
C1226 OUT_N.n1201 GND 0.01fF $ **FLOATING
C1227 OUT_N.n1202 GND 0.01fF $ **FLOATING
C1228 OUT_N.n1203 GND 0.01fF $ **FLOATING
C1229 OUT_N.n1204 GND 0.26fF $ **FLOATING
C1230 OUT_N.n1205 GND 0.26fF $ **FLOATING
C1231 OUT_N.n1206 GND 0.01fF $ **FLOATING
C1232 OUT_N.n1207 GND 0.01fF $ **FLOATING
C1233 OUT_N.n1208 GND 0.03fF $ **FLOATING
C1234 OUT_N.n1209 GND 0.03fF $ **FLOATING
C1235 OUT_N.n1210 GND 0.01fF $ **FLOATING
C1236 OUT_N.n1211 GND 0.07fF $ **FLOATING
C1237 OUT_N.n1212 GND 0.01fF $ **FLOATING
C1238 OUT_N.n1213 GND 0.01fF $ **FLOATING
C1239 OUT_N.n1214 GND 0.01fF $ **FLOATING
C1240 OUT_N.n1215 GND 0.01fF $ **FLOATING
C1241 OUT_N.n1216 GND 0.01fF $ **FLOATING
C1242 OUT_N.n1217 GND 0.22fF $ **FLOATING
C1243 OUT_N.n1218 GND 0.23fF $ **FLOATING
C1244 OUT_N.n1219 GND 0.01fF $ **FLOATING
C1245 OUT_N.n1220 GND 0.01fF $ **FLOATING
C1246 OUT_N.n1221 GND 0.01fF $ **FLOATING
C1247 OUT_N.n1222 GND 0.01fF $ **FLOATING
C1248 OUT_N.n1223 GND 0.01fF $ **FLOATING
C1249 OUT_N.n1224 GND 0.01fF $ **FLOATING
C1250 OUT_N.n1225 GND 0.00fF $ **FLOATING
C1251 OUT_N.n1226 GND 0.01fF $ **FLOATING
C1252 OUT_N.n1227 GND 0.01fF $ **FLOATING
C1253 OUT_N.n1228 GND 0.01fF $ **FLOATING
C1254 OUT_N.n1229 GND 0.01fF $ **FLOATING
C1255 OUT_N.n1230 GND 0.01fF $ **FLOATING
C1256 OUT_N.n1231 GND 0.01fF $ **FLOATING
C1257 OUT_N.n1232 GND 0.01fF $ **FLOATING
C1258 OUT_N.n1233 GND 0.03fF $ **FLOATING
C1259 OUT_N.n1234 GND 0.01fF $ **FLOATING
C1260 OUT_N.n1235 GND 0.01fF $ **FLOATING
C1261 OUT_N.n1236 GND 0.01fF $ **FLOATING
C1262 OUT_N.n1237 GND 0.01fF $ **FLOATING
C1263 OUT_N.n1238 GND 0.01fF $ **FLOATING
C1264 OUT_N.n1239 GND 0.14fF $ **FLOATING
C1265 OUT_N.n1240 GND 0.01fF $ **FLOATING
C1266 OUT_N.n1241 GND 0.03fF $ **FLOATING
C1267 OUT_N.n1242 GND 0.03fF $ **FLOATING
C1268 OUT_N.n1243 GND 0.01fF $ **FLOATING
C1269 OUT_N.t20 GND 0.25fF
C1270 OUT_N.n1244 GND 0.18fF $ **FLOATING
C1271 OUT_N.n1245 GND 0.06fF $ **FLOATING
C1272 OUT_N.n1246 GND 0.01fF $ **FLOATING
C1273 OUT_N.n1247 GND 0.01fF $ **FLOATING
C1274 OUT_N.n1248 GND 0.01fF $ **FLOATING
C1275 OUT_N.n1249 GND 0.01fF $ **FLOATING
C1276 OUT_N.n1250 GND 0.01fF $ **FLOATING
C1277 OUT_N.n1251 GND 0.00fF $ **FLOATING
C1278 OUT_N.t24 GND 0.25fF
C1279 OUT_N.n1252 GND 0.18fF $ **FLOATING
C1280 OUT_N.n1253 GND 0.03fF $ **FLOATING
C1281 OUT_N.n1254 GND 0.03fF $ **FLOATING
C1282 OUT_N.n1255 GND 0.00fF $ **FLOATING
C1283 OUT_N.n1256 GND 0.01fF $ **FLOATING
C1284 OUT_N.n1257 GND 0.01fF $ **FLOATING
C1285 OUT_N.n1258 GND 0.02fF $ **FLOATING
C1286 OUT_N.n1259 GND 0.02fF $ **FLOATING
C1287 OUT_N.n1260 GND 0.01fF $ **FLOATING
C1288 OUT_N.n1261 GND 0.05fF $ **FLOATING
C1289 OUT_N.n1262 GND 0.04fF $ **FLOATING
C1290 OUT_N.n1263 GND 0.01fF $ **FLOATING
C1291 OUT_N.n1264 GND 0.01fF $ **FLOATING
C1292 OUT_N.n1265 GND 0.03fF $ **FLOATING
C1293 OUT_N.n1266 GND 0.03fF $ **FLOATING
C1294 OUT_N.n1267 GND 0.05fF $ **FLOATING
C1295 OUT_N.n1268 GND 0.06fF $ **FLOATING
C1296 OUT_N.n1269 GND 0.01fF $ **FLOATING
C1297 OUT_N.n1270 GND 0.01fF $ **FLOATING
C1298 OUT_N.n1271 GND 0.01fF $ **FLOATING
C1299 OUT_N.n1272 GND 0.02fF $ **FLOATING
C1300 OUT_N.n1273 GND 0.01fF $ **FLOATING
C1301 OUT_N.n1274 GND 0.01fF $ **FLOATING
C1302 OUT_N.n1275 GND 0.01fF $ **FLOATING
C1303 OUT_N.n1276 GND 0.26fF $ **FLOATING
C1304 OUT_N.n1277 GND 0.26fF $ **FLOATING
C1305 OUT_N.n1278 GND 0.01fF $ **FLOATING
C1306 OUT_N.n1279 GND 0.01fF $ **FLOATING
C1307 OUT_N.n1280 GND 0.03fF $ **FLOATING
C1308 OUT_N.n1281 GND 0.03fF $ **FLOATING
C1309 OUT_N.n1282 GND 0.01fF $ **FLOATING
C1310 OUT_N.n1283 GND 0.07fF $ **FLOATING
C1311 OUT_N.n1284 GND 0.01fF $ **FLOATING
C1312 OUT_N.n1285 GND 0.01fF $ **FLOATING
C1313 OUT_N.n1286 GND 0.01fF $ **FLOATING
C1314 OUT_N.n1287 GND 0.01fF $ **FLOATING
C1315 OUT_N.n1288 GND 0.01fF $ **FLOATING
C1316 OUT_N.t22 GND 0.25fF
C1317 OUT_N.n1289 GND 0.18fF $ **FLOATING
C1318 OUT_N.n1290 GND 0.03fF $ **FLOATING
C1319 OUT_N.n1291 GND 0.03fF $ **FLOATING
C1320 OUT_N.n1292 GND 0.01fF $ **FLOATING
C1321 OUT_N.n1293 GND 0.01fF $ **FLOATING
C1322 OUT_N.n1294 GND 0.02fF $ **FLOATING
C1323 OUT_N.n1295 GND 0.02fF $ **FLOATING
C1324 OUT_N.n1296 GND 0.01fF $ **FLOATING
C1325 OUT_N.n1297 GND 0.01fF $ **FLOATING
C1326 OUT_N.n1298 GND 0.00fF $ **FLOATING
C1327 OUT_N.n1299 GND 0.05fF $ **FLOATING
C1328 OUT_N.n1300 GND 0.04fF $ **FLOATING
C1329 OUT_N.n1301 GND 0.01fF $ **FLOATING
C1330 OUT_N.n1302 GND 0.01fF $ **FLOATING
C1331 OUT_N.n1303 GND 0.02fF $ **FLOATING
C1332 OUT_N.n1304 GND 0.02fF $ **FLOATING
C1333 OUT_N.n1305 GND 0.01fF $ **FLOATING
C1334 OUT_N.n1306 GND 0.03fF $ **FLOATING
C1335 OUT_N.n1307 GND 0.01fF $ **FLOATING
C1336 OUT_N.n1308 GND 0.01fF $ **FLOATING
C1337 OUT_N.n1309 GND 0.01fF $ **FLOATING
C1338 OUT_N.n1310 GND 0.01fF $ **FLOATING
C1339 OUT_N.n1311 GND 0.01fF $ **FLOATING
C1340 OUT_N.t26 GND 0.25fF
C1341 OUT_N.n1312 GND 0.18fF $ **FLOATING
C1342 OUT_N.n1313 GND 0.03fF $ **FLOATING
C1343 OUT_N.n1314 GND 0.03fF $ **FLOATING
C1344 OUT_N.n1315 GND 0.00fF $ **FLOATING
C1345 OUT_N.n1316 GND 0.01fF $ **FLOATING
C1346 OUT_N.n1317 GND 0.00fF $ **FLOATING
C1347 OUT_N.n1318 GND 0.01fF $ **FLOATING
C1348 OUT_N.n1319 GND 0.01fF $ **FLOATING
C1349 OUT_N.n1320 GND 0.01fF $ **FLOATING
C1350 OUT_N.n1321 GND 0.01fF $ **FLOATING
C1351 OUT_P.t27 GND 0.25fF
C1352 OUT_P.n0 GND 0.18fF $ **FLOATING
C1353 OUT_P.n1 GND 0.03fF $ **FLOATING
C1354 OUT_P.n2 GND 0.04fF $ **FLOATING
C1355 OUT_P.n3 GND 0.10fF $ **FLOATING
C1356 OUT_P.n4 GND 0.01fF $ **FLOATING
C1357 OUT_P.n5 GND 0.04fF $ **FLOATING
C1358 OUT_P.n6 GND 0.07fF $ **FLOATING
C1359 OUT_P.n7 GND 0.08fF $ **FLOATING
C1360 OUT_P.n8 GND 0.07fF $ **FLOATING
C1361 OUT_P.n9 GND 0.08fF $ **FLOATING
C1362 OUT_P.n10 GND 0.07fF $ **FLOATING
C1363 OUT_P.n11 GND 0.48fF $ **FLOATING
C1364 OUT_P.n12 GND 0.19fF $ **FLOATING
C1365 OUT_P.n13 GND 0.02fF $ **FLOATING
C1366 OUT_P.t3 GND 0.23fF
C1367 OUT_P.n14 GND 0.01fF $ **FLOATING
C1368 OUT_P.t1 GND 0.23fF
C1369 OUT_P.n15 GND 0.66fF $ **FLOATING
C1370 OUT_P.n16 GND 0.07fF $ **FLOATING
C1371 OUT_P.n17 GND 0.52fF $ **FLOATING
C1372 OUT_P.n18 GND 0.02fF $ **FLOATING
C1373 OUT_P.n19 GND 0.00fF $ **FLOATING
C1374 OUT_P.n20 GND 0.01fF $ **FLOATING
C1375 OUT_P.n21 GND 0.01fF $ **FLOATING
C1376 OUT_P.n22 GND 0.01fF $ **FLOATING
C1377 OUT_P.n23 GND 0.04fF $ **FLOATING
C1378 OUT_P.n24 GND 0.07fF $ **FLOATING
C1379 OUT_P.n25 GND 0.04fF $ **FLOATING
C1380 OUT_P.n26 GND 0.04fF $ **FLOATING
C1381 OUT_P.n27 GND 0.05fF $ **FLOATING
C1382 OUT_P.n28 GND 0.01fF $ **FLOATING
C1383 OUT_P.n29 GND 0.00fF $ **FLOATING
C1384 OUT_P.n30 GND 0.01fF $ **FLOATING
C1385 OUT_P.n31 GND 0.01fF $ **FLOATING
C1386 OUT_P.n32 GND 0.01fF $ **FLOATING
C1387 OUT_P.n33 GND 0.01fF $ **FLOATING
C1388 OUT_P.n34 GND 0.01fF $ **FLOATING
C1389 OUT_P.n35 GND 0.01fF $ **FLOATING
C1390 OUT_P.n36 GND 0.01fF $ **FLOATING
C1391 OUT_P.n37 GND 0.01fF $ **FLOATING
C1392 OUT_P.n38 GND 0.03fF $ **FLOATING
C1393 OUT_P.n39 GND 0.00fF $ **FLOATING
C1394 OUT_P.n40 GND 0.00fF $ **FLOATING
C1395 OUT_P.n41 GND 0.00fF $ **FLOATING
C1396 OUT_P.n42 GND 0.00fF $ **FLOATING
C1397 OUT_P.n43 GND 0.00fF $ **FLOATING
C1398 OUT_P.n44 GND 0.00fF $ **FLOATING
C1399 OUT_P.n45 GND 0.00fF $ **FLOATING
C1400 OUT_P.n46 GND 0.02fF $ **FLOATING
C1401 OUT_P.n47 GND 0.02fF $ **FLOATING
C1402 OUT_P.n48 GND 0.00fF $ **FLOATING
C1403 OUT_P.n49 GND 0.00fF $ **FLOATING
C1404 OUT_P.n50 GND 0.01fF $ **FLOATING
C1405 OUT_P.n51 GND 0.02fF $ **FLOATING
C1406 OUT_P.n52 GND 0.01fF $ **FLOATING
C1407 OUT_P.n53 GND 0.01fF $ **FLOATING
C1408 OUT_P.n54 GND 0.02fF $ **FLOATING
C1409 OUT_P.n55 GND 0.01fF $ **FLOATING
C1410 OUT_P.n56 GND 0.01fF $ **FLOATING
C1411 OUT_P.n57 GND 0.00fF $ **FLOATING
C1412 OUT_P.n58 GND 0.01fF $ **FLOATING
C1413 OUT_P.n59 GND 0.02fF $ **FLOATING
C1414 OUT_P.n60 GND 0.01fF $ **FLOATING
C1415 OUT_P.n61 GND 0.01fF $ **FLOATING
C1416 OUT_P.n62 GND 0.02fF $ **FLOATING
C1417 OUT_P.n63 GND 0.01fF $ **FLOATING
C1418 OUT_P.n64 GND 0.01fF $ **FLOATING
C1419 OUT_P.n65 GND 0.01fF $ **FLOATING
C1420 OUT_P.n66 GND 0.00fF $ **FLOATING
C1421 OUT_P.n67 GND 0.00fF $ **FLOATING
C1422 OUT_P.n68 GND 0.01fF $ **FLOATING
C1423 OUT_P.n69 GND 0.00fF $ **FLOATING
C1424 OUT_P.n70 GND 0.01fF $ **FLOATING
C1425 OUT_P.n71 GND 0.01fF $ **FLOATING
C1426 OUT_P.n72 GND 0.01fF $ **FLOATING
C1427 OUT_P.n73 GND 0.02fF $ **FLOATING
C1428 OUT_P.n74 GND 0.01fF $ **FLOATING
C1429 OUT_P.n75 GND 0.01fF $ **FLOATING
C1430 OUT_P.n76 GND 0.01fF $ **FLOATING
C1431 OUT_P.n77 GND 0.01fF $ **FLOATING
C1432 OUT_P.n78 GND 0.01fF $ **FLOATING
C1433 OUT_P.n79 GND 0.00fF $ **FLOATING
C1434 OUT_P.n80 GND 0.01fF $ **FLOATING
C1435 OUT_P.n81 GND 0.01fF $ **FLOATING
C1436 OUT_P.n82 GND 0.01fF $ **FLOATING
C1437 OUT_P.n83 GND 0.01fF $ **FLOATING
C1438 OUT_P.n84 GND 0.01fF $ **FLOATING
C1439 OUT_P.n85 GND 0.01fF $ **FLOATING
C1440 OUT_P.n86 GND 0.00fF $ **FLOATING
C1441 OUT_P.n87 GND 0.01fF $ **FLOATING
C1442 OUT_P.n88 GND 0.00fF $ **FLOATING
C1443 OUT_P.n89 GND 0.01fF $ **FLOATING
C1444 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0/DRAIN GND 0.02fF $ **FLOATING
C1445 OUT_P.n90 GND 0.05fF $ **FLOATING
C1446 OUT_P.n91 GND 0.04fF $ **FLOATING
C1447 OUT_P.n92 GND 0.04fF $ **FLOATING
C1448 OUT_P.n93 GND 0.08fF $ **FLOATING
C1449 OUT_P.n94 GND 0.08fF $ **FLOATING
C1450 OUT_P.n95 GND 0.04fF $ **FLOATING
C1451 OUT_P.n96 GND 0.04fF $ **FLOATING
C1452 OUT_P.n97 GND 0.08fF $ **FLOATING
C1453 OUT_P.n98 GND 0.07fF $ **FLOATING
C1454 OUT_P.n99 GND 0.05fF $ **FLOATING
C1455 OUT_P.n100 GND 0.10fF $ **FLOATING
C1456 OUT_P.n101 GND 0.10fF $ **FLOATING
C1457 OUT_P.n102 GND 0.05fF $ **FLOATING
C1458 OUT_P.n103 GND 0.10fF $ **FLOATING
C1459 OUT_P.n104 GND 0.09fF $ **FLOATING
C1460 OUT_P.n105 GND 0.05fF $ **FLOATING
C1461 OUT_P.n106 GND 0.05fF $ **FLOATING
C1462 OUT_P.n107 GND 0.02fF $ **FLOATING
C1463 OUT_P.n108 GND 0.02fF $ **FLOATING
C1464 OUT_P.n109 GND 0.04fF $ **FLOATING
C1465 OUT_P.n110 GND 0.03fF $ **FLOATING
C1466 OUT_P.n111 GND 0.21fF $ **FLOATING
C1467 OUT_P.n112 GND 0.16fF $ **FLOATING
C1468 OUT_P.n114 GND 0.12fF $ **FLOATING
C1469 OUT_P.n115 GND 0.99fF $ **FLOATING
C1470 OUT_P.n116 GND 1.02fF $ **FLOATING
C1471 OUT_P.n117 GND 0.19fF $ **FLOATING
C1472 OUT_P.n118 GND 0.01fF $ **FLOATING
C1473 OUT_P.t8 GND 0.23fF
C1474 OUT_P.n119 GND 0.01fF $ **FLOATING
C1475 OUT_P.t10 GND 0.23fF
C1476 OUT_P.n120 GND 0.66fF $ **FLOATING
C1477 OUT_P.n121 GND 0.07fF $ **FLOATING
C1478 OUT_P.n122 GND 0.52fF $ **FLOATING
C1479 OUT_P.n123 GND 0.02fF $ **FLOATING
C1480 OUT_P.n124 GND 0.00fF $ **FLOATING
C1481 OUT_P.n125 GND 0.01fF $ **FLOATING
C1482 OUT_P.n126 GND 0.01fF $ **FLOATING
C1483 OUT_P.n127 GND 0.01fF $ **FLOATING
C1484 OUT_P.n128 GND 0.04fF $ **FLOATING
C1485 OUT_P.n129 GND 0.07fF $ **FLOATING
C1486 OUT_P.n130 GND 0.04fF $ **FLOATING
C1487 OUT_P.n131 GND 0.04fF $ **FLOATING
C1488 OUT_P.n132 GND 0.05fF $ **FLOATING
C1489 OUT_P.n133 GND 0.01fF $ **FLOATING
C1490 OUT_P.n134 GND 0.00fF $ **FLOATING
C1491 OUT_P.n135 GND 0.01fF $ **FLOATING
C1492 OUT_P.n136 GND 0.01fF $ **FLOATING
C1493 OUT_P.n137 GND 0.01fF $ **FLOATING
C1494 OUT_P.n138 GND 0.01fF $ **FLOATING
C1495 OUT_P.n139 GND 0.01fF $ **FLOATING
C1496 OUT_P.n140 GND 0.01fF $ **FLOATING
C1497 OUT_P.n141 GND 0.01fF $ **FLOATING
C1498 OUT_P.n142 GND 0.01fF $ **FLOATING
C1499 OUT_P.n143 GND 0.03fF $ **FLOATING
C1500 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2/DRAIN GND 0.02fF $ **FLOATING
C1501 OUT_P.n144 GND 0.05fF $ **FLOATING
C1502 OUT_P.n145 GND 0.04fF $ **FLOATING
C1503 OUT_P.n146 GND 0.04fF $ **FLOATING
C1504 OUT_P.n147 GND 0.08fF $ **FLOATING
C1505 OUT_P.n148 GND 0.08fF $ **FLOATING
C1506 OUT_P.n149 GND 0.04fF $ **FLOATING
C1507 OUT_P.n150 GND 0.04fF $ **FLOATING
C1508 OUT_P.n151 GND 0.08fF $ **FLOATING
C1509 OUT_P.n152 GND 0.07fF $ **FLOATING
C1510 OUT_P.n153 GND 0.05fF $ **FLOATING
C1511 OUT_P.n154 GND 0.10fF $ **FLOATING
C1512 OUT_P.n155 GND 0.10fF $ **FLOATING
C1513 OUT_P.n156 GND 0.05fF $ **FLOATING
C1514 OUT_P.n157 GND 0.10fF $ **FLOATING
C1515 OUT_P.n158 GND 0.09fF $ **FLOATING
C1516 OUT_P.n159 GND 0.05fF $ **FLOATING
C1517 OUT_P.n160 GND 0.05fF $ **FLOATING
C1518 OUT_P.n161 GND 0.00fF $ **FLOATING
C1519 OUT_P.n162 GND 0.00fF $ **FLOATING
C1520 OUT_P.n163 GND 0.00fF $ **FLOATING
C1521 OUT_P.n164 GND 0.00fF $ **FLOATING
C1522 OUT_P.n165 GND 0.00fF $ **FLOATING
C1523 OUT_P.n166 GND 0.00fF $ **FLOATING
C1524 OUT_P.n167 GND 0.00fF $ **FLOATING
C1525 OUT_P.n168 GND 0.00fF $ **FLOATING
C1526 OUT_P.n169 GND 0.02fF $ **FLOATING
C1527 OUT_P.n170 GND 0.02fF $ **FLOATING
C1528 OUT_P.n171 GND 0.00fF $ **FLOATING
C1529 OUT_P.n172 GND 0.01fF $ **FLOATING
C1530 OUT_P.n173 GND 0.02fF $ **FLOATING
C1531 OUT_P.n174 GND 0.01fF $ **FLOATING
C1532 OUT_P.n175 GND 0.01fF $ **FLOATING
C1533 OUT_P.n176 GND 0.02fF $ **FLOATING
C1534 OUT_P.n177 GND 0.01fF $ **FLOATING
C1535 OUT_P.n178 GND 0.01fF $ **FLOATING
C1536 OUT_P.n179 GND 0.00fF $ **FLOATING
C1537 OUT_P.n180 GND 0.01fF $ **FLOATING
C1538 OUT_P.n181 GND 0.02fF $ **FLOATING
C1539 OUT_P.n182 GND 0.01fF $ **FLOATING
C1540 OUT_P.n183 GND 0.01fF $ **FLOATING
C1541 OUT_P.n184 GND 0.02fF $ **FLOATING
C1542 OUT_P.n185 GND 0.01fF $ **FLOATING
C1543 OUT_P.n186 GND 0.01fF $ **FLOATING
C1544 OUT_P.n187 GND 0.01fF $ **FLOATING
C1545 OUT_P.n188 GND 0.00fF $ **FLOATING
C1546 OUT_P.n189 GND 0.01fF $ **FLOATING
C1547 OUT_P.n190 GND 0.00fF $ **FLOATING
C1548 OUT_P.n191 GND 0.01fF $ **FLOATING
C1549 OUT_P.n192 GND 0.01fF $ **FLOATING
C1550 OUT_P.n193 GND 0.01fF $ **FLOATING
C1551 OUT_P.n194 GND 0.02fF $ **FLOATING
C1552 OUT_P.n195 GND 0.01fF $ **FLOATING
C1553 OUT_P.n196 GND 0.01fF $ **FLOATING
C1554 OUT_P.n197 GND 0.01fF $ **FLOATING
C1555 OUT_P.n198 GND 0.01fF $ **FLOATING
C1556 OUT_P.n199 GND 0.00fF $ **FLOATING
C1557 OUT_P.n200 GND 0.01fF $ **FLOATING
C1558 OUT_P.n201 GND 0.00fF $ **FLOATING
C1559 OUT_P.n202 GND 0.01fF $ **FLOATING
C1560 OUT_P.n203 GND 0.01fF $ **FLOATING
C1561 OUT_P.n204 GND 0.01fF $ **FLOATING
C1562 OUT_P.n205 GND 0.01fF $ **FLOATING
C1563 OUT_P.n206 GND 0.01fF $ **FLOATING
C1564 OUT_P.n207 GND 0.01fF $ **FLOATING
C1565 OUT_P.n208 GND 0.00fF $ **FLOATING
C1566 OUT_P.n209 GND 0.01fF $ **FLOATING
C1567 OUT_P.n210 GND 0.00fF $ **FLOATING
C1568 OUT_P.n211 GND 0.01fF $ **FLOATING
C1569 OUT_P.n212 GND 0.02fF $ **FLOATING
C1570 OUT_P.n213 GND 0.02fF $ **FLOATING
C1571 OUT_P.n214 GND 0.04fF $ **FLOATING
C1572 OUT_P.n215 GND 0.03fF $ **FLOATING
C1573 OUT_P.n217 GND 0.16fF $ **FLOATING
C1574 OUT_P.n219 GND 0.12fF $ **FLOATING
C1575 OUT_P.n220 GND 0.99fF $ **FLOATING
C1576 OUT_P.n221 GND 1.02fF $ **FLOATING
C1577 OUT_P.n222 GND 0.19fF $ **FLOATING
C1578 OUT_P.n223 GND 0.01fF $ **FLOATING
C1579 OUT_P.t13 GND 0.23fF
C1580 OUT_P.n224 GND 0.01fF $ **FLOATING
C1581 OUT_P.t6 GND 0.23fF
C1582 OUT_P.n225 GND 0.66fF $ **FLOATING
C1583 OUT_P.n226 GND 0.07fF $ **FLOATING
C1584 OUT_P.n227 GND 0.52fF $ **FLOATING
C1585 OUT_P.n228 GND 0.02fF $ **FLOATING
C1586 OUT_P.n229 GND 0.00fF $ **FLOATING
C1587 OUT_P.n230 GND 0.01fF $ **FLOATING
C1588 OUT_P.n231 GND 0.01fF $ **FLOATING
C1589 OUT_P.n232 GND 0.01fF $ **FLOATING
C1590 OUT_P.n233 GND 0.04fF $ **FLOATING
C1591 OUT_P.n234 GND 0.07fF $ **FLOATING
C1592 OUT_P.n235 GND 0.04fF $ **FLOATING
C1593 OUT_P.n236 GND 0.04fF $ **FLOATING
C1594 OUT_P.n237 GND 0.05fF $ **FLOATING
C1595 OUT_P.n238 GND 0.01fF $ **FLOATING
C1596 OUT_P.n239 GND 0.00fF $ **FLOATING
C1597 OUT_P.n240 GND 0.01fF $ **FLOATING
C1598 OUT_P.n241 GND 0.01fF $ **FLOATING
C1599 OUT_P.n242 GND 0.01fF $ **FLOATING
C1600 OUT_P.n243 GND 0.01fF $ **FLOATING
C1601 OUT_P.n244 GND 0.01fF $ **FLOATING
C1602 OUT_P.n245 GND 0.01fF $ **FLOATING
C1603 OUT_P.n246 GND 0.01fF $ **FLOATING
C1604 OUT_P.n247 GND 0.01fF $ **FLOATING
C1605 OUT_P.n248 GND 0.03fF $ **FLOATING
C1606 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4/DRAIN GND 0.02fF $ **FLOATING
C1607 OUT_P.n249 GND 0.05fF $ **FLOATING
C1608 OUT_P.n250 GND 0.04fF $ **FLOATING
C1609 OUT_P.n251 GND 0.04fF $ **FLOATING
C1610 OUT_P.n252 GND 0.08fF $ **FLOATING
C1611 OUT_P.n253 GND 0.08fF $ **FLOATING
C1612 OUT_P.n254 GND 0.04fF $ **FLOATING
C1613 OUT_P.n255 GND 0.04fF $ **FLOATING
C1614 OUT_P.n256 GND 0.08fF $ **FLOATING
C1615 OUT_P.n257 GND 0.07fF $ **FLOATING
C1616 OUT_P.n258 GND 0.05fF $ **FLOATING
C1617 OUT_P.n259 GND 0.10fF $ **FLOATING
C1618 OUT_P.n260 GND 0.10fF $ **FLOATING
C1619 OUT_P.n261 GND 0.05fF $ **FLOATING
C1620 OUT_P.n262 GND 0.10fF $ **FLOATING
C1621 OUT_P.n263 GND 0.09fF $ **FLOATING
C1622 OUT_P.n264 GND 0.05fF $ **FLOATING
C1623 OUT_P.n265 GND 0.05fF $ **FLOATING
C1624 OUT_P.n266 GND 0.00fF $ **FLOATING
C1625 OUT_P.n267 GND 0.00fF $ **FLOATING
C1626 OUT_P.n268 GND 0.00fF $ **FLOATING
C1627 OUT_P.n269 GND 0.00fF $ **FLOATING
C1628 OUT_P.n270 GND 0.00fF $ **FLOATING
C1629 OUT_P.n271 GND 0.00fF $ **FLOATING
C1630 OUT_P.n272 GND 0.00fF $ **FLOATING
C1631 OUT_P.n273 GND 0.00fF $ **FLOATING
C1632 OUT_P.n274 GND 0.02fF $ **FLOATING
C1633 OUT_P.n275 GND 0.02fF $ **FLOATING
C1634 OUT_P.n276 GND 0.00fF $ **FLOATING
C1635 OUT_P.n277 GND 0.01fF $ **FLOATING
C1636 OUT_P.n278 GND 0.02fF $ **FLOATING
C1637 OUT_P.n279 GND 0.01fF $ **FLOATING
C1638 OUT_P.n280 GND 0.01fF $ **FLOATING
C1639 OUT_P.n281 GND 0.02fF $ **FLOATING
C1640 OUT_P.n282 GND 0.01fF $ **FLOATING
C1641 OUT_P.n283 GND 0.01fF $ **FLOATING
C1642 OUT_P.n284 GND 0.00fF $ **FLOATING
C1643 OUT_P.n285 GND 0.01fF $ **FLOATING
C1644 OUT_P.n286 GND 0.02fF $ **FLOATING
C1645 OUT_P.n287 GND 0.01fF $ **FLOATING
C1646 OUT_P.n288 GND 0.01fF $ **FLOATING
C1647 OUT_P.n289 GND 0.02fF $ **FLOATING
C1648 OUT_P.n290 GND 0.01fF $ **FLOATING
C1649 OUT_P.n291 GND 0.01fF $ **FLOATING
C1650 OUT_P.n292 GND 0.01fF $ **FLOATING
C1651 OUT_P.n293 GND 0.00fF $ **FLOATING
C1652 OUT_P.n294 GND 0.01fF $ **FLOATING
C1653 OUT_P.n295 GND 0.00fF $ **FLOATING
C1654 OUT_P.n296 GND 0.01fF $ **FLOATING
C1655 OUT_P.n297 GND 0.01fF $ **FLOATING
C1656 OUT_P.n298 GND 0.01fF $ **FLOATING
C1657 OUT_P.n299 GND 0.02fF $ **FLOATING
C1658 OUT_P.n300 GND 0.01fF $ **FLOATING
C1659 OUT_P.n301 GND 0.01fF $ **FLOATING
C1660 OUT_P.n302 GND 0.01fF $ **FLOATING
C1661 OUT_P.n303 GND 0.01fF $ **FLOATING
C1662 OUT_P.n304 GND 0.00fF $ **FLOATING
C1663 OUT_P.n305 GND 0.01fF $ **FLOATING
C1664 OUT_P.n306 GND 0.00fF $ **FLOATING
C1665 OUT_P.n307 GND 0.01fF $ **FLOATING
C1666 OUT_P.n308 GND 0.01fF $ **FLOATING
C1667 OUT_P.n309 GND 0.01fF $ **FLOATING
C1668 OUT_P.n310 GND 0.01fF $ **FLOATING
C1669 OUT_P.n311 GND 0.01fF $ **FLOATING
C1670 OUT_P.n312 GND 0.01fF $ **FLOATING
C1671 OUT_P.n313 GND 0.00fF $ **FLOATING
C1672 OUT_P.n314 GND 0.01fF $ **FLOATING
C1673 OUT_P.n315 GND 0.00fF $ **FLOATING
C1674 OUT_P.n316 GND 0.01fF $ **FLOATING
C1675 OUT_P.n317 GND 0.02fF $ **FLOATING
C1676 OUT_P.n318 GND 0.02fF $ **FLOATING
C1677 OUT_P.n319 GND 0.04fF $ **FLOATING
C1678 OUT_P.n320 GND 0.03fF $ **FLOATING
C1679 OUT_P.n322 GND 0.16fF $ **FLOATING
C1680 OUT_P.n324 GND 0.12fF $ **FLOATING
C1681 OUT_P.n325 GND 0.99fF $ **FLOATING
C1682 OUT_P.n326 GND 1.02fF $ **FLOATING
C1683 OUT_P.n327 GND 0.19fF $ **FLOATING
C1684 OUT_P.n328 GND 0.01fF $ **FLOATING
C1685 OUT_P.t11 GND 0.23fF
C1686 OUT_P.n329 GND 0.01fF $ **FLOATING
C1687 OUT_P.t7 GND 0.23fF
C1688 OUT_P.n330 GND 0.66fF $ **FLOATING
C1689 OUT_P.n331 GND 0.07fF $ **FLOATING
C1690 OUT_P.n332 GND 0.52fF $ **FLOATING
C1691 OUT_P.n333 GND 0.02fF $ **FLOATING
C1692 OUT_P.n334 GND 0.00fF $ **FLOATING
C1693 OUT_P.n335 GND 0.01fF $ **FLOATING
C1694 OUT_P.n336 GND 0.01fF $ **FLOATING
C1695 OUT_P.n337 GND 0.01fF $ **FLOATING
C1696 OUT_P.n338 GND 0.04fF $ **FLOATING
C1697 OUT_P.n339 GND 0.07fF $ **FLOATING
C1698 OUT_P.n340 GND 0.04fF $ **FLOATING
C1699 OUT_P.n341 GND 0.04fF $ **FLOATING
C1700 OUT_P.n342 GND 0.05fF $ **FLOATING
C1701 OUT_P.n343 GND 0.01fF $ **FLOATING
C1702 OUT_P.n344 GND 0.00fF $ **FLOATING
C1703 OUT_P.n345 GND 0.01fF $ **FLOATING
C1704 OUT_P.n346 GND 0.01fF $ **FLOATING
C1705 OUT_P.n347 GND 0.01fF $ **FLOATING
C1706 OUT_P.n348 GND 0.01fF $ **FLOATING
C1707 OUT_P.n349 GND 0.01fF $ **FLOATING
C1708 OUT_P.n350 GND 0.01fF $ **FLOATING
C1709 OUT_P.n351 GND 0.01fF $ **FLOATING
C1710 OUT_P.n352 GND 0.01fF $ **FLOATING
C1711 OUT_P.n353 GND 0.03fF $ **FLOATING
C1712 OUT_P.n354 GND 0.05fF $ **FLOATING
C1713 OUT_P.n355 GND 0.04fF $ **FLOATING
C1714 OUT_P.n356 GND 0.04fF $ **FLOATING
C1715 OUT_P.n357 GND 0.08fF $ **FLOATING
C1716 OUT_P.n358 GND 0.08fF $ **FLOATING
C1717 OUT_P.n359 GND 0.04fF $ **FLOATING
C1718 OUT_P.n360 GND 0.04fF $ **FLOATING
C1719 OUT_P.n361 GND 0.08fF $ **FLOATING
C1720 OUT_P.n362 GND 0.07fF $ **FLOATING
C1721 OUT_P.n363 GND 0.05fF $ **FLOATING
C1722 OUT_P.n364 GND 0.10fF $ **FLOATING
C1723 OUT_P.n365 GND 0.10fF $ **FLOATING
C1724 OUT_P.n366 GND 0.05fF $ **FLOATING
C1725 OUT_P.n367 GND 0.10fF $ **FLOATING
C1726 OUT_P.n368 GND 0.09fF $ **FLOATING
C1727 OUT_P.n369 GND 0.05fF $ **FLOATING
C1728 OUT_P.n370 GND 0.05fF $ **FLOATING
C1729 OUT_P.n371 GND 0.00fF $ **FLOATING
C1730 OUT_P.n372 GND 0.00fF $ **FLOATING
C1731 OUT_P.n373 GND 0.00fF $ **FLOATING
C1732 OUT_P.n374 GND 0.00fF $ **FLOATING
C1733 OUT_P.n375 GND 0.00fF $ **FLOATING
C1734 OUT_P.n376 GND 0.00fF $ **FLOATING
C1735 OUT_P.n377 GND 0.00fF $ **FLOATING
C1736 OUT_P.n378 GND 0.00fF $ **FLOATING
C1737 OUT_P.n379 GND 0.02fF $ **FLOATING
C1738 OUT_P.n380 GND 0.02fF $ **FLOATING
C1739 OUT_P.n381 GND 0.00fF $ **FLOATING
C1740 OUT_P.n382 GND 0.01fF $ **FLOATING
C1741 OUT_P.n383 GND 0.02fF $ **FLOATING
C1742 OUT_P.n384 GND 0.01fF $ **FLOATING
C1743 OUT_P.n385 GND 0.01fF $ **FLOATING
C1744 OUT_P.n386 GND 0.02fF $ **FLOATING
C1745 OUT_P.n387 GND 0.01fF $ **FLOATING
C1746 OUT_P.n388 GND 0.01fF $ **FLOATING
C1747 OUT_P.n389 GND 0.00fF $ **FLOATING
C1748 OUT_P.n390 GND 0.01fF $ **FLOATING
C1749 OUT_P.n391 GND 0.02fF $ **FLOATING
C1750 OUT_P.n392 GND 0.01fF $ **FLOATING
C1751 OUT_P.n393 GND 0.01fF $ **FLOATING
C1752 OUT_P.n394 GND 0.02fF $ **FLOATING
C1753 OUT_P.n395 GND 0.01fF $ **FLOATING
C1754 OUT_P.n396 GND 0.01fF $ **FLOATING
C1755 OUT_P.n397 GND 0.01fF $ **FLOATING
C1756 OUT_P.n398 GND 0.00fF $ **FLOATING
C1757 OUT_P.n399 GND 0.01fF $ **FLOATING
C1758 OUT_P.n400 GND 0.00fF $ **FLOATING
C1759 OUT_P.n401 GND 0.01fF $ **FLOATING
C1760 OUT_P.n402 GND 0.01fF $ **FLOATING
C1761 OUT_P.n403 GND 0.01fF $ **FLOATING
C1762 OUT_P.n404 GND 0.02fF $ **FLOATING
C1763 OUT_P.n405 GND 0.01fF $ **FLOATING
C1764 OUT_P.n406 GND 0.01fF $ **FLOATING
C1765 OUT_P.n407 GND 0.01fF $ **FLOATING
C1766 OUT_P.n408 GND 0.01fF $ **FLOATING
C1767 OUT_P.n409 GND 0.00fF $ **FLOATING
C1768 OUT_P.n410 GND 0.01fF $ **FLOATING
C1769 OUT_P.n411 GND 0.00fF $ **FLOATING
C1770 OUT_P.n412 GND 0.01fF $ **FLOATING
C1771 OUT_P.n413 GND 0.01fF $ **FLOATING
C1772 OUT_P.n414 GND 0.01fF $ **FLOATING
C1773 OUT_P.n415 GND 0.01fF $ **FLOATING
C1774 OUT_P.n416 GND 0.01fF $ **FLOATING
C1775 OUT_P.n417 GND 0.01fF $ **FLOATING
C1776 OUT_P.n418 GND 0.00fF $ **FLOATING
C1777 OUT_P.n419 GND 0.01fF $ **FLOATING
C1778 OUT_P.n420 GND 0.00fF $ **FLOATING
C1779 OUT_P.n421 GND 0.01fF $ **FLOATING
C1780 OUT_P.n422 GND 0.02fF $ **FLOATING
C1781 OUT_P.n423 GND 0.02fF $ **FLOATING
C1782 OUT_P.n424 GND 0.04fF $ **FLOATING
C1783 OUT_P.n425 GND 0.03fF $ **FLOATING
C1784 OUT_P.n427 GND 0.16fF $ **FLOATING
C1785 OUT_P.n429 GND 0.12fF $ **FLOATING
C1786 OUT_P.n430 GND 0.96fF $ **FLOATING
C1787 OUT_P.n431 GND 1.00fF $ **FLOATING
C1788 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5/GATE GND 0.00fF $ **FLOATING
C1789 OUT_P.n433 GND 0.01fF $ **FLOATING
C1790 OUT_P.n434 GND 0.01fF $ **FLOATING
C1791 OUT_P.n435 GND 0.01fF $ **FLOATING
C1792 OUT_P.n436 GND 0.01fF $ **FLOATING
C1793 OUT_P.n437 GND 0.01fF $ **FLOATING
C1794 OUT_P.n438 GND 0.00fF $ **FLOATING
C1795 OUT_P.n439 GND 0.18fF $ **FLOATING
C1796 OUT_P.n440 GND 0.03fF $ **FLOATING
C1797 OUT_P.n441 GND 0.03fF $ **FLOATING
C1798 OUT_P.n442 GND 0.00fF $ **FLOATING
C1799 OUT_P.n443 GND 0.01fF $ **FLOATING
C1800 OUT_P.n444 GND 0.01fF $ **FLOATING
C1801 OUT_P.n445 GND 0.02fF $ **FLOATING
C1802 OUT_P.n446 GND 0.02fF $ **FLOATING
C1803 OUT_P.n447 GND 0.01fF $ **FLOATING
C1804 OUT_P.n448 GND 0.05fF $ **FLOATING
C1805 OUT_P.n449 GND 0.04fF $ **FLOATING
C1806 OUT_P.n450 GND 0.01fF $ **FLOATING
C1807 OUT_P.n451 GND 0.00fF $ **FLOATING
C1808 OUT_P.n452 GND 0.01fF $ **FLOATING
C1809 OUT_P.n453 GND 0.01fF $ **FLOATING
C1810 OUT_P.n454 GND 0.02fF $ **FLOATING
C1811 OUT_P.n455 GND 0.03fF $ **FLOATING
C1812 OUT_P.n456 GND 0.18fF $ **FLOATING
C1813 OUT_P.n457 GND 0.06fF $ **FLOATING
C1814 OUT_P.n458 GND 0.06fF $ **FLOATING
C1815 OUT_P.n459 GND 0.06fF $ **FLOATING
C1816 OUT_P.n460 GND 0.01fF $ **FLOATING
C1817 OUT_P.n461 GND 0.01fF $ **FLOATING
C1818 OUT_P.n462 GND 0.00fF $ **FLOATING
C1819 OUT_P.n463 GND 0.01fF $ **FLOATING
C1820 OUT_P.n464 GND 0.01fF $ **FLOATING
C1821 OUT_P.n465 GND 0.01fF $ **FLOATING
C1822 OUT_P.n466 GND 0.01fF $ **FLOATING
C1823 OUT_P.n467 GND 0.01fF $ **FLOATING
C1824 OUT_P.n468 GND 0.01fF $ **FLOATING
C1825 OUT_P.n469 GND 0.01fF $ **FLOATING
C1826 OUT_P.n470 GND 0.01fF $ **FLOATING
C1827 OUT_P.n471 GND 0.04fF $ **FLOATING
C1828 OUT_P.n472 GND 0.01fF $ **FLOATING
C1829 OUT_P.n473 GND 0.01fF $ **FLOATING
C1830 OUT_P.n474 GND 0.01fF $ **FLOATING
C1831 OUT_P.n475 GND 0.01fF $ **FLOATING
C1832 OUT_P.n476 GND 0.01fF $ **FLOATING
C1833 OUT_P.n477 GND 0.01fF $ **FLOATING
C1834 OUT_P.n478 GND 0.01fF $ **FLOATING
C1835 OUT_P.n479 GND 0.00fF $ **FLOATING
C1836 OUT_P.n480 GND 0.01fF $ **FLOATING
C1837 OUT_P.n481 GND 0.03fF $ **FLOATING
C1838 OUT_P.n482 GND 0.01fF $ **FLOATING
C1839 OUT_P.n483 GND 0.01fF $ **FLOATING
C1840 OUT_P.n484 GND 0.01fF $ **FLOATING
C1841 OUT_P.n485 GND 0.00fF $ **FLOATING
C1842 OUT_P.n486 GND 0.18fF $ **FLOATING
C1843 OUT_P.n487 GND 0.03fF $ **FLOATING
C1844 OUT_P.n488 GND 0.03fF $ **FLOATING
C1845 OUT_P.n489 GND 0.01fF $ **FLOATING
C1846 OUT_P.n490 GND 0.01fF $ **FLOATING
C1847 OUT_P.n491 GND 0.02fF $ **FLOATING
C1848 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9/GATE GND 0.00fF $ **FLOATING
C1849 OUT_P.n492 GND 0.01fF $ **FLOATING
C1850 OUT_P.n493 GND 0.02fF $ **FLOATING
C1851 OUT_P.n494 GND 0.01fF $ **FLOATING
C1852 OUT_P.n495 GND 0.01fF $ **FLOATING
C1853 OUT_P.n496 GND 0.00fF $ **FLOATING
C1854 OUT_P.n497 GND 0.18fF $ **FLOATING
C1855 OUT_P.n498 GND 0.03fF $ **FLOATING
C1856 OUT_P.n499 GND 0.03fF $ **FLOATING
C1857 OUT_P.n500 GND 0.01fF $ **FLOATING
C1858 OUT_P.n501 GND 0.01fF $ **FLOATING
C1859 OUT_P.n502 GND 0.01fF $ **FLOATING
C1860 OUT_P.n503 GND 0.02fF $ **FLOATING
C1861 OUT_P.n504 GND 0.02fF $ **FLOATING
C1862 OUT_P.n505 GND 0.01fF $ **FLOATING
C1863 OUT_P.n506 GND 0.05fF $ **FLOATING
C1864 OUT_P.n507 GND 0.04fF $ **FLOATING
C1865 OUT_P.n508 GND 0.01fF $ **FLOATING
C1866 OUT_P.n509 GND 0.00fF $ **FLOATING
C1867 OUT_P.n510 GND 0.01fF $ **FLOATING
C1868 OUT_P.n511 GND 0.03fF $ **FLOATING
C1869 OUT_P.n512 GND 0.02fF $ **FLOATING
C1870 OUT_P.n513 GND 0.01fF $ **FLOATING
C1871 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3/GATE GND 0.00fF $ **FLOATING
C1872 OUT_P.n514 GND 0.01fF $ **FLOATING
C1873 OUT_P.n515 GND 0.01fF $ **FLOATING
C1874 OUT_P.n516 GND 0.01fF $ **FLOATING
C1875 OUT_P.n517 GND 0.01fF $ **FLOATING
C1876 OUT_P.n518 GND 0.01fF $ **FLOATING
C1877 OUT_P.n519 GND 0.00fF $ **FLOATING
C1878 OUT_P.n520 GND 0.18fF $ **FLOATING
C1879 OUT_P.n521 GND 0.03fF $ **FLOATING
C1880 OUT_P.n522 GND 0.03fF $ **FLOATING
C1881 OUT_P.n523 GND 0.00fF $ **FLOATING
C1882 OUT_P.n524 GND 0.01fF $ **FLOATING
C1883 OUT_P.n525 GND 0.01fF $ **FLOATING
C1884 OUT_P.n526 GND 0.02fF $ **FLOATING
C1885 OUT_P.n527 GND 0.02fF $ **FLOATING
C1886 OUT_P.n528 GND 0.01fF $ **FLOATING
C1887 OUT_P.n529 GND 0.05fF $ **FLOATING
C1888 OUT_P.n530 GND 0.04fF $ **FLOATING
C1889 OUT_P.n531 GND 0.01fF $ **FLOATING
C1890 OUT_P.n532 GND 0.00fF $ **FLOATING
C1891 OUT_P.n533 GND 0.01fF $ **FLOATING
C1892 OUT_P.n534 GND 0.01fF $ **FLOATING
C1893 OUT_P.n535 GND 0.02fF $ **FLOATING
C1894 OUT_P.n536 GND 0.03fF $ **FLOATING
C1895 OUT_P.n537 GND 0.18fF $ **FLOATING
C1896 OUT_P.n538 GND 0.06fF $ **FLOATING
C1897 OUT_P.n539 GND 0.06fF $ **FLOATING
C1898 OUT_P.n540 GND 0.06fF $ **FLOATING
C1899 OUT_P.n541 GND 0.01fF $ **FLOATING
C1900 OUT_P.n542 GND 0.01fF $ **FLOATING
C1901 OUT_P.n543 GND 0.00fF $ **FLOATING
C1902 OUT_P.n544 GND 0.01fF $ **FLOATING
C1903 OUT_P.n545 GND 0.01fF $ **FLOATING
C1904 OUT_P.n546 GND 0.01fF $ **FLOATING
C1905 OUT_P.n547 GND 0.01fF $ **FLOATING
C1906 OUT_P.n548 GND 0.01fF $ **FLOATING
C1907 OUT_P.n549 GND 0.01fF $ **FLOATING
C1908 OUT_P.n550 GND 0.01fF $ **FLOATING
C1909 OUT_P.n551 GND 0.01fF $ **FLOATING
C1910 OUT_P.n552 GND 0.03fF $ **FLOATING
C1911 OUT_P.n553 GND 0.01fF $ **FLOATING
C1912 OUT_P.n554 GND 0.01fF $ **FLOATING
C1913 OUT_P.n555 GND 0.01fF $ **FLOATING
C1914 OUT_P.n556 GND 0.01fF $ **FLOATING
C1915 OUT_P.n557 GND 0.01fF $ **FLOATING
C1916 OUT_P.n558 GND 0.01fF $ **FLOATING
C1917 OUT_P.n559 GND 0.01fF $ **FLOATING
C1918 OUT_P.n560 GND 0.01fF $ **FLOATING
C1919 OUT_P.n561 GND 0.01fF $ **FLOATING
C1920 OUT_P.n562 GND 0.01fF $ **FLOATING
C1921 OUT_P.n563 GND 0.02fF $ **FLOATING
C1922 OUT_P.n564 GND 0.01fF $ **FLOATING
C1923 OUT_P.n565 GND 0.01fF $ **FLOATING
C1924 OUT_P.n566 GND 0.01fF $ **FLOATING
C1925 OUT_P.n567 GND 0.18fF $ **FLOATING
C1926 OUT_P.n568 GND 0.03fF $ **FLOATING
C1927 OUT_P.n569 GND 0.03fF $ **FLOATING
C1928 OUT_P.n570 GND 0.00fF $ **FLOATING
C1929 OUT_P.n571 GND 0.01fF $ **FLOATING
C1930 OUT_P.n572 GND 0.01fF $ **FLOATING
C1931 OUT_P.n573 GND 0.02fF $ **FLOATING
C1932 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11/GATE GND 0.01fF $ **FLOATING
C1933 OUT_P.n574 GND 0.01fF $ **FLOATING
C1934 OUT_P.n575 GND 0.01fF $ **FLOATING
C1935 OUT_P.n576 GND 0.01fF $ **FLOATING
C1936 OUT_P.n577 GND 0.01fF $ **FLOATING
C1937 OUT_P.n578 GND 0.01fF $ **FLOATING
C1938 OUT_P.n579 GND 0.18fF $ **FLOATING
C1939 OUT_P.n580 GND 0.03fF $ **FLOATING
C1940 OUT_P.n581 GND 0.03fF $ **FLOATING
C1941 OUT_P.n582 GND 0.00fF $ **FLOATING
C1942 OUT_P.n583 GND 0.01fF $ **FLOATING
C1943 OUT_P.n584 GND 0.01fF $ **FLOATING
C1944 OUT_P.n585 GND 0.02fF $ **FLOATING
C1945 OUT_P.n586 GND 0.02fF $ **FLOATING
C1946 OUT_P.n587 GND 0.01fF $ **FLOATING
C1947 OUT_P.n588 GND 0.05fF $ **FLOATING
C1948 OUT_P.n589 GND 0.04fF $ **FLOATING
C1949 OUT_P.n590 GND 0.01fF $ **FLOATING
C1950 OUT_P.n591 GND 0.01fF $ **FLOATING
C1951 OUT_P.n592 GND 0.02fF $ **FLOATING
C1952 OUT_P.n593 GND 0.02fF $ **FLOATING
C1953 OUT_P.n594 GND 0.01fF $ **FLOATING
C1954 OUT_P.n595 GND 0.01fF $ **FLOATING
C1955 OUT_P.n596 GND 0.01fF $ **FLOATING
C1956 OUT_P.n597 GND 0.01fF $ **FLOATING
C1957 OUT_P.n598 GND 0.03fF $ **FLOATING
C1958 OUT_P.n599 GND 0.01fF $ **FLOATING
C1959 OUT_P.n600 GND 0.01fF $ **FLOATING
C1960 OUT_P.n601 GND 0.01fF $ **FLOATING
C1961 OUT_P.n602 GND 0.01fF $ **FLOATING
C1962 OUT_P.n603 GND 0.01fF $ **FLOATING
C1963 OUT_P.n604 GND 0.01fF $ **FLOATING
C1964 OUT_P.n605 GND 0.01fF $ **FLOATING
C1965 OUT_P.n606 GND 0.01fF $ **FLOATING
C1966 OUT_P.n607 GND 0.01fF $ **FLOATING
C1967 OUT_P.n608 GND 0.01fF $ **FLOATING
C1968 OUT_P.n609 GND 0.02fF $ **FLOATING
C1969 OUT_P.n610 GND 0.01fF $ **FLOATING
C1970 OUT_P.n611 GND 0.01fF $ **FLOATING
C1971 OUT_P.n612 GND 0.01fF $ **FLOATING
C1972 OUT_P.n613 GND 0.18fF $ **FLOATING
C1973 OUT_P.n614 GND 0.03fF $ **FLOATING
C1974 OUT_P.n615 GND 0.03fF $ **FLOATING
C1975 OUT_P.n616 GND 0.00fF $ **FLOATING
C1976 OUT_P.n617 GND 0.01fF $ **FLOATING
C1977 OUT_P.n618 GND 0.01fF $ **FLOATING
C1978 OUT_P.n619 GND 0.02fF $ **FLOATING
C1979 vco_pair_base_0/rf_nfet_01v8_aM02W5p00L0p15_0/GATE GND 0.01fF $ **FLOATING
C1980 OUT_P.n620 GND 0.01fF $ **FLOATING
C1981 OUT_P.n621 GND 0.01fF $ **FLOATING
C1982 OUT_P.n622 GND 0.01fF $ **FLOATING
C1983 OUT_P.n623 GND 0.01fF $ **FLOATING
C1984 OUT_P.n624 GND 0.01fF $ **FLOATING
C1985 OUT_P.n625 GND 0.18fF $ **FLOATING
C1986 OUT_P.n626 GND 0.03fF $ **FLOATING
C1987 OUT_P.n627 GND 0.03fF $ **FLOATING
C1988 OUT_P.n628 GND 0.00fF $ **FLOATING
C1989 OUT_P.n629 GND 0.01fF $ **FLOATING
C1990 OUT_P.n630 GND 0.01fF $ **FLOATING
C1991 OUT_P.n631 GND 0.02fF $ **FLOATING
C1992 OUT_P.n632 GND 0.02fF $ **FLOATING
C1993 OUT_P.n633 GND 0.01fF $ **FLOATING
C1994 OUT_P.n634 GND 0.05fF $ **FLOATING
C1995 OUT_P.n635 GND 0.04fF $ **FLOATING
C1996 OUT_P.n636 GND 0.01fF $ **FLOATING
C1997 OUT_P.n637 GND 0.01fF $ **FLOATING
C1998 OUT_P.n638 GND 0.02fF $ **FLOATING
C1999 OUT_P.n639 GND 0.02fF $ **FLOATING
C2000 OUT_P.n640 GND 0.01fF $ **FLOATING
C2001 OUT_P.n641 GND 0.14fF $ **FLOATING
C2002 OUT_P.n642 GND 0.01fF $ **FLOATING
C2003 OUT_P.n643 GND 0.03fF $ **FLOATING
C2004 OUT_P.n644 GND 0.03fF $ **FLOATING
C2005 OUT_P.n645 GND 0.01fF $ **FLOATING
C2006 OUT_P.n646 GND 0.07fF $ **FLOATING
C2007 OUT_P.n647 GND 0.01fF $ **FLOATING
C2008 OUT_P.n648 GND 0.01fF $ **FLOATING
C2009 OUT_P.n649 GND 0.01fF $ **FLOATING
C2010 OUT_P.n650 GND 0.01fF $ **FLOATING
C2011 OUT_P.n651 GND 0.01fF $ **FLOATING
C2012 OUT_P.n652 GND 0.01fF $ **FLOATING
C2013 OUT_P.n653 GND 0.22fF $ **FLOATING
C2014 OUT_P.n654 GND 0.22fF $ **FLOATING
C2015 OUT_P.n655 GND 0.01fF $ **FLOATING
C2016 OUT_P.n656 GND 0.01fF $ **FLOATING
C2017 OUT_P.n657 GND 0.01fF $ **FLOATING
C2018 OUT_P.n658 GND 0.01fF $ **FLOATING
C2019 OUT_P.n659 GND 0.01fF $ **FLOATING
C2020 OUT_P.n660 GND 0.01fF $ **FLOATING
C2021 OUT_P.n661 GND 0.07fF $ **FLOATING
C2022 OUT_P.n662 GND 0.01fF $ **FLOATING
C2023 OUT_P.n663 GND 0.03fF $ **FLOATING
C2024 OUT_P.n664 GND 0.03fF $ **FLOATING
C2025 OUT_P.n665 GND 0.01fF $ **FLOATING
C2026 OUT_P.n666 GND 0.18fF $ **FLOATING
C2027 OUT_P.n667 GND 0.06fF $ **FLOATING
C2028 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1/GATE GND 0.00fF $ **FLOATING
C2029 OUT_P.n668 GND 0.01fF $ **FLOATING
C2030 OUT_P.n669 GND 0.01fF $ **FLOATING
C2031 OUT_P.n670 GND 0.01fF $ **FLOATING
C2032 OUT_P.n671 GND 0.01fF $ **FLOATING
C2033 OUT_P.n672 GND 0.01fF $ **FLOATING
C2034 OUT_P.n673 GND 0.00fF $ **FLOATING
C2035 OUT_P.n674 GND 0.18fF $ **FLOATING
C2036 OUT_P.n675 GND 0.03fF $ **FLOATING
C2037 OUT_P.n676 GND 0.03fF $ **FLOATING
C2038 OUT_P.n677 GND 0.00fF $ **FLOATING
C2039 OUT_P.n678 GND 0.01fF $ **FLOATING
C2040 OUT_P.n679 GND 0.01fF $ **FLOATING
C2041 OUT_P.n680 GND 0.02fF $ **FLOATING
C2042 OUT_P.n681 GND 0.02fF $ **FLOATING
C2043 OUT_P.n682 GND 0.01fF $ **FLOATING
C2044 OUT_P.n683 GND 0.05fF $ **FLOATING
C2045 OUT_P.n684 GND 0.04fF $ **FLOATING
C2046 OUT_P.n685 GND 0.01fF $ **FLOATING
C2047 OUT_P.n686 GND 0.00fF $ **FLOATING
C2048 OUT_P.n687 GND 0.01fF $ **FLOATING
C2049 OUT_P.n688 GND 0.01fF $ **FLOATING
C2050 OUT_P.n689 GND 0.02fF $ **FLOATING
C2051 OUT_P.n690 GND 0.03fF $ **FLOATING
C2052 OUT_P.n691 GND 0.06fF $ **FLOATING
C2053 OUT_P.n692 GND 0.06fF $ **FLOATING
C2054 OUT_P.n693 GND 0.01fF $ **FLOATING
C2055 OUT_P.n694 GND 0.01fF $ **FLOATING
C2056 OUT_P.n695 GND 0.00fF $ **FLOATING
C2057 OUT_P.n696 GND 0.01fF $ **FLOATING
C2058 OUT_P.n697 GND 0.01fF $ **FLOATING
C2059 OUT_P.n698 GND 0.01fF $ **FLOATING
C2060 OUT_P.n699 GND 0.01fF $ **FLOATING
C2061 OUT_P.n700 GND 0.01fF $ **FLOATING
C2062 OUT_P.n701 GND 0.01fF $ **FLOATING
C2063 OUT_P.n702 GND 0.26fF $ **FLOATING
C2064 OUT_P.n703 GND 0.26fF $ **FLOATING
C2065 OUT_P.n704 GND 0.01fF $ **FLOATING
C2066 OUT_P.n705 GND 0.01fF $ **FLOATING
C2067 OUT_P.n706 GND 0.03fF $ **FLOATING
C2068 OUT_P.n707 GND 0.03fF $ **FLOATING
C2069 OUT_P.n708 GND 0.01fF $ **FLOATING
C2070 OUT_P.n709 GND 0.07fF $ **FLOATING
C2071 OUT_P.n710 GND 0.01fF $ **FLOATING
C2072 OUT_P.n711 GND 0.01fF $ **FLOATING
C2073 OUT_P.n712 GND 0.01fF $ **FLOATING
C2074 OUT_P.n713 GND 0.01fF $ **FLOATING
C2075 OUT_P.n714 GND 0.01fF $ **FLOATING
C2076 OUT_P.n715 GND 0.01fF $ **FLOATING
C2077 OUT_P.n716 GND 0.22fF $ **FLOATING
C2078 OUT_P.n717 GND 0.22fF $ **FLOATING
C2079 OUT_P.n718 GND 0.01fF $ **FLOATING
C2080 OUT_P.n719 GND 0.01fF $ **FLOATING
C2081 OUT_P.n720 GND 0.01fF $ **FLOATING
C2082 OUT_P.n721 GND 0.01fF $ **FLOATING
C2083 OUT_P.n722 GND 0.01fF $ **FLOATING
C2084 OUT_P.n723 GND 0.01fF $ **FLOATING
C2085 OUT_P.n724 GND 0.07fF $ **FLOATING
C2086 OUT_P.n725 GND 0.01fF $ **FLOATING
C2087 OUT_P.n726 GND 0.03fF $ **FLOATING
C2088 OUT_P.n727 GND 0.03fF $ **FLOATING
C2089 OUT_P.n728 GND 0.01fF $ **FLOATING
C2090 OUT_P.n729 GND 0.01fF $ **FLOATING
C2091 OUT_P.n730 GND 0.26fF $ **FLOATING
C2092 OUT_P.n731 GND 0.26fF $ **FLOATING
C2093 OUT_P.n732 GND 0.01fF $ **FLOATING
C2094 OUT_P.n733 GND 0.01fF $ **FLOATING
C2095 OUT_P.n734 GND 0.03fF $ **FLOATING
C2096 OUT_P.n735 GND 0.03fF $ **FLOATING
C2097 OUT_P.n736 GND 0.01fF $ **FLOATING
C2098 OUT_P.n737 GND 0.07fF $ **FLOATING
C2099 OUT_P.n738 GND 0.01fF $ **FLOATING
C2100 OUT_P.n739 GND 0.01fF $ **FLOATING
C2101 OUT_P.n740 GND 0.01fF $ **FLOATING
C2102 OUT_P.n741 GND 0.01fF $ **FLOATING
C2103 OUT_P.n742 GND 0.01fF $ **FLOATING
C2104 OUT_P.n743 GND 0.01fF $ **FLOATING
C2105 OUT_P.n744 GND 0.22fF $ **FLOATING
C2106 OUT_P.n745 GND 0.22fF $ **FLOATING
C2107 OUT_P.n746 GND 0.01fF $ **FLOATING
C2108 OUT_P.n747 GND 0.01fF $ **FLOATING
C2109 OUT_P.n748 GND 0.01fF $ **FLOATING
C2110 OUT_P.n749 GND 0.01fF $ **FLOATING
C2111 OUT_P.n750 GND 0.01fF $ **FLOATING
C2112 OUT_P.n751 GND 0.01fF $ **FLOATING
C2113 OUT_P.n752 GND 0.07fF $ **FLOATING
C2114 OUT_P.n753 GND 0.01fF $ **FLOATING
C2115 OUT_P.n754 GND 0.03fF $ **FLOATING
C2116 OUT_P.n755 GND 0.03fF $ **FLOATING
C2117 OUT_P.n756 GND 0.01fF $ **FLOATING
C2118 OUT_P.n757 GND 0.01fF $ **FLOATING
C2119 OUT_P.n758 GND 0.26fF $ **FLOATING
C2120 OUT_P.n759 GND 0.26fF $ **FLOATING
C2121 OUT_P.n760 GND 0.01fF $ **FLOATING
C2122 OUT_P.n761 GND 0.01fF $ **FLOATING
C2123 OUT_P.n762 GND 0.01fF $ **FLOATING
C2124 OUT_P.n763 GND 0.04fF $ **FLOATING
C2125 OUT_P.n764 GND 0.01fF $ **FLOATING
C2126 OUT_P.n765 GND 0.01fF $ **FLOATING
C2127 OUT_P.n766 GND 0.01fF $ **FLOATING
C2128 OUT_P.n767 GND 0.01fF $ **FLOATING
C2129 OUT_P.n768 GND 0.01fF $ **FLOATING
C2130 OUT_P.n769 GND 0.03fF $ **FLOATING
C2131 OUT_P.n770 GND 0.03fF $ **FLOATING
C2132 OUT_P.n771 GND 0.01fF $ **FLOATING
C2133 OUT_P.n772 GND 0.18fF $ **FLOATING
C2134 OUT_P.n773 GND 0.06fF $ **FLOATING
C2135 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7/GATE GND 0.00fF $ **FLOATING
C2136 OUT_P.n774 GND 0.01fF $ **FLOATING
C2137 OUT_P.n775 GND 0.02fF $ **FLOATING
C2138 OUT_P.n776 GND 0.01fF $ **FLOATING
C2139 OUT_P.n777 GND 0.01fF $ **FLOATING
C2140 OUT_P.n778 GND 0.00fF $ **FLOATING
C2141 OUT_P.n779 GND 0.18fF $ **FLOATING
C2142 OUT_P.n780 GND 0.03fF $ **FLOATING
C2143 OUT_P.n781 GND 0.03fF $ **FLOATING
C2144 OUT_P.n782 GND 0.01fF $ **FLOATING
C2145 OUT_P.n783 GND 0.01fF $ **FLOATING
C2146 OUT_P.n784 GND 0.01fF $ **FLOATING
C2147 OUT_P.n785 GND 0.02fF $ **FLOATING
C2148 OUT_P.n786 GND 0.02fF $ **FLOATING
C2149 OUT_P.n787 GND 0.01fF $ **FLOATING
C2150 OUT_P.n788 GND 0.05fF $ **FLOATING
C2151 OUT_P.n789 GND 0.04fF $ **FLOATING
C2152 OUT_P.n790 GND 0.01fF $ **FLOATING
C2153 OUT_P.n791 GND 0.00fF $ **FLOATING
C2154 OUT_P.n792 GND 0.01fF $ **FLOATING
C2155 OUT_P.n793 GND 0.03fF $ **FLOATING
C2156 OUT_P.n794 GND 0.03fF $ **FLOATING
C2157 OUT_P.n795 GND 0.07fF $ **FLOATING
C2158 OUT_P.n796 GND 0.06fF $ **FLOATING
C2159 OUT_P.n797 GND 0.01fF $ **FLOATING
C2160 OUT_P.n798 GND 0.01fF $ **FLOATING
C2161 OUT_P.n799 GND 0.00fF $ **FLOATING
C2162 OUT_P.n800 GND 0.01fF $ **FLOATING
C2163 OUT_P.n801 GND 0.02fF $ **FLOATING
C2164 OUT_P.n802 GND 0.01fF $ **FLOATING
C2165 OUT_P.n803 GND 0.01fF $ **FLOATING
C2166 OUT_P.n804 GND 0.01fF $ **FLOATING
C2167 OUT_P.n805 GND 0.35fF $ **FLOATING
C2168 OUT_P.n806 GND 0.21fF $ **FLOATING
C2169 OUT_P.n807 GND 0.00fF $ **FLOATING
C2170 OUT_P.n808 GND 0.00fF $ **FLOATING
C2171 OUT_P.n809 GND 0.00fF $ **FLOATING
C2172 OUT_P.n810 GND 0.01fF $ **FLOATING
C2173 OUT_P.n811 GND 0.00fF $ **FLOATING
C2174 OUT_P.n812 GND 0.01fF $ **FLOATING
C2175 OUT_P.n813 GND 0.02fF $ **FLOATING
C2176 OUT_P.t5 GND 0.23fF
C2177 OUT_P.t0 GND 0.23fF
C2178 OUT_P.n814 GND 0.66fF $ **FLOATING
C2179 OUT_P.n815 GND 0.07fF $ **FLOATING
C2180 OUT_P.n816 GND 0.52fF $ **FLOATING
C2181 OUT_P.n817 GND 0.01fF $ **FLOATING
C2182 OUT_P.n818 GND 0.01fF $ **FLOATING
C2183 OUT_P.n819 GND 0.00fF $ **FLOATING
C2184 OUT_P.n820 GND 0.01fF $ **FLOATING
C2185 OUT_P.n821 GND 0.01fF $ **FLOATING
C2186 OUT_P.n822 GND 0.01fF $ **FLOATING
C2187 OUT_P.n823 GND 0.02fF $ **FLOATING
C2188 OUT_P.n824 GND 0.01fF $ **FLOATING
C2189 OUT_P.n825 GND 0.01fF $ **FLOATING
C2190 OUT_P.n826 GND 0.00fF $ **FLOATING
C2191 OUT_P.n827 GND 0.00fF $ **FLOATING
C2192 OUT_P.n828 GND 0.00fF $ **FLOATING
C2193 OUT_P.n829 GND 0.01fF $ **FLOATING
C2194 OUT_P.n830 GND 0.00fF $ **FLOATING
C2195 OUT_P.n831 GND 0.01fF $ **FLOATING
C2196 OUT_P.n832 GND 0.01fF $ **FLOATING
C2197 OUT_P.n833 GND 0.00fF $ **FLOATING
C2198 OUT_P.n834 GND 0.01fF $ **FLOATING
C2199 OUT_P.n835 GND 0.01fF $ **FLOATING
C2200 OUT_P.n836 GND 0.01fF $ **FLOATING
C2201 OUT_P.n837 GND 0.01fF $ **FLOATING
C2202 OUT_P.n838 GND 0.01fF $ **FLOATING
C2203 OUT_P.n839 GND 0.00fF $ **FLOATING
C2204 OUT_P.n840 GND 0.01fF $ **FLOATING
C2205 OUT_P.n841 GND 0.01fF $ **FLOATING
C2206 OUT_P.n842 GND 0.01fF $ **FLOATING
C2207 OUT_P.n843 GND 0.01fF $ **FLOATING
C2208 OUT_P.n844 GND 0.01fF $ **FLOATING
C2209 OUT_P.n845 GND 0.01fF $ **FLOATING
C2210 OUT_P.n846 GND 0.02fF $ **FLOATING
C2211 OUT_P.n847 GND 0.01fF $ **FLOATING
C2212 OUT_P.n848 GND 0.01fF $ **FLOATING
C2213 OUT_P.n849 GND 0.00fF $ **FLOATING
C2214 OUT_P.n850 GND 0.01fF $ **FLOATING
C2215 OUT_P.n851 GND 0.01fF $ **FLOATING
C2216 OUT_P.n852 GND 0.01fF $ **FLOATING
C2217 OUT_P.n853 GND 0.01fF $ **FLOATING
C2218 OUT_P.n854 GND 0.00fF $ **FLOATING
C2219 OUT_P.n855 GND 0.01fF $ **FLOATING
C2220 OUT_P.n856 GND 0.02fF $ **FLOATING
C2221 OUT_P.n857 GND 0.01fF $ **FLOATING
C2222 OUT_P.n858 GND 0.00fF $ **FLOATING
C2223 OUT_P.n859 GND 0.02fF $ **FLOATING
C2224 OUT_P.n860 GND 0.01fF $ **FLOATING
C2225 OUT_P.n861 GND 0.01fF $ **FLOATING
C2226 OUT_P.n862 GND 0.01fF $ **FLOATING
C2227 OUT_P.n863 GND 0.01fF $ **FLOATING
C2228 OUT_P.n864 GND 0.01fF $ **FLOATING
C2229 OUT_P.n865 GND 0.01fF $ **FLOATING
C2230 OUT_P.n866 GND 0.01fF $ **FLOATING
C2231 OUT_P.n867 GND 0.01fF $ **FLOATING
C2232 OUT_P.n868 GND 0.01fF $ **FLOATING
C2233 OUT_P.n869 GND 0.02fF $ **FLOATING
C2234 OUT_P.n870 GND 0.01fF $ **FLOATING
C2235 OUT_P.n871 GND 0.00fF $ **FLOATING
C2236 OUT_P.n872 GND 0.01fF $ **FLOATING
C2237 OUT_P.n873 GND 0.02fF $ **FLOATING
C2238 OUT_P.n874 GND 0.02fF $ **FLOATING
C2239 OUT_P.n875 GND 0.19fF $ **FLOATING
C2240 OUT_P.n876 GND 0.02fF $ **FLOATING
C2241 OUT_P.n877 GND 0.03fF $ **FLOATING
C2242 OUT_P.n878 GND 0.04fF $ **FLOATING
C2243 OUT_P.n879 GND 0.03fF $ **FLOATING
C2244 OUT_P.n881 GND 0.04fF $ **FLOATING
C2245 OUT_P.n882 GND 0.05fF $ **FLOATING
C2246 OUT_P.n883 GND 0.03fF $ **FLOATING
C2247 OUT_P.n884 GND 0.02fF $ **FLOATING
C2248 OUT_P.n885 GND 0.05fF $ **FLOATING
C2249 OUT_P.n886 GND 0.05fF $ **FLOATING
C2250 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12/DRAIN GND 0.09fF $ **FLOATING
C2251 OUT_P.n887 GND 0.10fF $ **FLOATING
C2252 OUT_P.n888 GND 0.05fF $ **FLOATING
C2253 OUT_P.n889 GND 0.08fF $ **FLOATING
C2254 OUT_P.n890 GND 0.08fF $ **FLOATING
C2255 OUT_P.n891 GND 0.08fF $ **FLOATING
C2256 OUT_P.n892 GND 0.08fF $ **FLOATING
C2257 OUT_P.n893 GND 0.08fF $ **FLOATING
C2258 OUT_P.n894 GND 0.05fF $ **FLOATING
C2259 OUT_P.n895 GND 0.09fF $ **FLOATING
C2260 OUT_P.n896 GND 0.10fF $ **FLOATING
C2261 OUT_P.n897 GND 0.05fF $ **FLOATING
C2262 OUT_P.n898 GND 0.07fF $ **FLOATING
C2263 OUT_P.n899 GND 0.08fF $ **FLOATING
C2264 OUT_P.n900 GND 0.05fF $ **FLOATING
C2265 OUT_P.n901 GND 0.05fF $ **FLOATING
C2266 OUT_P.n902 GND 1.34fF $ **FLOATING
C2267 OUT_P.n903 GND 0.16fF $ **FLOATING
C2268 OUT_P.n905 GND 0.12fF $ **FLOATING
C2269 OUT_P.n906 GND 0.99fF $ **FLOATING
C2270 OUT_P.n907 GND 1.02fF $ **FLOATING
C2271 OUT_P.n908 GND 0.00fF $ **FLOATING
C2272 OUT_P.n909 GND 0.00fF $ **FLOATING
C2273 OUT_P.n910 GND 0.00fF $ **FLOATING
C2274 OUT_P.n911 GND 0.00fF $ **FLOATING
C2275 OUT_P.n912 GND 0.01fF $ **FLOATING
C2276 OUT_P.n913 GND 0.00fF $ **FLOATING
C2277 OUT_P.n914 GND 0.01fF $ **FLOATING
C2278 OUT_P.n915 GND 0.02fF $ **FLOATING
C2279 OUT_P.t9 GND 0.23fF
C2280 OUT_P.t4 GND 0.23fF
C2281 OUT_P.n916 GND 0.66fF $ **FLOATING
C2282 OUT_P.n917 GND 0.07fF $ **FLOATING
C2283 OUT_P.n918 GND 0.52fF $ **FLOATING
C2284 OUT_P.n919 GND 0.01fF $ **FLOATING
C2285 OUT_P.n920 GND 0.01fF $ **FLOATING
C2286 OUT_P.n921 GND 0.00fF $ **FLOATING
C2287 OUT_P.n922 GND 0.01fF $ **FLOATING
C2288 OUT_P.n923 GND 0.01fF $ **FLOATING
C2289 OUT_P.n924 GND 0.01fF $ **FLOATING
C2290 OUT_P.n925 GND 0.02fF $ **FLOATING
C2291 OUT_P.n926 GND 0.01fF $ **FLOATING
C2292 OUT_P.n927 GND 0.01fF $ **FLOATING
C2293 OUT_P.n928 GND 0.00fF $ **FLOATING
C2294 OUT_P.n929 GND 0.00fF $ **FLOATING
C2295 OUT_P.n930 GND 0.00fF $ **FLOATING
C2296 OUT_P.n931 GND 0.01fF $ **FLOATING
C2297 OUT_P.n932 GND 0.01fF $ **FLOATING
C2298 OUT_P.n933 GND 0.01fF $ **FLOATING
C2299 OUT_P.n934 GND 0.00fF $ **FLOATING
C2300 OUT_P.n935 GND 0.01fF $ **FLOATING
C2301 OUT_P.n936 GND 0.01fF $ **FLOATING
C2302 OUT_P.n937 GND 0.01fF $ **FLOATING
C2303 OUT_P.n938 GND 0.01fF $ **FLOATING
C2304 OUT_P.n939 GND 0.01fF $ **FLOATING
C2305 OUT_P.n940 GND 0.00fF $ **FLOATING
C2306 OUT_P.n941 GND 0.01fF $ **FLOATING
C2307 OUT_P.n942 GND 0.00fF $ **FLOATING
C2308 OUT_P.n943 GND 0.01fF $ **FLOATING
C2309 OUT_P.n944 GND 0.01fF $ **FLOATING
C2310 OUT_P.n945 GND 0.01fF $ **FLOATING
C2311 OUT_P.n946 GND 0.01fF $ **FLOATING
C2312 OUT_P.n947 GND 0.01fF $ **FLOATING
C2313 OUT_P.n948 GND 0.02fF $ **FLOATING
C2314 OUT_P.n949 GND 0.01fF $ **FLOATING
C2315 OUT_P.n950 GND 0.01fF $ **FLOATING
C2316 OUT_P.n951 GND 0.00fF $ **FLOATING
C2317 OUT_P.n952 GND 0.01fF $ **FLOATING
C2318 OUT_P.n953 GND 0.01fF $ **FLOATING
C2319 OUT_P.n954 GND 0.01fF $ **FLOATING
C2320 OUT_P.n955 GND 0.01fF $ **FLOATING
C2321 OUT_P.n956 GND 0.00fF $ **FLOATING
C2322 OUT_P.n957 GND 0.01fF $ **FLOATING
C2323 OUT_P.n958 GND 0.02fF $ **FLOATING
C2324 OUT_P.n959 GND 0.01fF $ **FLOATING
C2325 OUT_P.n960 GND 0.00fF $ **FLOATING
C2326 OUT_P.n961 GND 0.02fF $ **FLOATING
C2327 OUT_P.n962 GND 0.01fF $ **FLOATING
C2328 OUT_P.n963 GND 0.01fF $ **FLOATING
C2329 OUT_P.n964 GND 0.01fF $ **FLOATING
C2330 OUT_P.n965 GND 0.01fF $ **FLOATING
C2331 OUT_P.n966 GND 0.01fF $ **FLOATING
C2332 OUT_P.n967 GND 0.01fF $ **FLOATING
C2333 OUT_P.n968 GND 0.01fF $ **FLOATING
C2334 OUT_P.n969 GND 0.01fF $ **FLOATING
C2335 OUT_P.n970 GND 0.01fF $ **FLOATING
C2336 OUT_P.n971 GND 0.02fF $ **FLOATING
C2337 OUT_P.n972 GND 0.01fF $ **FLOATING
C2338 OUT_P.n973 GND 0.01fF $ **FLOATING
C2339 OUT_P.n974 GND 0.02fF $ **FLOATING
C2340 OUT_P.n975 GND 0.02fF $ **FLOATING
C2341 OUT_P.n976 GND 0.19fF $ **FLOATING
C2342 OUT_P.n977 GND 0.02fF $ **FLOATING
C2343 OUT_P.n978 GND 0.03fF $ **FLOATING
C2344 OUT_P.n979 GND 0.04fF $ **FLOATING
C2345 OUT_P.n980 GND 0.02fF $ **FLOATING
C2346 OUT_P.n982 GND 0.04fF $ **FLOATING
C2347 OUT_P.n983 GND 0.05fF $ **FLOATING
C2348 OUT_P.n984 GND 0.03fF $ **FLOATING
C2349 OUT_P.n985 GND 0.02fF $ **FLOATING
C2350 OUT_P.n986 GND 0.05fF $ **FLOATING
C2351 OUT_P.n987 GND 0.05fF $ **FLOATING
C2352 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10/DRAIN GND 0.09fF $ **FLOATING
C2353 OUT_P.n988 GND 0.10fF $ **FLOATING
C2354 OUT_P.n989 GND 0.05fF $ **FLOATING
C2355 OUT_P.n990 GND 0.08fF $ **FLOATING
C2356 OUT_P.n991 GND 0.08fF $ **FLOATING
C2357 OUT_P.n992 GND 0.08fF $ **FLOATING
C2358 OUT_P.n993 GND 0.08fF $ **FLOATING
C2359 OUT_P.n994 GND 0.08fF $ **FLOATING
C2360 OUT_P.n995 GND 0.05fF $ **FLOATING
C2361 OUT_P.n996 GND 0.09fF $ **FLOATING
C2362 OUT_P.n997 GND 0.10fF $ **FLOATING
C2363 OUT_P.n998 GND 0.05fF $ **FLOATING
C2364 OUT_P.n999 GND 0.07fF $ **FLOATING
C2365 OUT_P.n1000 GND 0.08fF $ **FLOATING
C2366 OUT_P.n1001 GND 0.05fF $ **FLOATING
C2367 OUT_P.n1002 GND 0.05fF $ **FLOATING
C2368 OUT_P.n1004 GND 0.16fF $ **FLOATING
C2369 OUT_P.n1006 GND 0.12fF $ **FLOATING
C2370 OUT_P.n1007 GND 0.99fF $ **FLOATING
C2371 OUT_P.n1008 GND 1.02fF $ **FLOATING
C2372 OUT_P.n1009 GND 0.00fF $ **FLOATING
C2373 OUT_P.n1010 GND 0.00fF $ **FLOATING
C2374 OUT_P.n1011 GND 0.00fF $ **FLOATING
C2375 OUT_P.n1012 GND 0.00fF $ **FLOATING
C2376 OUT_P.n1013 GND 0.01fF $ **FLOATING
C2377 OUT_P.n1014 GND 0.00fF $ **FLOATING
C2378 OUT_P.n1015 GND 0.01fF $ **FLOATING
C2379 OUT_P.n1016 GND 0.02fF $ **FLOATING
C2380 OUT_P.t12 GND 0.23fF
C2381 OUT_P.t2 GND 0.23fF
C2382 OUT_P.n1017 GND 0.66fF $ **FLOATING
C2383 OUT_P.n1018 GND 0.07fF $ **FLOATING
C2384 OUT_P.n1019 GND 0.52fF $ **FLOATING
C2385 OUT_P.n1020 GND 0.01fF $ **FLOATING
C2386 OUT_P.n1021 GND 0.01fF $ **FLOATING
C2387 OUT_P.n1022 GND 0.00fF $ **FLOATING
C2388 OUT_P.n1023 GND 0.01fF $ **FLOATING
C2389 OUT_P.n1024 GND 0.01fF $ **FLOATING
C2390 OUT_P.n1025 GND 0.01fF $ **FLOATING
C2391 OUT_P.n1026 GND 0.02fF $ **FLOATING
C2392 OUT_P.n1027 GND 0.01fF $ **FLOATING
C2393 OUT_P.n1028 GND 0.01fF $ **FLOATING
C2394 OUT_P.n1029 GND 0.00fF $ **FLOATING
C2395 OUT_P.n1030 GND 0.00fF $ **FLOATING
C2396 OUT_P.n1031 GND 0.00fF $ **FLOATING
C2397 OUT_P.n1032 GND 0.01fF $ **FLOATING
C2398 OUT_P.n1033 GND 0.01fF $ **FLOATING
C2399 OUT_P.n1034 GND 0.01fF $ **FLOATING
C2400 OUT_P.n1035 GND 0.00fF $ **FLOATING
C2401 OUT_P.n1036 GND 0.01fF $ **FLOATING
C2402 OUT_P.n1037 GND 0.01fF $ **FLOATING
C2403 OUT_P.n1038 GND 0.01fF $ **FLOATING
C2404 OUT_P.n1039 GND 0.01fF $ **FLOATING
C2405 OUT_P.n1040 GND 0.01fF $ **FLOATING
C2406 OUT_P.n1041 GND 0.00fF $ **FLOATING
C2407 OUT_P.n1042 GND 0.01fF $ **FLOATING
C2408 OUT_P.n1043 GND 0.00fF $ **FLOATING
C2409 OUT_P.n1044 GND 0.01fF $ **FLOATING
C2410 OUT_P.n1045 GND 0.01fF $ **FLOATING
C2411 OUT_P.n1046 GND 0.01fF $ **FLOATING
C2412 OUT_P.n1047 GND 0.01fF $ **FLOATING
C2413 OUT_P.n1048 GND 0.01fF $ **FLOATING
C2414 OUT_P.n1049 GND 0.02fF $ **FLOATING
C2415 OUT_P.n1050 GND 0.01fF $ **FLOATING
C2416 OUT_P.n1051 GND 0.01fF $ **FLOATING
C2417 OUT_P.n1052 GND 0.00fF $ **FLOATING
C2418 OUT_P.n1053 GND 0.01fF $ **FLOATING
C2419 OUT_P.n1054 GND 0.01fF $ **FLOATING
C2420 OUT_P.n1055 GND 0.01fF $ **FLOATING
C2421 OUT_P.n1056 GND 0.01fF $ **FLOATING
C2422 OUT_P.n1057 GND 0.00fF $ **FLOATING
C2423 OUT_P.n1058 GND 0.01fF $ **FLOATING
C2424 OUT_P.n1059 GND 0.02fF $ **FLOATING
C2425 OUT_P.n1060 GND 0.01fF $ **FLOATING
C2426 OUT_P.n1061 GND 0.00fF $ **FLOATING
C2427 OUT_P.n1062 GND 0.02fF $ **FLOATING
C2428 OUT_P.n1063 GND 0.01fF $ **FLOATING
C2429 OUT_P.n1064 GND 0.01fF $ **FLOATING
C2430 OUT_P.n1065 GND 0.01fF $ **FLOATING
C2431 OUT_P.n1066 GND 0.01fF $ **FLOATING
C2432 OUT_P.n1067 GND 0.01fF $ **FLOATING
C2433 OUT_P.n1068 GND 0.01fF $ **FLOATING
C2434 OUT_P.n1069 GND 0.01fF $ **FLOATING
C2435 OUT_P.n1070 GND 0.01fF $ **FLOATING
C2436 OUT_P.n1071 GND 0.01fF $ **FLOATING
C2437 OUT_P.n1072 GND 0.02fF $ **FLOATING
C2438 OUT_P.n1073 GND 0.01fF $ **FLOATING
C2439 OUT_P.n1074 GND 0.01fF $ **FLOATING
C2440 OUT_P.n1075 GND 0.02fF $ **FLOATING
C2441 OUT_P.n1076 GND 0.02fF $ **FLOATING
C2442 OUT_P.n1077 GND 0.19fF $ **FLOATING
C2443 OUT_P.n1078 GND 0.02fF $ **FLOATING
C2444 OUT_P.n1079 GND 0.03fF $ **FLOATING
C2445 OUT_P.n1080 GND 0.04fF $ **FLOATING
C2446 OUT_P.n1081 GND 0.02fF $ **FLOATING
C2447 OUT_P.n1083 GND 0.04fF $ **FLOATING
C2448 OUT_P.n1084 GND 0.05fF $ **FLOATING
C2449 OUT_P.n1085 GND 0.03fF $ **FLOATING
C2450 OUT_P.n1086 GND 0.02fF $ **FLOATING
C2451 OUT_P.n1087 GND 0.05fF $ **FLOATING
C2452 OUT_P.n1088 GND 0.05fF $ **FLOATING
C2453 vco_pair_base_0/sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8/DRAIN GND 0.09fF $ **FLOATING
C2454 OUT_P.n1089 GND 0.10fF $ **FLOATING
C2455 OUT_P.n1090 GND 0.05fF $ **FLOATING
C2456 OUT_P.n1091 GND 0.08fF $ **FLOATING
C2457 OUT_P.n1092 GND 0.08fF $ **FLOATING
C2458 OUT_P.n1093 GND 0.08fF $ **FLOATING
C2459 OUT_P.n1094 GND 0.08fF $ **FLOATING
C2460 OUT_P.n1095 GND 0.08fF $ **FLOATING
C2461 OUT_P.n1096 GND 0.05fF $ **FLOATING
C2462 OUT_P.n1097 GND 0.09fF $ **FLOATING
C2463 OUT_P.n1098 GND 0.10fF $ **FLOATING
C2464 OUT_P.n1099 GND 0.05fF $ **FLOATING
C2465 OUT_P.n1100 GND 0.07fF $ **FLOATING
C2466 OUT_P.n1101 GND 0.08fF $ **FLOATING
C2467 OUT_P.n1102 GND 0.05fF $ **FLOATING
C2468 OUT_P.n1103 GND 0.05fF $ **FLOATING
C2469 OUT_P.n1105 GND 0.16fF $ **FLOATING
C2470 OUT_P.n1107 GND 0.12fF $ **FLOATING
C2471 OUT_P.n1108 GND 1.53fF $ **FLOATING
C2472 OUT_P.n1109 GND 1.51fF $ **FLOATING
C2473 OUT_P.n1110 GND 0.35fF $ **FLOATING
C2474 OUT_P.n1111 GND 0.44fF $ **FLOATING
C2475 OUT_P.n1112 GND 0.03fF $ **FLOATING
C2476 OUT_P.n1113 GND 0.00fF $ **FLOATING
C2477 OUT_P.n1114 GND 0.00fF $ **FLOATING
C2478 OUT_P.n1115 GND 0.01fF $ **FLOATING
C2479 OUT_P.n1116 GND 0.02fF $ **FLOATING
C2480 OUT_P.n1117 GND 0.02fF $ **FLOATING
C2481 OUT_P.n1118 GND 0.02fF $ **FLOATING
C2482 OUT_P.n1119 GND 0.02fF $ **FLOATING
C2483 OUT_P.n1120 GND 0.02fF $ **FLOATING
C2484 OUT_P.n1121 GND 0.01fF $ **FLOATING
C2485 OUT_P.n1122 GND 0.01fF $ **FLOATING
C2486 OUT_P.n1123 GND 0.11fF $ **FLOATING
C2487 OUT_P.n1124 GND 0.06fF $ **FLOATING
C2488 OUT_P.t21 GND 0.25fF
C2489 OUT_P.n1125 GND 0.18fF $ **FLOATING
C2490 OUT_P.n1126 GND 0.06fF $ **FLOATING
C2491 OUT_P.n1127 GND 0.02fF $ **FLOATING
C2492 OUT_P.t19 GND 0.25fF
C2493 OUT_P.n1128 GND 0.18fF $ **FLOATING
C2494 OUT_P.n1129 GND 0.03fF $ **FLOATING
C2495 OUT_P.n1130 GND 0.04fF $ **FLOATING
C2496 OUT_P.n1131 GND 0.01fF $ **FLOATING
C2497 OUT_P.n1132 GND 0.01fF $ **FLOATING
C2498 OUT_P.n1133 GND 0.00fF $ **FLOATING
C2499 OUT_P.n1134 GND 0.01fF $ **FLOATING
C2500 OUT_P.n1135 GND 0.03fF $ **FLOATING
C2501 OUT_P.n1136 GND 0.03fF $ **FLOATING
C2502 OUT_P.n1137 GND 0.05fF $ **FLOATING
C2503 OUT_P.n1138 GND 0.04fF $ **FLOATING
C2504 OUT_P.n1139 GND 0.02fF $ **FLOATING
C2505 OUT_P.n1140 GND 0.03fF $ **FLOATING
C2506 OUT_P.n1141 GND 0.03fF $ **FLOATING
C2507 OUT_P.n1142 GND 0.06fF $ **FLOATING
C2508 OUT_P.n1143 GND 0.04fF $ **FLOATING
C2509 OUT_P.n1144 GND 0.01fF $ **FLOATING
C2510 OUT_P.n1145 GND 0.02fF $ **FLOATING
C2511 OUT_P.n1146 GND 0.36fF $ **FLOATING
C2512 OUT_P.n1147 GND 0.36fF $ **FLOATING
C2513 OUT_P.n1148 GND 0.02fF $ **FLOATING
C2514 OUT_P.n1149 GND 0.01fF $ **FLOATING
C2515 OUT_P.n1150 GND 0.03fF $ **FLOATING
C2516 OUT_P.n1151 GND 0.00fF $ **FLOATING
C2517 OUT_P.n1152 GND 0.00fF $ **FLOATING
C2518 OUT_P.n1153 GND 0.01fF $ **FLOATING
C2519 OUT_P.n1154 GND 0.02fF $ **FLOATING
C2520 OUT_P.n1155 GND 0.06fF $ **FLOATING
C2521 OUT_P.n1156 GND 0.06fF $ **FLOATING
C2522 OUT_P.n1157 GND 0.02fF $ **FLOATING
C2523 OUT_P.t15 GND 0.25fF
C2524 OUT_P.n1158 GND 0.18fF $ **FLOATING
C2525 OUT_P.n1159 GND 0.03fF $ **FLOATING
C2526 OUT_P.n1160 GND 0.04fF $ **FLOATING
C2527 OUT_P.n1161 GND 0.01fF $ **FLOATING
C2528 OUT_P.n1162 GND 0.01fF $ **FLOATING
C2529 OUT_P.n1163 GND 0.00fF $ **FLOATING
C2530 OUT_P.n1164 GND 0.01fF $ **FLOATING
C2531 OUT_P.n1165 GND 0.03fF $ **FLOATING
C2532 OUT_P.n1166 GND 0.03fF $ **FLOATING
C2533 OUT_P.n1167 GND 0.05fF $ **FLOATING
C2534 OUT_P.n1168 GND 0.04fF $ **FLOATING
C2535 OUT_P.n1169 GND 0.02fF $ **FLOATING
C2536 OUT_P.n1170 GND 0.03fF $ **FLOATING
C2537 OUT_P.n1171 GND 0.03fF $ **FLOATING
C2538 OUT_P.t18 GND 0.25fF
C2539 OUT_P.n1172 GND 0.18fF $ **FLOATING
C2540 OUT_P.n1173 GND 0.06fF $ **FLOATING
C2541 OUT_P.n1174 GND 0.06fF $ **FLOATING
C2542 OUT_P.n1175 GND 0.04fF $ **FLOATING
C2543 OUT_P.n1176 GND 0.02fF $ **FLOATING
C2544 OUT_P.n1177 GND 0.02fF $ **FLOATING
C2545 OUT_P.n1178 GND 0.02fF $ **FLOATING
C2546 OUT_P.n1179 GND 0.02fF $ **FLOATING
C2547 OUT_P.n1180 GND 0.01fF $ **FLOATING
C2548 OUT_P.n1181 GND 0.01fF $ **FLOATING
C2549 OUT_P.n1182 GND 0.02fF $ **FLOATING
C2550 OUT_P.n1183 GND 0.36fF $ **FLOATING
C2551 OUT_P.n1184 GND 0.36fF $ **FLOATING
C2552 OUT_P.n1185 GND 0.02fF $ **FLOATING
C2553 OUT_P.n1186 GND 0.01fF $ **FLOATING
C2554 OUT_P.n1187 GND 0.03fF $ **FLOATING
C2555 OUT_P.n1188 GND 0.00fF $ **FLOATING
C2556 OUT_P.n1189 GND 0.00fF $ **FLOATING
C2557 OUT_P.n1190 GND 0.01fF $ **FLOATING
C2558 OUT_P.n1191 GND 0.02fF $ **FLOATING
C2559 OUT_P.n1192 GND 0.06fF $ **FLOATING
C2560 OUT_P.n1193 GND 0.06fF $ **FLOATING
C2561 OUT_P.n1194 GND 0.02fF $ **FLOATING
C2562 OUT_P.t20 GND 0.25fF
C2563 OUT_P.n1195 GND 0.18fF $ **FLOATING
C2564 OUT_P.n1196 GND 0.03fF $ **FLOATING
C2565 OUT_P.n1197 GND 0.04fF $ **FLOATING
C2566 OUT_P.n1198 GND 0.01fF $ **FLOATING
C2567 OUT_P.n1199 GND 0.01fF $ **FLOATING
C2568 OUT_P.n1200 GND 0.00fF $ **FLOATING
C2569 OUT_P.n1201 GND 0.01fF $ **FLOATING
C2570 OUT_P.n1202 GND 0.03fF $ **FLOATING
C2571 OUT_P.n1203 GND 0.03fF $ **FLOATING
C2572 OUT_P.n1204 GND 0.05fF $ **FLOATING
C2573 OUT_P.n1205 GND 0.04fF $ **FLOATING
C2574 OUT_P.n1206 GND 0.02fF $ **FLOATING
C2575 OUT_P.n1207 GND 0.03fF $ **FLOATING
C2576 OUT_P.n1208 GND 0.03fF $ **FLOATING
C2577 OUT_P.t26 GND 0.25fF
C2578 OUT_P.n1209 GND 0.18fF $ **FLOATING
C2579 OUT_P.n1210 GND 0.06fF $ **FLOATING
C2580 OUT_P.n1211 GND 0.06fF $ **FLOATING
C2581 OUT_P.n1212 GND 0.04fF $ **FLOATING
C2582 OUT_P.n1213 GND 0.02fF $ **FLOATING
C2583 OUT_P.n1214 GND 0.02fF $ **FLOATING
C2584 OUT_P.n1215 GND 0.02fF $ **FLOATING
C2585 OUT_P.n1216 GND 0.02fF $ **FLOATING
C2586 OUT_P.n1217 GND 0.01fF $ **FLOATING
C2587 OUT_P.n1218 GND 0.01fF $ **FLOATING
C2588 OUT_P.n1219 GND 0.02fF $ **FLOATING
C2589 OUT_P.n1220 GND 0.36fF $ **FLOATING
C2590 OUT_P.n1221 GND 0.36fF $ **FLOATING
C2591 OUT_P.n1222 GND 0.02fF $ **FLOATING
C2592 OUT_P.n1223 GND 0.01fF $ **FLOATING
C2593 OUT_P.n1224 GND 0.03fF $ **FLOATING
C2594 OUT_P.n1225 GND 0.00fF $ **FLOATING
C2595 OUT_P.n1226 GND 0.00fF $ **FLOATING
C2596 OUT_P.n1227 GND 0.01fF $ **FLOATING
C2597 OUT_P.n1228 GND 0.02fF $ **FLOATING
C2598 OUT_P.n1229 GND 0.06fF $ **FLOATING
C2599 OUT_P.n1230 GND 0.06fF $ **FLOATING
C2600 OUT_P.n1231 GND 0.05fF $ **FLOATING
C2601 OUT_P.n1232 GND 0.04fF $ **FLOATING
C2602 OUT_P.t22 GND 0.25fF
C2603 OUT_P.n1233 GND 0.18fF $ **FLOATING
C2604 OUT_P.n1234 GND 0.03fF $ **FLOATING
C2605 OUT_P.n1235 GND 0.04fF $ **FLOATING
C2606 OUT_P.n1236 GND 0.02fF $ **FLOATING
C2607 OUT_P.n1237 GND 0.01fF $ **FLOATING
C2608 OUT_P.n1238 GND 0.01fF $ **FLOATING
C2609 OUT_P.n1239 GND 0.00fF $ **FLOATING
C2610 OUT_P.n1240 GND 0.01fF $ **FLOATING
C2611 OUT_P.n1241 GND 0.03fF $ **FLOATING
C2612 OUT_P.n1242 GND 0.03fF $ **FLOATING
C2613 OUT_P.n1243 GND 0.02fF $ **FLOATING
C2614 OUT_P.n1244 GND 0.03fF $ **FLOATING
C2615 OUT_P.n1245 GND 0.03fF $ **FLOATING
C2616 OUT_P.t17 GND 0.25fF
C2617 OUT_P.n1246 GND 0.18fF $ **FLOATING
C2618 OUT_P.n1247 GND 0.06fF $ **FLOATING
C2619 OUT_P.n1248 GND 0.06fF $ **FLOATING
C2620 OUT_P.n1249 GND 0.04fF $ **FLOATING
C2621 OUT_P.n1250 GND 0.02fF $ **FLOATING
C2622 OUT_P.n1251 GND 0.02fF $ **FLOATING
C2623 OUT_P.n1252 GND 0.02fF $ **FLOATING
C2624 OUT_P.n1253 GND 0.02fF $ **FLOATING
C2625 OUT_P.n1254 GND 0.01fF $ **FLOATING
C2626 OUT_P.n1255 GND 0.01fF $ **FLOATING
C2627 OUT_P.n1256 GND 0.02fF $ **FLOATING
C2628 OUT_P.n1257 GND 1.14fF $ **FLOATING
C2629 OUT_P.n1258 GND 2.83fF $ **FLOATING
C2630 OUT_P.n1260 GND 0.23fF $ **FLOATING
C2631 OUT_P.n1261 GND 1.09fF $ **FLOATING
C2632 OUT_P.n1262 GND 1.09fF $ **FLOATING
C2633 OUT_P.n1264 GND 3.07fF $ **FLOATING
C2634 OUT_P.n1265 GND 1.35fF $ **FLOATING
C2635 OUT_P.t24 GND 0.25fF
C2636 OUT_P.n1266 GND 0.18fF $ **FLOATING
C2637 OUT_P.n1267 GND 0.06fF $ **FLOATING
C2638 OUT_P.n1268 GND 0.02fF $ **FLOATING
C2639 OUT_P.t14 GND 0.25fF
C2640 OUT_P.n1269 GND 0.18fF $ **FLOATING
C2641 OUT_P.n1270 GND 0.03fF $ **FLOATING
C2642 OUT_P.n1271 GND 0.04fF $ **FLOATING
C2643 OUT_P.n1272 GND 0.01fF $ **FLOATING
C2644 OUT_P.n1273 GND 0.01fF $ **FLOATING
C2645 OUT_P.n1274 GND 0.01fF $ **FLOATING
C2646 OUT_P.n1275 GND 0.03fF $ **FLOATING
C2647 OUT_P.n1276 GND 0.03fF $ **FLOATING
C2648 OUT_P.n1277 GND 0.05fF $ **FLOATING
C2649 OUT_P.n1278 GND 0.04fF $ **FLOATING
C2650 OUT_P.n1279 GND 0.02fF $ **FLOATING
C2651 OUT_P.n1280 GND 0.03fF $ **FLOATING
C2652 OUT_P.n1281 GND 0.03fF $ **FLOATING
C2653 OUT_P.n1282 GND 0.06fF $ **FLOATING
C2654 OUT_P.n1283 GND 0.14fF $ **FLOATING
C2655 OUT_P.n1284 GND 0.07fF $ **FLOATING
C2656 OUT_P.n1285 GND 0.08fF $ **FLOATING
C2657 OUT_P.n1286 GND 0.07fF $ **FLOATING
C2658 OUT_P.n1287 GND 0.08fF $ **FLOATING
C2659 OUT_P.n1288 GND 0.07fF $ **FLOATING
C2660 OUT_P.n1289 GND 0.10fF $ **FLOATING
C2661 OUT_P.n1290 GND 0.01fF $ **FLOATING
C2662 OUT_P.n1291 GND 0.03fF $ **FLOATING
C2663 OUT_P.n1292 GND 0.43fF $ **FLOATING
C2664 OUT_P.n1293 GND 0.43fF $ **FLOATING
C2665 OUT_P.t25 GND 0.25fF
C2666 OUT_P.n1294 GND 0.18fF $ **FLOATING
C2667 OUT_P.n1295 GND 0.06fF $ **FLOATING
C2668 OUT_P.n1296 GND 0.02fF $ **FLOATING
C2669 OUT_P.t23 GND 0.25fF
C2670 OUT_P.n1297 GND 0.18fF $ **FLOATING
C2671 OUT_P.n1298 GND 0.03fF $ **FLOATING
C2672 OUT_P.n1299 GND 0.04fF $ **FLOATING
C2673 OUT_P.n1300 GND 0.01fF $ **FLOATING
C2674 OUT_P.n1301 GND 0.01fF $ **FLOATING
C2675 OUT_P.n1302 GND 0.01fF $ **FLOATING
C2676 OUT_P.n1303 GND 0.03fF $ **FLOATING
C2677 OUT_P.n1304 GND 0.03fF $ **FLOATING
C2678 OUT_P.n1305 GND 0.05fF $ **FLOATING
C2679 OUT_P.n1306 GND 0.04fF $ **FLOATING
C2680 OUT_P.n1307 GND 0.02fF $ **FLOATING
C2681 OUT_P.n1308 GND 0.03fF $ **FLOATING
C2682 OUT_P.n1309 GND 0.03fF $ **FLOATING
C2683 OUT_P.n1310 GND 0.06fF $ **FLOATING
C2684 OUT_P.n1311 GND 0.14fF $ **FLOATING
C2685 OUT_P.n1312 GND 0.07fF $ **FLOATING
C2686 OUT_P.n1313 GND 0.08fF $ **FLOATING
C2687 OUT_P.n1314 GND 0.07fF $ **FLOATING
C2688 OUT_P.n1315 GND 0.08fF $ **FLOATING
C2689 OUT_P.n1316 GND 0.07fF $ **FLOATING
C2690 OUT_P.n1317 GND 0.10fF $ **FLOATING
C2691 OUT_P.n1318 GND 0.01fF $ **FLOATING
C2692 OUT_P.n1319 GND 0.03fF $ **FLOATING
C2693 OUT_P.n1320 GND 0.43fF $ **FLOATING
C2694 OUT_P.n1321 GND 0.54fF $ **FLOATING
C2695 OUT_P.n1322 GND 0.14fF $ **FLOATING
C2696 OUT_P.t16 GND 0.25fF
C2697 OUT_P.n1323 GND 0.18fF $ **FLOATING
C2698 OUT_P.n1324 GND 0.06fF $ **FLOATING
C2699 OUT_P.n1325 GND 0.06fF $ **FLOATING
C2700 OUT_P.n1326 GND 0.03fF $ **FLOATING
C2701 OUT_P.n1327 GND 0.03fF $ **FLOATING
C2702 OUT_P.n1328 GND 0.05fF $ **FLOATING
C2703 OUT_P.n1329 GND 0.04fF $ **FLOATING
C2704 OUT_P.n1330 GND 0.02fF $ **FLOATING
C2705 OUT_P.n1331 GND 0.03fF $ **FLOATING
C2706 OUT_P.n1332 GND 0.03fF $ **FLOATING
C2707 OUT_P.n1333 GND 0.01fF $ **FLOATING
C2708 OUT_P.n1334 GND 0.01fF $ **FLOATING
C2709 OUT_P.n1335 GND 0.01fF $ **FLOATING
C2710 OUT_P.n1336 GND 0.02fF $ **FLOATING
.ends

