** sch_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_wo_ind_tb.sch
**.subckt vco_wo_ind_tb
V1 VDD GND 1.8
Vbit0 net1 GND 0
Vbit1 net2 GND 0
Vbit2 net3 GND 0
Vbit3 net4 GND 0
Vbit4 net5 GND 0
Vbit5 net6 GND 0
Vtune net8 GND 1.8
L1 net7 OUTP 1.1n m=1
L2 net7 OUTN 1.1n m=1
R1 OUTN OUTP 350 m=1
R2 BUFN BUFP 100 m=1
C1 BUFP GND 50f m=1
C2 BUFN GND 50f m=1
E1 BUFOUT GND BUFP BUFN 1
E2 VCOOUT GND OUTP OUTN 1
X1 OUTP GND net7 VDD OUTN net1 net2 net3 net4 net5 net6 GND net8 BUFP BUFN VDD vco_wo_ind
**** begin user architecture code


.save BUFOUT
.control
    *intial value of code sweeps
    let code = 63 
    let j = 0
    let start_vtune = 0
    let end_vtune = 1.8
    let delta_vtune = 0.1
    let vtune_act = start_vtune
    
    *creating plot to store amplitude and freq data
    setplot new
    set scratch = $curplot 
    set curplottitle = "Frequency and Amplitude for each code"
    let vtune_scale = delta_vtune*vector(19) $ x axis of lot
    settype voltage vtune_scale
    *let freq = vector(1216)
    let freq = unitvec(19)
    *reshape freq [64][19]
    settype frequency freq
    *let amplitude = vector(1216)
    let amplitude = unitvec(19)
    *reshape amplitude [64][19]
    settype voltage amplitude

    *setting printing data
    set wr_singlescale
    set wr_vecnames

    while code < 64
    * setting the cap bank code
        while vtune_act <= end_vtune
            *do tran sim
            alter Vtune vtune_act
            tran 100p 85n 50n
            meas tran period trig bufout val=50m rise=1 targ bufout val=50m rise=2 $ measuring period
            let {$scratch}.freq[j] = 1/period
            let {$scratch}.amplitude[j] = vecmax(bufout)
            let j = j + 1
            let vtune_act = vtune_act + delta_vtune
            wrdata data.csv {$scratch}.freq {$scratch}.amplitude
        end
        *reset variables
        let vtune_act = start_vtune
        let j = 0
        let code = code + 1
    end

    *plotting
    setplot {$scratch}
    plot freq
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/shpeccy/ntfs_drive/Linux_Programs/skywater-pdk/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/shpeccy/ntfs_drive/Linux_Programs/skywater-pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/shpeccy/ntfs_drive/Linux_Programs/skywater-pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/shpeccy/ntfs_drive/Linux_Programs/skywater-pdk/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  vco_wo_ind.sym # of pins=16
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_wo_ind.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_wo_ind.sch
.subckt vco_wo_ind  OUT_P GND IND_CT VDD OUT_N freq<0> freq<1> freq<2> freq<3> freq<4> freq<5> VBIAS
+ Vtune BUF_P BUF_N VBIAS_BUF
*.iopin OUT_P
*.iopin IND_CT
*.iopin Vtune
*.ipin freq<0>
*.ipin freq<1>
*.ipin freq<2>
*.ipin freq<3>
*.ipin freq<4>
*.ipin freq<5>
*.iopin GND
*.opin BUF_P
*.opin BUF_N
*.iopin OUT_N
*.iopin VBIAS_BUF
*.iopin VDD
*.iopin VBIAS
X1 OUT_P OUT_N GND Vtune cap_var
X2 OUT_P OUT_N VDD GND freq<0> freq<1> freq<2> freq<3> freq<4> freq<5> capbank
XC1 OUT_P OUT_N sky130_fd_pr__cap_mim_m3_1 W=13.3 L=13.3 MF=1 m=1
R2 net1 VBIAS_BUF sky130_fd_pr__res_generic_po W=1 L=6 m=1
x1 VDD IND_CT GND VBIAS vco_pmirr
x2 OUT_P OUT_N GND vco_pair
X3 net1 VDD GND BUF_N BUF_P OUT_P OUT_N buffer
.ends


* expanding   symbol:  cap_var.sym # of pins=4
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/cap_var.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/cap_var.sch
.subckt cap_var  OUT_P OUT_N GND Vtune
*.iopin OUT_P
*.iopin OUT_N
*.iopin Vtune
*.iopin GND
XC1 OUT_P Vtune GND sky130_fd_pr__cap_var_lvt W=4 L=0.6 VM=14 m=14
XC2 OUT_N Vtune GND sky130_fd_pr__cap_var_lvt W=4 L=0.6 VM=14 m=14
.ends


* expanding   symbol:  capbank.sym # of pins=10
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/capbank.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/capbank.sch
.subckt capbank  OUT_P OUT_N VDD GND bit0 bit1 bit2 bit3 bit4 bit5
*.iopin VDD
*.iopin GND
*.ipin bit0
*.ipin bit1
*.ipin bit2
*.ipin bit3
*.ipin bit4
*.ipin bit5
*.iopin OUT_P
*.iopin OUT_N
X1 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X2 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X3 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X4 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X5 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X6 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X7 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X8 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X9 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X10 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X11 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X12 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X13 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X14 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X15 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X16 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X17 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X18 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X19 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X20 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X21 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X22 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X23 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X24 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X25 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X26 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X27 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X28 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X29 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X30 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X31 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X32 w_inv5 bit5 OUT_P GND OUT_N cell_unit
X33 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X34 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X35 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X36 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X37 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X38 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X39 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X40 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X41 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X42 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X43 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X44 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X45 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X46 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X47 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X48 w_inv4 bit4 OUT_P GND OUT_N cell_unit
X49 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X50 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X51 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X52 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X53 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X54 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X55 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X56 w_inv3 bit3 OUT_P GND OUT_N cell_unit
X57 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X58 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X59 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X60 w_inv2 bit2 OUT_P GND OUT_N cell_unit
X61 w_inv1 bit1 OUT_P GND OUT_N cell_unit
X62 w_inv1 bit1 OUT_P GND OUT_N cell_unit
X63 w_inv0 bit0 OUT_P GND OUT_N cell_unit
X64 bit0 w_inv0 VDD GND inv
X65 bit1 w_inv1 VDD GND inv
X66 bit2 w_inv2 VDD GND inv
X67 bit3 w_inv3 VDD GND inv
X68 bit4 w_inv4 VDD GND inv
X69 bit5 w_inv5 VDD GND inv
.ends


* expanding   symbol:  vco_pmirr.sym # of pins=4
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_pmirr.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_pmirr.sch
.subckt vco_pmirr  VDD IND_CT GND VBIAS
*.iopin IND_CT
*.iopin VBIAS
*.iopin VDD
*.iopin GND
X25 VDD net1 net1 VDD rf_pfet_01v8_aM02W3p00L0p15
X17 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X18 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X19 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X20 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X21 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X22 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X23 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X24 VDD net1 IND_CT VDD rf_pfet_01v8_aM02W3p00L0p15
X1 VDD VDD VDD VDD rf_pfet_01v8_aM02W3p00L0p15
X2 VDD VDD VDD VDD rf_pfet_01v8_aM02W3p00L0p15
X3 VDD VDD VDD VDD rf_pfet_01v8_aM02W3p00L0p15
X4 VDD VDD VDD VDD rf_pfet_01v8_aM02W3p00L0p15
X5 VDD VDD VDD VDD rf_pfet_01v8_aM02W3p00L0p15
XR1 VBIAS net1 GND sky130_fd_pr__res_high_po_2p85 L=3.5 mult=1 m=1
.ends


* expanding   symbol:  vco_pair.sym # of pins=3
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_pair.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/vco_pair.sch
.subckt vco_pair  OUT_P OUT_N GND
*.iopin GND
*.iopin OUT_P
*.iopin OUT_N
X1 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X2 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X3 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X4 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X5 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X6 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X7 OUT_P OUT_N GND GND rf_nfet_01v8_aM02W5p00L0p15
X8 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X9 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X10 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X11 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X12 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X13 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X14 OUT_N OUT_P GND GND rf_nfet_01v8_aM02W5p00L0p15
X16 GND GND GND GND rf_nfet_01v8_aM02W5p00L0p15
X17 GND GND GND GND rf_nfet_01v8_aM02W5p00L0p15
X18 GND GND GND GND rf_nfet_01v8_aM02W5p00L0p15
X19 GND GND GND GND rf_nfet_01v8_aM02W5p00L0p15
.ends


* expanding   symbol:  buffer.sym # of pins=7
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/buffer.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/buffer.sch
.subckt buffer  VBIAS VDD GND OUT_N OUT_P IN_P IN_N
*.iopin VBIAS
*.iopin VDD
*.iopin GND
*.opin OUT_P
*.opin OUT_N
*.ipin IN_P
*.ipin IN_N
X10 OUT_N IN_P W_D GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X11 OUT_P IN_N W_D GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X12 OUT_N IN_P W_D GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X13 OUT_P IN_N W_D GND rf_nfet_01v8_lvt_aM04W5p00L0p15
R1 OUT_N VDD sky130_fd_pr__res_generic_po W=3.5 L=3.5 m=1
R2 OUT_P VDD sky130_fd_pr__res_generic_po W=3.5 L=3.5 m=1
X9 VBIAS VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X1 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X2 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X3 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X4 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X5 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X6 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X7 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X8 W_D VBIAS GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X14 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X15 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X16 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X17 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X18 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X19 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X20 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X21 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
X22 GND GND GND GND rf_nfet_01v8_lvt_aM04W5p00L0p15
.ends


* expanding   symbol:  cell_unit.sym # of pins=5
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/cell_unit.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/cell_unit.sch
.subckt cell_unit  V_bias ON OUT_N GND OUT_P
*.iopin OUT_N
*.iopin OUT_P
*.iopin GND
*.ipin ON
*.ipin V_bias
XC1 OUT_N net1 sky130_fd_pr__cap_mim_m3_1 W=3.3 L=3.3 MF=1 m=1
XC2 OUT_P net2 sky130_fd_pr__cap_mim_m3_1 W=3.3 L=3.3 MF=1 m=1
XR1 net1 V_bias GND sky130_fd_pr__res_xhigh_po_0p35 L=1.5 mult=1 m=1
XR2 net2 V_bias GND sky130_fd_pr__res_xhigh_po_0p35 L=1.5 mult=1 m=1
X1 net2 ON net1 GND rf_nfet_01v8_aM02W1p65L0p15
.ends


* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/inv.sym
** sch_path: /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/inv.sch
.subckt inv  IN OUT VDD GND
*.ipin IN
*.opin OUT
*.iopin VDD
*.iopin GND
XM1 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  rf_pfet_01v8_aM02W3p00L0p15.sym # of pins=4
** sym_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_pfet_01v8_aM02W3p00L0p15.sym
** sch_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_pfet_01v8_aM02W3p00L0p15.sch
.subckt rf_pfet_01v8_aM02W3p00L0p15  SOURCE GATE DRAIN BULK
*.iopin DRAIN
*.iopin SOURCE
*.ipin GATE
*.ipin BULK
**** begin user architecture code


X0 SOURCE GATE DRAIN BULK sky130_fd_pr__pfet_01v8 w=3.01e+06u l=150000u
X1 DRAIN GATE SOURCE BULK sky130_fd_pr__pfet_01v8 w=3.01e+06u l=150000u


**** end user architecture code
.ends


* expanding   symbol:  rf_nfet_01v8_aM02W5p00L0p15.sym # of pins=4
** sym_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_nfet_01v8_aM02W5p00L0p15.sym
** sch_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_nfet_01v8_aM02W5p00L0p15.sch
.subckt rf_nfet_01v8_aM02W5p00L0p15  DRAIN GATE SOURCE SUBSTRATE
*.iopin SOURCE
*.iopin DRAIN
*.ipin GATE
*.ipin SUBSTRATE
**** begin user architecture code


X0 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.05e+06u l=150000u
X1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 w=5.05e+06u l=150000u


**** end user architecture code
.ends


* expanding   symbol:  rf_nfet_01v8_lvt_aM04W5p00L0p15.sym # of pins=4
** sym_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_nfet_01v8_lvt_aM04W5p00L0p15.sym
** sch_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_nfet_01v8_lvt_aM04W5p00L0p15.sch
.subckt rf_nfet_01v8_lvt_aM04W5p00L0p15  DRAIN GATE SOURCE SUBSTRATE
*.iopin SOURCE
*.iopin DRAIN
*.ipin GATE
*.ipin SUBSTRATE
**** begin user architecture code


X0 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=150000u
X1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=150000u
X2 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=150000u
X3 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8_lvt w=5.05e+06u l=150000u


**** end user architecture code
.ends


* expanding   symbol:  rf_nfet_01v8_aM02W1p65L0p15.sym # of pins=4
** sym_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_nfet_01v8_aM02W1p65L0p15.sym
** sch_path:
*+ /home/shpeccy/ntfs_drive/Documents/Database/ESIC/caravel_asic_one/xschem/rf_nfet_01v8_aM02W1p65L0p15.sch
.subckt rf_nfet_01v8_aM02W1p65L0p15  DRAIN GATE SOURCE SUBSTRATE
*.iopin SOURCE
*.iopin DRAIN
*.ipin GATE
*.ipin SUBSTRATE
**** begin user architecture code


X0 SOURCE GATE DRAIN SUBSTRATE sky130_fd_pr__nfet_01v8 w=1.65e+06u l=150000u
X1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 w=1.65e+06u l=150000u


**** end user architecture code
.ends

.GLOBAL GND
.GLOBAL VDD
.end
