* NGSPICE file created from cell_unit_pex.ext - technology: sky130B

.subckt cell_unit_pex ON V_bias OUT_P OUT_N GND
X0 OUT_P.t0 a_n44_16.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X1 a_n44_16.t3 V_bias.t1 GND.t3 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X2 a_246_92.t1 V_bias.t0 GND.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X3 a_n44_16.t1 ON.t0 a_246_92.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X4 OUT_N.t0 a_246_92.t0 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X5 a_246_92.t2 ON.t1 a_n44_16.t0 GND.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
C0 OUT_P V_bias 2.36fF
C1 OUT_N ON 3.36fF
C2 OUT_N V_bias 2.36fF
C3 OUT_P ON 3.36fF
R0 OUT_P OUT_P.t0 0.21
R1 a_n44_16.n10 a_n44_16.t0 10.181
R2 a_n44_16.n10 a_n44_16.t1 10.181
R3 a_n44_16.t3 a_n44_16.n18 9.68
R4 a_n44_16.n1 a_n44_16.n0 9.302
R5 a_n44_16.n7 a_n44_16.n6 9.3
R6 a_n44_16.n5 a_n44_16.n4 9.3
R7 a_n44_16.n9 a_n44_16.n8 9
R8 a_n44_16.n13 a_n44_16.n12 7.729
R9 a_n44_16.n13 a_n44_16.n10 6.296
R10 a_n44_16.n16 a_n44_16.n1 4.508
R11 a_n44_16.n15 a_n44_16.n14 4.501
R12 a_n44_16.n15 a_n44_16.n9 4.501
R13 a_n44_16.n16 a_n44_16.n3 4.494
R14 a_n44_16.n18 a_n44_16.t2 1.259
R15 a_n44_16.n12 a_n44_16.n11 0.536
R16 a_n44_16.n18 a_n44_16.n17 0.415
R17 a_n44_16.n14 a_n44_16.n13 0.151
R18 a_n44_16.n7 a_n44_16.n5 0.028
R19 a_n44_16.n3 a_n44_16.n2 0.025
R20 a_n44_16.n17 a_n44_16.n16 0.021
R21 a_n44_16.n9 a_n44_16.n7 0.012
R22 a_n44_16.n16 a_n44_16.n15 0.006
R23 V_bias.n0 V_bias.t1 9.633
R24 V_bias.n0 V_bias.t0 9.587
R25 V_bias V_bias.n0 0.265
R26 GND.n5 GND.t0 650.171
R27 GND.n45 GND.t3 650.171
R28 GND.n5 GND.t1 582.13
R29 GND.n45 GND.t2 582.13
R30 GND.n69 GND.n68 55.353
R31 GND.n29 GND.n28 55.353
R32 GND.n61 GND.n60 54.344
R33 GND.n70 GND.n69 54.344
R34 GND.n21 GND.n20 54.344
R35 GND.n30 GND.n29 54.344
R36 GND.n51 GND.n50 47.551
R37 GND.n11 GND.n10 47.551
R38 GND.n43 GND.n42 22.848
R39 GND.n44 GND.n43 22.848
R40 GND.n3 GND.n2 22.848
R41 GND.n4 GND.n3 22.848
R42 GND.n46 GND.n44 10.189
R43 GND.n6 GND.n4 10.189
R44 GND.n52 GND.n51 9.861
R45 GND.n12 GND.n11 9.861
R46 GND.n53 GND.n52 9.457
R47 GND.n13 GND.n12 9.457
R48 GND.n76 GND.n75 9.3
R49 GND.n78 GND.n77 9.3
R50 GND.n57 GND.n56 9.3
R51 GND.n55 GND.n54 9.3
R52 GND.n65 GND.n64 9.3
R53 GND.n64 GND.n63 9.3
R54 GND.n74 GND.n73 9.3
R55 GND.n73 GND.n72 9.3
R56 GND.n47 GND.n46 9.3
R57 GND.n46 GND.n45 9.3
R58 GND.n36 GND.n35 9.3
R59 GND.n17 GND.n16 9.3
R60 GND.n15 GND.n14 9.3
R61 GND.n25 GND.n24 9.3
R62 GND.n24 GND.n23 9.3
R63 GND.n34 GND.n33 9.3
R64 GND.n33 GND.n32 9.3
R65 GND.n38 GND.n37 9.3
R66 GND.n7 GND.n6 9.3
R67 GND.n6 GND.n5 9.3
R68 GND.n59 GND.n58 6.023
R69 GND.n67 GND.n66 6.023
R70 GND.n19 GND.n18 6.023
R71 GND.n27 GND.n26 6.023
R72 GND.n49 GND.n48 5.27
R73 GND.n41 GND.n40 5.27
R74 GND.n9 GND.n8 5.27
R75 GND.n1 GND.n0 5.27
R76 GND.n55 GND.n53 4.048
R77 GND.n15 GND.n13 4.048
R78 GND.n79 GND.n47 3.924
R79 GND.n39 GND.n7 3.924
R80 GND.n71 GND.n70 3.324
R81 GND.n62 GND.n61 3.324
R82 GND.n31 GND.n30 3.324
R83 GND.n22 GND.n21 3.324
R84 GND.n53 GND.n49 1.129
R85 GND.n47 GND.n41 1.129
R86 GND.n13 GND.n9 1.129
R87 GND.n7 GND.n1 1.129
R88 GND GND.n80 1.091
R89 GND.n80 GND.n79 0.919
R90 GND.n80 GND.n39 0.919
R91 GND.n64 GND.n59 0.376
R92 GND.n73 GND.n67 0.376
R93 GND.n24 GND.n19 0.376
R94 GND.n33 GND.n27 0.376
R95 GND.n74 GND.n65 0.15
R96 GND.n34 GND.n25 0.15
R97 GND.n79 GND.n78 0.125
R98 GND.n39 GND.n38 0.125
R99 GND.n63 GND.n62 0.053
R100 GND.n72 GND.n71 0.053
R101 GND.n23 GND.n22 0.053
R102 GND.n32 GND.n31 0.053
R103 GND.n57 GND.n55 0.034
R104 GND.n78 GND.n76 0.034
R105 GND.n17 GND.n15 0.034
R106 GND.n38 GND.n36 0.034
R107 GND.n65 GND.n57 0.002
R108 GND.n76 GND.n74 0.002
R109 GND.n25 GND.n17 0.002
R110 GND.n36 GND.n34 0.002
R111 a_246_92.n26 a_246_92.t2 10.181
R112 a_246_92.n18 a_246_92.t3 10.181
R113 a_246_92.t1 a_246_92.n39 9.68
R114 a_246_92.n3 a_246_92.n2 9.302
R115 a_246_92.n13 a_246_92.n12 9.302
R116 a_246_92.n32 a_246_92.n31 9.3
R117 a_246_92.n34 a_246_92.n33 9.3
R118 a_246_92.n7 a_246_92.n6 9.3
R119 a_246_92.n5 a_246_92.n4 9.3
R120 a_246_92.n36 a_246_92.n35 9
R121 a_246_92.n9 a_246_92.n8 9
R122 a_246_92.n27 a_246_92.n25 7.729
R123 a_246_92.n19 a_246_92.n17 7.729
R124 a_246_92.n27 a_246_92.n26 6.296
R125 a_246_92.n19 a_246_92.n18 6.296
R126 a_246_92.n30 a_246_92.n3 4.508
R127 a_246_92.n14 a_246_92.n13 4.508
R128 a_246_92.n37 a_246_92.n36 4.496
R129 a_246_92.n21 a_246_92.n20 4.496
R130 a_246_92.n29 a_246_92.n28 4.495
R131 a_246_92.n10 a_246_92.n9 4.495
R132 a_246_92.n14 a_246_92.n11 4.494
R133 a_246_92.n30 a_246_92.n1 4.494
R134 a_246_92.n39 a_246_92.t0 1.087
R135 a_246_92.n25 a_246_92.n24 0.536
R136 a_246_92.n17 a_246_92.n16 0.536
R137 a_246_92.n39 a_246_92.n38 0.255
R138 a_246_92.n28 a_246_92.n27 0.151
R139 a_246_92.n20 a_246_92.n19 0.151
R140 a_246_92.n23 a_246_92.n22 0.125
R141 a_246_92.n34 a_246_92.n32 0.028
R142 a_246_92.n7 a_246_92.n5 0.028
R143 a_246_92.n1 a_246_92.n0 0.025
R144 a_246_92.n20 a_246_92.n15 0.024
R145 a_246_92.n36 a_246_92.n34 0.012
R146 a_246_92.n9 a_246_92.n7 0.012
R147 a_246_92.n29 a_246_92.n23 0.011
R148 a_246_92.n30 a_246_92.n29 0.011
R149 a_246_92.n14 a_246_92.n10 0.011
R150 a_246_92.n38 a_246_92.n37 0.01
R151 a_246_92.n22 a_246_92.n21 0.01
R152 a_246_92.n21 a_246_92.n14 0.01
R153 a_246_92.n37 a_246_92.n30 0.01
R154 ON.n4 ON.t1 300.446
R155 ON.n2 ON.t0 300.446
R156 ON.n3 ON.n2 27.537
R157 ON.n5 ON.n4 24.127
R158 ON.n1 ON.n0 8.764
R159 ON.n6 ON.n5 4.661
R160 ON.n3 ON.n1 3.401
R161 ON.n6 ON.n3 0.626
R162 ON ON.n6 0.586
R163 OUT_N OUT_N.t0 0.211
C4 OUT_N GND 14.65fF
C5 OUT_P GND 13.53fF
C6 ON GND 25.76fF
C7 V_bias GND 22.38fF
C8 OUT_N.t0 GND 2.95fF $ **FLOATING
C9 ON.n0 GND 0.00fF
C10 ON.n1 GND 0.00fF
C11 ON.t0 GND 0.03fF $ **FLOATING
C12 ON.n2 GND 0.01fF
C13 ON.n3 GND 0.00fF
C14 ON.t1 GND 0.03fF $ **FLOATING
C15 ON.n4 GND 0.01fF
C16 ON.n5 GND 0.00fF
C17 ON.n6 GND 7.37fF
C18 a_246_92.n0 GND 0.00fF
C19 a_246_92.n1 GND 0.00fF
C20 a_246_92.n2 GND 0.01fF
C21 a_246_92.n3 GND 0.01fF
C22 a_246_92.n4 GND 0.00fF
C23 a_246_92.n5 GND 0.00fF
C24 a_246_92.n6 GND 0.00fF
C25 a_246_92.n7 GND 0.00fF
C26 a_246_92.n8 GND 0.00fF
C27 a_246_92.n9 GND 0.00fF
C28 a_246_92.n10 GND 0.09fF
C29 a_246_92.n11 GND 0.00fF
C30 a_246_92.n12 GND 0.01fF
C31 a_246_92.n13 GND 0.01fF
C32 a_246_92.n14 GND 0.01fF
C33 a_246_92.n15 GND 0.00fF
C34 a_246_92.n16 GND 0.00fF
C35 a_246_92.n17 GND 0.00fF
C36 a_246_92.t3 GND 0.02fF $ **FLOATING
C37 a_246_92.n18 GND 0.07fF
C38 a_246_92.n19 GND 0.02fF
C39 a_246_92.n20 GND 0.05fF
C40 a_246_92.n22 GND 0.04fF
C41 a_246_92.n23 GND 0.04fF
C42 a_246_92.n24 GND 0.00fF
C43 a_246_92.n25 GND 0.00fF
C44 a_246_92.t2 GND 0.02fF $ **FLOATING
C45 a_246_92.n26 GND 0.07fF
C46 a_246_92.n27 GND 0.02fF
C47 a_246_92.n28 GND 0.05fF
C48 a_246_92.n30 GND 0.01fF
C49 a_246_92.n31 GND 0.00fF
C50 a_246_92.n32 GND 0.00fF
C51 a_246_92.n33 GND 0.00fF
C52 a_246_92.n34 GND 0.00fF
C53 a_246_92.n35 GND 0.00fF
C54 a_246_92.n36 GND 0.00fF
C55 a_246_92.n38 GND 0.08fF
C56 a_246_92.t0 GND 4.19fF $ **FLOATING
C57 a_246_92.n39 GND 0.61fF
C58 a_246_92.t1 GND 0.26fF $ **FLOATING
C59 V_bias.t0 GND 0.07fF $ **FLOATING
C60 V_bias.t1 GND 0.12fF $ **FLOATING
C61 V_bias.n0 GND 16.80fF
C62 a_n44_16.n0 GND 0.01fF
C63 a_n44_16.n1 GND 0.01fF
C64 a_n44_16.n2 GND 0.00fF
C65 a_n44_16.n3 GND 0.00fF
C66 a_n44_16.n4 GND 0.00fF
C67 a_n44_16.n5 GND 0.00fF
C68 a_n44_16.n6 GND 0.00fF
C69 a_n44_16.n7 GND 0.00fF
C70 a_n44_16.n8 GND 0.00fF
C71 a_n44_16.n9 GND 0.00fF
C72 a_n44_16.t0 GND 0.02fF $ **FLOATING
C73 a_n44_16.t1 GND 0.02fF $ **FLOATING
C74 a_n44_16.n10 GND 0.05fF
C75 a_n44_16.n11 GND 0.00fF
C76 a_n44_16.n12 GND 0.00fF
C77 a_n44_16.n13 GND 0.02fF
C78 a_n44_16.n14 GND 0.04fF
C79 a_n44_16.n15 GND 0.12fF
C80 a_n44_16.n16 GND 0.01fF
C81 a_n44_16.n17 GND 0.12fF
C82 a_n44_16.t2 GND 3.87fF $ **FLOATING
C83 a_n44_16.n18 GND 0.52fF
C84 a_n44_16.t3 GND 0.24fF $ **FLOATING
C85 OUT_P.t0 GND 4.04fF $ **FLOATING
.ends
