magic
tech sky130B
magscale 1 2
timestamp 1654467620
<< psubdiff >>
rect 26 2720 4874 2732
rect 26 2686 72 2720
rect 106 2686 146 2720
rect 180 2686 220 2720
rect 254 2686 294 2720
rect 328 2686 368 2720
rect 402 2686 442 2720
rect 476 2686 516 2720
rect 550 2686 590 2720
rect 624 2686 664 2720
rect 698 2686 738 2720
rect 772 2686 812 2720
rect 846 2686 886 2720
rect 920 2686 960 2720
rect 994 2686 1034 2720
rect 1068 2686 1108 2720
rect 1142 2686 1182 2720
rect 1216 2686 1256 2720
rect 1290 2686 1330 2720
rect 1364 2686 1404 2720
rect 1438 2686 1478 2720
rect 1512 2686 1552 2720
rect 1586 2686 1626 2720
rect 1660 2686 1700 2720
rect 1734 2686 1774 2720
rect 1808 2686 1848 2720
rect 1882 2686 1922 2720
rect 1956 2686 1996 2720
rect 2030 2686 2070 2720
rect 2104 2686 2144 2720
rect 2178 2686 2218 2720
rect 2252 2686 2292 2720
rect 2326 2686 2366 2720
rect 2400 2686 2440 2720
rect 2474 2686 2514 2720
rect 2548 2686 2588 2720
rect 2622 2686 2662 2720
rect 2696 2686 2736 2720
rect 2770 2686 2810 2720
rect 2844 2686 2884 2720
rect 2918 2686 2958 2720
rect 2992 2686 3032 2720
rect 3066 2686 3106 2720
rect 3140 2686 3180 2720
rect 3214 2686 3254 2720
rect 3288 2686 3328 2720
rect 3362 2686 3402 2720
rect 3436 2686 3476 2720
rect 3510 2686 3550 2720
rect 3584 2686 3624 2720
rect 3658 2686 3698 2720
rect 3732 2686 3772 2720
rect 3806 2686 3846 2720
rect 3880 2686 3920 2720
rect 3954 2686 3994 2720
rect 4028 2686 4068 2720
rect 4102 2686 4142 2720
rect 4176 2686 4216 2720
rect 4250 2686 4290 2720
rect 4324 2686 4364 2720
rect 4398 2686 4438 2720
rect 4472 2686 4512 2720
rect 4546 2686 4586 2720
rect 4620 2686 4660 2720
rect 4694 2686 4734 2720
rect 4768 2686 4808 2720
rect 4842 2686 4874 2720
rect 26 2666 4874 2686
rect 26 92 84 2666
rect 592 92 650 2666
rect 730 92 788 2666
rect 1296 92 1354 2666
rect 1434 92 1492 2666
rect 2000 92 2058 2666
rect 2138 92 2196 2666
rect 2704 92 2762 2666
rect 2842 92 2900 2666
rect 3408 92 3466 2666
rect 3546 92 3604 2666
rect 4112 92 4170 2666
rect 4250 92 4308 2666
rect 4816 2546 4874 2666
rect 4816 92 4874 218
rect 26 72 4874 92
rect 26 38 72 72
rect 106 38 146 72
rect 180 38 220 72
rect 254 38 294 72
rect 328 38 368 72
rect 402 38 442 72
rect 476 38 516 72
rect 550 38 590 72
rect 624 38 664 72
rect 698 38 738 72
rect 772 38 812 72
rect 846 38 886 72
rect 920 38 960 72
rect 994 38 1034 72
rect 1068 38 1108 72
rect 1142 38 1182 72
rect 1216 38 1256 72
rect 1290 38 1330 72
rect 1364 38 1404 72
rect 1438 38 1478 72
rect 1512 38 1552 72
rect 1586 38 1626 72
rect 1660 38 1700 72
rect 1734 38 1774 72
rect 1808 38 1848 72
rect 1882 38 1922 72
rect 1956 38 1996 72
rect 2030 38 2070 72
rect 2104 38 2144 72
rect 2178 38 2218 72
rect 2252 38 2292 72
rect 2326 38 2366 72
rect 2400 38 2440 72
rect 2474 38 2514 72
rect 2548 38 2588 72
rect 2622 38 2662 72
rect 2696 38 2736 72
rect 2770 38 2810 72
rect 2844 38 2884 72
rect 2918 38 2958 72
rect 2992 38 3032 72
rect 3066 38 3106 72
rect 3140 38 3180 72
rect 3214 38 3254 72
rect 3288 38 3328 72
rect 3362 38 3402 72
rect 3436 38 3476 72
rect 3510 38 3550 72
rect 3584 38 3624 72
rect 3658 38 3698 72
rect 3732 38 3772 72
rect 3806 38 3846 72
rect 3880 38 3920 72
rect 3954 38 3994 72
rect 4028 38 4068 72
rect 4102 38 4142 72
rect 4176 38 4216 72
rect 4250 38 4290 72
rect 4324 38 4364 72
rect 4398 38 4438 72
rect 4472 38 4512 72
rect 4546 38 4586 72
rect 4620 38 4660 72
rect 4694 38 4734 72
rect 4768 38 4808 72
rect 4842 38 4874 72
rect 26 26 4874 38
<< psubdiffcont >>
rect 72 2686 106 2720
rect 146 2686 180 2720
rect 220 2686 254 2720
rect 294 2686 328 2720
rect 368 2686 402 2720
rect 442 2686 476 2720
rect 516 2686 550 2720
rect 590 2686 624 2720
rect 664 2686 698 2720
rect 738 2686 772 2720
rect 812 2686 846 2720
rect 886 2686 920 2720
rect 960 2686 994 2720
rect 1034 2686 1068 2720
rect 1108 2686 1142 2720
rect 1182 2686 1216 2720
rect 1256 2686 1290 2720
rect 1330 2686 1364 2720
rect 1404 2686 1438 2720
rect 1478 2686 1512 2720
rect 1552 2686 1586 2720
rect 1626 2686 1660 2720
rect 1700 2686 1734 2720
rect 1774 2686 1808 2720
rect 1848 2686 1882 2720
rect 1922 2686 1956 2720
rect 1996 2686 2030 2720
rect 2070 2686 2104 2720
rect 2144 2686 2178 2720
rect 2218 2686 2252 2720
rect 2292 2686 2326 2720
rect 2366 2686 2400 2720
rect 2440 2686 2474 2720
rect 2514 2686 2548 2720
rect 2588 2686 2622 2720
rect 2662 2686 2696 2720
rect 2736 2686 2770 2720
rect 2810 2686 2844 2720
rect 2884 2686 2918 2720
rect 2958 2686 2992 2720
rect 3032 2686 3066 2720
rect 3106 2686 3140 2720
rect 3180 2686 3214 2720
rect 3254 2686 3288 2720
rect 3328 2686 3362 2720
rect 3402 2686 3436 2720
rect 3476 2686 3510 2720
rect 3550 2686 3584 2720
rect 3624 2686 3658 2720
rect 3698 2686 3732 2720
rect 3772 2686 3806 2720
rect 3846 2686 3880 2720
rect 3920 2686 3954 2720
rect 3994 2686 4028 2720
rect 4068 2686 4102 2720
rect 4142 2686 4176 2720
rect 4216 2686 4250 2720
rect 4290 2686 4324 2720
rect 4364 2686 4398 2720
rect 4438 2686 4472 2720
rect 4512 2686 4546 2720
rect 4586 2686 4620 2720
rect 4660 2686 4694 2720
rect 4734 2686 4768 2720
rect 4808 2686 4842 2720
rect 72 38 106 72
rect 146 38 180 72
rect 220 38 254 72
rect 294 38 328 72
rect 368 38 402 72
rect 442 38 476 72
rect 516 38 550 72
rect 590 38 624 72
rect 664 38 698 72
rect 738 38 772 72
rect 812 38 846 72
rect 886 38 920 72
rect 960 38 994 72
rect 1034 38 1068 72
rect 1108 38 1142 72
rect 1182 38 1216 72
rect 1256 38 1290 72
rect 1330 38 1364 72
rect 1404 38 1438 72
rect 1478 38 1512 72
rect 1552 38 1586 72
rect 1626 38 1660 72
rect 1700 38 1734 72
rect 1774 38 1808 72
rect 1848 38 1882 72
rect 1922 38 1956 72
rect 1996 38 2030 72
rect 2070 38 2104 72
rect 2144 38 2178 72
rect 2218 38 2252 72
rect 2292 38 2326 72
rect 2366 38 2400 72
rect 2440 38 2474 72
rect 2514 38 2548 72
rect 2588 38 2622 72
rect 2662 38 2696 72
rect 2736 38 2770 72
rect 2810 38 2844 72
rect 2884 38 2918 72
rect 2958 38 2992 72
rect 3032 38 3066 72
rect 3106 38 3140 72
rect 3180 38 3214 72
rect 3254 38 3288 72
rect 3328 38 3362 72
rect 3402 38 3436 72
rect 3476 38 3510 72
rect 3550 38 3584 72
rect 3624 38 3658 72
rect 3698 38 3732 72
rect 3772 38 3806 72
rect 3846 38 3880 72
rect 3920 38 3954 72
rect 3994 38 4028 72
rect 4068 38 4102 72
rect 4142 38 4176 72
rect 4216 38 4250 72
rect 4290 38 4324 72
rect 4364 38 4398 72
rect 4438 38 4472 72
rect 4512 38 4546 72
rect 4586 38 4620 72
rect 4660 38 4694 72
rect 4734 38 4768 72
rect 4808 38 4842 72
<< locali >>
rect 38 2526 72 2720
rect 106 2686 146 2720
rect 180 2686 220 2720
rect 254 2686 294 2720
rect 328 2686 368 2720
rect 402 2686 442 2720
rect 476 2686 516 2720
rect 550 2686 590 2720
rect 624 2686 664 2720
rect 698 2686 738 2720
rect 772 2686 812 2720
rect 846 2686 886 2720
rect 920 2686 960 2720
rect 994 2686 1034 2720
rect 1068 2686 1108 2720
rect 1142 2686 1182 2720
rect 1216 2686 1256 2720
rect 1290 2686 1330 2720
rect 1364 2686 1404 2720
rect 1438 2686 1478 2720
rect 1512 2686 1552 2720
rect 1586 2686 1626 2720
rect 1660 2686 1700 2720
rect 1734 2686 1774 2720
rect 1808 2686 1848 2720
rect 1882 2686 1922 2720
rect 1956 2686 1996 2720
rect 2030 2686 2070 2720
rect 2104 2686 2144 2720
rect 2178 2686 2218 2720
rect 2252 2686 2292 2720
rect 2326 2686 2366 2720
rect 2400 2686 2440 2720
rect 2474 2686 2514 2720
rect 2548 2686 2588 2720
rect 2622 2686 2662 2720
rect 2696 2686 2736 2720
rect 2770 2686 2810 2720
rect 2844 2686 2884 2720
rect 2918 2686 2958 2720
rect 2992 2686 3032 2720
rect 3066 2686 3106 2720
rect 3140 2686 3180 2720
rect 3214 2686 3254 2720
rect 3288 2686 3328 2720
rect 3362 2686 3402 2720
rect 3436 2686 3476 2720
rect 3510 2686 3550 2720
rect 3584 2686 3624 2720
rect 3658 2686 3698 2720
rect 3732 2686 3772 2720
rect 3806 2686 3846 2720
rect 3880 2686 3920 2720
rect 3954 2686 3994 2720
rect 4028 2686 4068 2720
rect 4102 2686 4142 2720
rect 4176 2686 4216 2720
rect 4250 2686 4290 2720
rect 4324 2686 4364 2720
rect 4398 2686 4438 2720
rect 4472 2686 4512 2720
rect 4546 2686 4586 2720
rect 4620 2686 4660 2720
rect 4694 2686 4734 2720
rect 4768 2686 4808 2720
rect 4842 2686 4862 2720
rect 38 38 72 232
rect 604 72 638 2686
rect 742 72 776 2686
rect 1308 72 1342 2686
rect 1446 72 1480 2686
rect 2012 72 2046 2686
rect 2150 72 2184 2686
rect 2716 72 2750 2686
rect 2854 72 2888 2686
rect 3420 72 3454 2686
rect 3558 72 3592 2686
rect 4124 72 4158 2686
rect 4262 72 4296 2686
rect 4828 72 4862 2686
rect 106 38 146 72
rect 180 38 220 72
rect 254 38 294 72
rect 328 38 368 72
rect 402 38 442 72
rect 476 38 516 72
rect 550 38 590 72
rect 624 38 664 72
rect 698 38 738 72
rect 772 38 812 72
rect 846 38 886 72
rect 920 38 960 72
rect 994 38 1034 72
rect 1068 38 1108 72
rect 1142 38 1182 72
rect 1216 38 1256 72
rect 1290 38 1330 72
rect 1364 38 1404 72
rect 1438 38 1478 72
rect 1512 38 1552 72
rect 1586 38 1626 72
rect 1660 38 1700 72
rect 1734 38 1774 72
rect 1808 38 1848 72
rect 1882 38 1922 72
rect 1956 38 1996 72
rect 2030 38 2070 72
rect 2104 38 2144 72
rect 2178 38 2218 72
rect 2252 38 2292 72
rect 2326 38 2366 72
rect 2400 38 2440 72
rect 2474 38 2514 72
rect 2548 38 2588 72
rect 2622 38 2662 72
rect 2696 38 2736 72
rect 2770 38 2810 72
rect 2844 38 2884 72
rect 2918 38 2958 72
rect 2992 38 3032 72
rect 3066 38 3106 72
rect 3140 38 3180 72
rect 3214 38 3254 72
rect 3288 38 3328 72
rect 3362 38 3402 72
rect 3436 38 3476 72
rect 3510 38 3550 72
rect 3584 38 3624 72
rect 3658 38 3698 72
rect 3732 38 3772 72
rect 3806 38 3846 72
rect 3880 38 3920 72
rect 3954 38 3994 72
rect 4028 38 4068 72
rect 4102 38 4142 72
rect 4176 38 4216 72
rect 4250 38 4290 72
rect 4324 38 4364 72
rect 4398 38 4438 72
rect 4472 38 4512 72
rect 4546 38 4586 72
rect 4620 38 4660 72
rect 4694 38 4734 72
rect 4768 38 4808 72
rect 4842 38 4862 72
<< viali >>
rect 72 2686 106 2720
rect 146 2686 180 2720
rect 220 2686 254 2720
rect 294 2686 328 2720
rect 368 2686 402 2720
rect 442 2686 476 2720
rect 516 2686 550 2720
rect 590 2686 624 2720
rect 664 2686 698 2720
rect 738 2686 772 2720
rect 812 2686 846 2720
rect 886 2686 920 2720
rect 960 2686 994 2720
rect 1034 2686 1068 2720
rect 1108 2686 1142 2720
rect 1182 2686 1216 2720
rect 1256 2686 1290 2720
rect 1330 2686 1364 2720
rect 1404 2686 1438 2720
rect 1478 2686 1512 2720
rect 1552 2686 1586 2720
rect 1626 2686 1660 2720
rect 1700 2686 1734 2720
rect 1774 2686 1808 2720
rect 1848 2686 1882 2720
rect 1922 2686 1956 2720
rect 1996 2686 2030 2720
rect 2070 2686 2104 2720
rect 2144 2686 2178 2720
rect 2218 2686 2252 2720
rect 2292 2686 2326 2720
rect 2366 2686 2400 2720
rect 2440 2686 2474 2720
rect 2514 2686 2548 2720
rect 2588 2686 2622 2720
rect 2662 2686 2696 2720
rect 2736 2686 2770 2720
rect 2810 2686 2844 2720
rect 2884 2686 2918 2720
rect 2958 2686 2992 2720
rect 3032 2686 3066 2720
rect 3106 2686 3140 2720
rect 3180 2686 3214 2720
rect 3254 2686 3288 2720
rect 3328 2686 3362 2720
rect 3402 2686 3436 2720
rect 3476 2686 3510 2720
rect 3550 2686 3584 2720
rect 3624 2686 3658 2720
rect 3698 2686 3732 2720
rect 3772 2686 3806 2720
rect 3846 2686 3880 2720
rect 3920 2686 3954 2720
rect 3994 2686 4028 2720
rect 4068 2686 4102 2720
rect 4142 2686 4176 2720
rect 4216 2686 4250 2720
rect 4290 2686 4324 2720
rect 4364 2686 4398 2720
rect 4438 2686 4472 2720
rect 4512 2686 4546 2720
rect 4586 2686 4620 2720
rect 4660 2686 4694 2720
rect 4734 2686 4768 2720
rect 4808 2686 4842 2720
rect 72 38 106 72
rect 146 38 180 72
rect 220 38 254 72
rect 294 38 328 72
rect 368 38 402 72
rect 442 38 476 72
rect 516 38 550 72
rect 590 38 624 72
rect 664 38 698 72
rect 738 38 772 72
rect 812 38 846 72
rect 886 38 920 72
rect 960 38 994 72
rect 1034 38 1068 72
rect 1108 38 1142 72
rect 1182 38 1216 72
rect 1256 38 1290 72
rect 1330 38 1364 72
rect 1404 38 1438 72
rect 1478 38 1512 72
rect 1552 38 1586 72
rect 1626 38 1660 72
rect 1700 38 1734 72
rect 1774 38 1808 72
rect 1848 38 1882 72
rect 1922 38 1956 72
rect 1996 38 2030 72
rect 2070 38 2104 72
rect 2144 38 2178 72
rect 2218 38 2252 72
rect 2292 38 2326 72
rect 2366 38 2400 72
rect 2440 38 2474 72
rect 2514 38 2548 72
rect 2588 38 2622 72
rect 2662 38 2696 72
rect 2736 38 2770 72
rect 2810 38 2844 72
rect 2884 38 2918 72
rect 2958 38 2992 72
rect 3032 38 3066 72
rect 3106 38 3140 72
rect 3180 38 3214 72
rect 3254 38 3288 72
rect 3328 38 3362 72
rect 3402 38 3436 72
rect 3476 38 3510 72
rect 3550 38 3584 72
rect 3624 38 3658 72
rect 3698 38 3732 72
rect 3772 38 3806 72
rect 3846 38 3880 72
rect 3920 38 3954 72
rect 3994 38 4028 72
rect 4068 38 4102 72
rect 4142 38 4176 72
rect 4216 38 4250 72
rect 4290 38 4324 72
rect 4364 38 4398 72
rect 4438 38 4472 72
rect 4512 38 4546 72
rect 4586 38 4620 72
rect 4660 38 4694 72
rect 4734 38 4768 72
rect 4808 38 4842 72
<< metal1 >>
rect 26 2720 4874 2732
rect 26 2686 72 2720
rect 106 2686 146 2720
rect 180 2686 220 2720
rect 254 2686 294 2720
rect 328 2686 368 2720
rect 402 2686 442 2720
rect 476 2686 516 2720
rect 550 2686 590 2720
rect 624 2686 664 2720
rect 698 2686 738 2720
rect 772 2686 812 2720
rect 846 2686 886 2720
rect 920 2686 960 2720
rect 994 2686 1034 2720
rect 1068 2686 1108 2720
rect 1142 2686 1182 2720
rect 1216 2686 1256 2720
rect 1290 2686 1330 2720
rect 1364 2686 1404 2720
rect 1438 2686 1478 2720
rect 1512 2686 1552 2720
rect 1586 2686 1626 2720
rect 1660 2686 1700 2720
rect 1734 2686 1774 2720
rect 1808 2686 1848 2720
rect 1882 2686 1922 2720
rect 1956 2686 1996 2720
rect 2030 2686 2070 2720
rect 2104 2686 2144 2720
rect 2178 2686 2218 2720
rect 2252 2686 2292 2720
rect 2326 2686 2366 2720
rect 2400 2686 2440 2720
rect 2474 2686 2514 2720
rect 2548 2686 2588 2720
rect 2622 2686 2662 2720
rect 2696 2686 2736 2720
rect 2770 2686 2810 2720
rect 2844 2686 2884 2720
rect 2918 2686 2958 2720
rect 2992 2686 3032 2720
rect 3066 2686 3106 2720
rect 3140 2686 3180 2720
rect 3214 2686 3254 2720
rect 3288 2686 3328 2720
rect 3362 2686 3402 2720
rect 3436 2686 3476 2720
rect 3510 2686 3550 2720
rect 3584 2686 3624 2720
rect 3658 2686 3698 2720
rect 3732 2686 3772 2720
rect 3806 2686 3846 2720
rect 3880 2686 3920 2720
rect 3954 2686 3994 2720
rect 4028 2686 4068 2720
rect 4102 2686 4142 2720
rect 4176 2686 4216 2720
rect 4250 2686 4290 2720
rect 4324 2686 4364 2720
rect 4398 2686 4438 2720
rect 4472 2686 4512 2720
rect 4546 2686 4586 2720
rect 4620 2686 4660 2720
rect 4694 2686 4734 2720
rect 4768 2686 4808 2720
rect 4842 2686 4874 2720
rect 26 2666 4874 2686
rect 26 2572 650 2666
rect 26 2520 84 2572
rect 140 2538 192 2572
rect 226 2538 278 2572
rect 312 2538 364 2572
rect 398 2538 450 2572
rect 484 2538 536 2572
rect 592 2534 650 2572
rect 730 2520 788 2666
rect 866 2632 1214 2638
rect 866 2580 888 2632
rect 940 2580 974 2632
rect 1026 2580 1052 2632
rect 1104 2580 1134 2632
rect 1186 2580 1214 2632
rect 866 2572 1214 2580
rect 1296 2534 1354 2666
rect 1434 2520 1492 2666
rect 1570 2632 1918 2638
rect 1570 2580 1592 2632
rect 1644 2580 1678 2632
rect 1730 2580 1756 2632
rect 1808 2580 1838 2632
rect 1890 2580 1918 2632
rect 1570 2572 1918 2580
rect 2000 2534 2058 2666
rect 2138 2520 2196 2666
rect 2276 2632 2624 2638
rect 2276 2580 2298 2632
rect 2350 2580 2384 2632
rect 2436 2580 2462 2632
rect 2514 2580 2544 2632
rect 2596 2580 2624 2632
rect 2276 2572 2624 2580
rect 2704 2534 2762 2666
rect 2842 2520 2900 2666
rect 2980 2632 3328 2638
rect 2980 2580 3002 2632
rect 3054 2580 3088 2632
rect 3140 2580 3166 2632
rect 3218 2580 3248 2632
rect 3300 2580 3328 2632
rect 2980 2572 3328 2580
rect 3408 2534 3466 2666
rect 3546 2520 3604 2666
rect 3684 2632 4032 2638
rect 3684 2580 3706 2632
rect 3758 2580 3792 2632
rect 3844 2580 3870 2632
rect 3922 2580 3952 2632
rect 4004 2580 4032 2632
rect 3684 2572 4032 2580
rect 4112 2534 4170 2666
rect 4250 2572 4874 2666
rect 4250 2538 4308 2572
rect 4364 2538 4416 2572
rect 4450 2538 4502 2572
rect 4536 2538 4588 2572
rect 4622 2538 4674 2572
rect 4708 2538 4760 2572
rect 4816 2538 4874 2572
rect 26 1510 84 1544
rect 140 1510 192 1544
rect 226 1510 278 1544
rect 312 1510 364 1544
rect 398 1510 450 1544
rect 484 1510 536 1544
rect 592 1510 650 1546
rect 26 1444 650 1510
rect 592 1314 650 1444
rect 26 1248 650 1314
rect 26 1214 84 1248
rect 140 1214 192 1248
rect 226 1214 278 1248
rect 312 1214 364 1248
rect 398 1214 450 1248
rect 484 1214 536 1248
rect 592 1212 650 1248
rect 730 1210 788 1544
rect 868 1490 1216 1508
rect 868 1438 890 1490
rect 942 1438 976 1490
rect 1028 1438 1054 1490
rect 1106 1438 1136 1490
rect 1188 1438 1216 1490
rect 868 1414 1216 1438
rect 868 1324 1216 1342
rect 868 1272 890 1324
rect 942 1272 976 1324
rect 1028 1272 1054 1324
rect 1106 1272 1136 1324
rect 1188 1272 1216 1324
rect 868 1248 1216 1272
rect 1296 1212 1354 1546
rect 1434 1210 1492 1544
rect 1572 1490 1920 1508
rect 1572 1438 1594 1490
rect 1646 1438 1680 1490
rect 1732 1438 1758 1490
rect 1810 1438 1840 1490
rect 1892 1438 1920 1490
rect 1572 1414 1920 1438
rect 1572 1324 1920 1342
rect 1572 1272 1594 1324
rect 1646 1272 1680 1324
rect 1732 1272 1758 1324
rect 1810 1272 1840 1324
rect 1892 1272 1920 1324
rect 1572 1248 1920 1272
rect 2000 1212 2058 1546
rect 2138 1314 2196 1544
rect 2276 1490 2624 1508
rect 2276 1438 2298 1490
rect 2350 1438 2384 1490
rect 2436 1438 2462 1490
rect 2514 1438 2544 1490
rect 2596 1438 2624 1490
rect 2276 1414 2624 1438
rect 2704 1314 2762 1546
rect 2138 1248 2762 1314
rect 2138 1210 2196 1248
rect 2252 1214 2304 1248
rect 2338 1214 2390 1248
rect 2424 1214 2476 1248
rect 2510 1214 2562 1248
rect 2596 1214 2648 1248
rect 2704 1212 2762 1248
rect 2842 1210 2900 1544
rect 2980 1490 3328 1508
rect 2980 1438 3002 1490
rect 3054 1438 3088 1490
rect 3140 1438 3166 1490
rect 3218 1438 3248 1490
rect 3300 1438 3328 1490
rect 2980 1414 3328 1438
rect 2980 1324 3328 1342
rect 2980 1272 3002 1324
rect 3054 1272 3088 1324
rect 3140 1272 3166 1324
rect 3218 1272 3248 1324
rect 3300 1272 3328 1324
rect 2980 1248 3328 1272
rect 3408 1212 3466 1546
rect 3546 1210 3604 1544
rect 3684 1490 4032 1508
rect 3684 1438 3706 1490
rect 3758 1438 3792 1490
rect 3844 1438 3870 1490
rect 3922 1438 3952 1490
rect 4004 1438 4032 1490
rect 3684 1414 4032 1438
rect 3684 1324 4032 1342
rect 3684 1272 3706 1324
rect 3758 1272 3792 1324
rect 3844 1272 3870 1324
rect 3922 1272 3952 1324
rect 4004 1272 4032 1324
rect 3684 1248 4032 1272
rect 4112 1212 4170 1544
rect 4250 1510 4308 1544
rect 4364 1510 4416 1544
rect 4450 1510 4502 1544
rect 4536 1510 4588 1544
rect 4622 1510 4674 1544
rect 4708 1510 4760 1544
rect 4816 1510 4874 1560
rect 4250 1444 4874 1510
rect 4250 1314 4308 1444
rect 4816 1314 4874 1444
rect 4250 1248 4874 1314
rect 4250 1210 4308 1248
rect 4364 1214 4416 1248
rect 4450 1214 4502 1248
rect 4536 1214 4588 1248
rect 4622 1214 4674 1248
rect 4708 1214 4760 1248
rect 4816 1214 4874 1248
rect 26 186 84 222
rect 140 186 192 220
rect 226 186 278 220
rect 312 186 364 220
rect 398 186 450 220
rect 484 186 536 220
rect 592 186 650 250
rect 26 140 180 186
rect 510 140 650 186
rect 26 92 650 140
rect 730 92 788 246
rect 868 180 1216 186
rect 868 128 890 180
rect 942 128 976 180
rect 1028 128 1054 180
rect 1106 128 1136 180
rect 1188 128 1216 180
rect 868 120 1216 128
rect 1296 92 1354 250
rect 1434 92 1492 246
rect 1572 180 1920 186
rect 1572 128 1594 180
rect 1646 128 1680 180
rect 1732 128 1758 180
rect 1810 128 1840 180
rect 1892 128 1920 180
rect 1572 120 1920 128
rect 2000 92 2058 250
rect 2138 186 2196 246
rect 2252 186 2304 220
rect 2338 186 2390 220
rect 2424 186 2476 220
rect 2510 186 2562 220
rect 2596 186 2648 220
rect 2704 186 2762 250
rect 2138 148 2278 186
rect 2618 148 2762 186
rect 2138 92 2762 148
rect 2842 92 2900 246
rect 2980 180 3328 186
rect 2980 128 3002 180
rect 3054 128 3088 180
rect 3140 128 3166 180
rect 3218 128 3248 180
rect 3300 128 3328 180
rect 2980 120 3328 128
rect 3408 92 3466 250
rect 3546 92 3604 246
rect 3684 180 4032 186
rect 3684 128 3706 180
rect 3758 128 3792 180
rect 3844 128 3870 180
rect 3922 128 3952 180
rect 4004 128 4032 180
rect 3684 120 4032 128
rect 4112 92 4170 250
rect 4250 186 4308 220
rect 4364 186 4416 220
rect 4450 186 4502 220
rect 4536 186 4588 220
rect 4622 186 4674 220
rect 4708 186 4760 220
rect 4816 186 4874 220
rect 4250 128 4390 186
rect 4732 128 4874 186
rect 4250 92 4874 128
rect 26 72 4874 92
rect 26 38 72 72
rect 106 38 146 72
rect 180 38 220 72
rect 254 38 294 72
rect 328 38 368 72
rect 402 38 442 72
rect 476 38 516 72
rect 550 38 590 72
rect 624 38 664 72
rect 698 38 738 72
rect 772 38 812 72
rect 846 38 886 72
rect 920 38 960 72
rect 994 38 1034 72
rect 1068 38 1108 72
rect 1142 38 1182 72
rect 1216 38 1256 72
rect 1290 38 1330 72
rect 1364 38 1404 72
rect 1438 38 1478 72
rect 1512 38 1552 72
rect 1586 38 1626 72
rect 1660 38 1700 72
rect 1734 38 1774 72
rect 1808 38 1848 72
rect 1882 38 1922 72
rect 1956 38 1996 72
rect 2030 38 2070 72
rect 2104 38 2144 72
rect 2178 38 2218 72
rect 2252 38 2292 72
rect 2326 38 2366 72
rect 2400 38 2440 72
rect 2474 38 2514 72
rect 2548 38 2588 72
rect 2622 38 2662 72
rect 2696 38 2736 72
rect 2770 38 2810 72
rect 2844 38 2884 72
rect 2918 38 2958 72
rect 2992 38 3032 72
rect 3066 38 3106 72
rect 3140 38 3180 72
rect 3214 38 3254 72
rect 3288 38 3328 72
rect 3362 38 3402 72
rect 3436 38 3476 72
rect 3510 38 3550 72
rect 3584 38 3624 72
rect 3658 38 3698 72
rect 3732 38 3772 72
rect 3806 38 3846 72
rect 3880 38 3920 72
rect 3954 38 3994 72
rect 4028 38 4068 72
rect 4102 38 4142 72
rect 4176 38 4216 72
rect 4250 38 4290 72
rect 4324 38 4364 72
rect 4398 38 4438 72
rect 4472 38 4512 72
rect 4546 38 4586 72
rect 4620 38 4660 72
rect 4694 38 4734 72
rect 4768 38 4808 72
rect 4842 38 4874 72
rect 26 26 4874 38
rect 834 -132 1058 26
rect 834 -188 856 -132
rect 912 -188 982 -132
rect 1038 -188 1058 -132
rect 834 -236 1058 -188
rect 834 -292 856 -236
rect 912 -292 982 -236
rect 1038 -292 1058 -236
rect 834 -320 1058 -292
rect 834 -376 856 -320
rect 912 -376 982 -320
rect 1038 -376 1058 -320
rect 834 -406 1058 -376
rect 834 -462 856 -406
rect 912 -462 982 -406
rect 1038 -462 1058 -406
rect 834 -500 1058 -462
rect 834 -556 856 -500
rect 912 -556 982 -500
rect 1038 -556 1058 -500
rect 834 -600 1058 -556
rect 834 -656 856 -600
rect 912 -656 982 -600
rect 1038 -656 1058 -600
rect 834 -684 1058 -656
rect 834 -740 856 -684
rect 912 -740 982 -684
rect 1038 -740 1058 -684
rect 834 -772 1058 -740
rect 1684 -132 1908 26
rect 1684 -188 1706 -132
rect 1762 -188 1832 -132
rect 1888 -188 1908 -132
rect 1684 -236 1908 -188
rect 1684 -292 1706 -236
rect 1762 -292 1832 -236
rect 1888 -292 1908 -236
rect 1684 -320 1908 -292
rect 1684 -376 1706 -320
rect 1762 -376 1832 -320
rect 1888 -376 1908 -320
rect 1684 -406 1908 -376
rect 1684 -462 1706 -406
rect 1762 -462 1832 -406
rect 1888 -462 1908 -406
rect 1684 -500 1908 -462
rect 1684 -556 1706 -500
rect 1762 -556 1832 -500
rect 1888 -556 1908 -500
rect 1684 -600 1908 -556
rect 1684 -656 1706 -600
rect 1762 -656 1832 -600
rect 1888 -656 1908 -600
rect 1684 -684 1908 -656
rect 1684 -740 1706 -684
rect 1762 -740 1832 -684
rect 1888 -740 1908 -684
rect 1684 -772 1908 -740
rect 2868 -132 3092 26
rect 2868 -188 2890 -132
rect 2946 -188 3016 -132
rect 3072 -188 3092 -132
rect 2868 -236 3092 -188
rect 2868 -292 2890 -236
rect 2946 -292 3016 -236
rect 3072 -292 3092 -236
rect 2868 -320 3092 -292
rect 2868 -376 2890 -320
rect 2946 -376 3016 -320
rect 3072 -376 3092 -320
rect 2868 -406 3092 -376
rect 2868 -462 2890 -406
rect 2946 -462 3016 -406
rect 3072 -462 3092 -406
rect 2868 -500 3092 -462
rect 2868 -556 2890 -500
rect 2946 -556 3016 -500
rect 3072 -556 3092 -500
rect 2868 -600 3092 -556
rect 2868 -656 2890 -600
rect 2946 -656 3016 -600
rect 3072 -656 3092 -600
rect 2868 -684 3092 -656
rect 2868 -740 2890 -684
rect 2946 -740 3016 -684
rect 3072 -740 3092 -684
rect 2868 -772 3092 -740
rect 3688 -132 3912 26
rect 3688 -188 3710 -132
rect 3766 -188 3836 -132
rect 3892 -188 3912 -132
rect 3688 -236 3912 -188
rect 3688 -292 3710 -236
rect 3766 -292 3836 -236
rect 3892 -292 3912 -236
rect 3688 -320 3912 -292
rect 3688 -376 3710 -320
rect 3766 -376 3836 -320
rect 3892 -376 3912 -320
rect 3688 -406 3912 -376
rect 3688 -462 3710 -406
rect 3766 -462 3836 -406
rect 3892 -462 3912 -406
rect 3688 -500 3912 -462
rect 3688 -556 3710 -500
rect 3766 -556 3836 -500
rect 3892 -556 3912 -500
rect 3688 -600 3912 -556
rect 3688 -656 3710 -600
rect 3766 -656 3836 -600
rect 3892 -656 3912 -600
rect 3688 -684 3912 -656
rect 3688 -740 3710 -684
rect 3766 -740 3836 -684
rect 3892 -740 3912 -684
rect 3688 -772 3912 -740
<< via1 >>
rect 888 2580 940 2632
rect 974 2580 1026 2632
rect 1052 2580 1104 2632
rect 1134 2580 1186 2632
rect 1592 2580 1644 2632
rect 1678 2580 1730 2632
rect 1756 2580 1808 2632
rect 1838 2580 1890 2632
rect 2298 2580 2350 2632
rect 2384 2580 2436 2632
rect 2462 2580 2514 2632
rect 2544 2580 2596 2632
rect 3002 2580 3054 2632
rect 3088 2580 3140 2632
rect 3166 2580 3218 2632
rect 3248 2580 3300 2632
rect 3706 2580 3758 2632
rect 3792 2580 3844 2632
rect 3870 2580 3922 2632
rect 3952 2580 4004 2632
rect 890 1438 942 1490
rect 976 1438 1028 1490
rect 1054 1438 1106 1490
rect 1136 1438 1188 1490
rect 890 1272 942 1324
rect 976 1272 1028 1324
rect 1054 1272 1106 1324
rect 1136 1272 1188 1324
rect 1594 1438 1646 1490
rect 1680 1438 1732 1490
rect 1758 1438 1810 1490
rect 1840 1438 1892 1490
rect 1594 1272 1646 1324
rect 1680 1272 1732 1324
rect 1758 1272 1810 1324
rect 1840 1272 1892 1324
rect 2298 1438 2350 1490
rect 2384 1438 2436 1490
rect 2462 1438 2514 1490
rect 2544 1438 2596 1490
rect 3002 1438 3054 1490
rect 3088 1438 3140 1490
rect 3166 1438 3218 1490
rect 3248 1438 3300 1490
rect 3002 1272 3054 1324
rect 3088 1272 3140 1324
rect 3166 1272 3218 1324
rect 3248 1272 3300 1324
rect 3706 1438 3758 1490
rect 3792 1438 3844 1490
rect 3870 1438 3922 1490
rect 3952 1438 4004 1490
rect 3706 1272 3758 1324
rect 3792 1272 3844 1324
rect 3870 1272 3922 1324
rect 3952 1272 4004 1324
rect 890 128 942 180
rect 976 128 1028 180
rect 1054 128 1106 180
rect 1136 128 1188 180
rect 1594 128 1646 180
rect 1680 128 1732 180
rect 1758 128 1810 180
rect 1840 128 1892 180
rect 3002 128 3054 180
rect 3088 128 3140 180
rect 3166 128 3218 180
rect 3248 128 3300 180
rect 3706 128 3758 180
rect 3792 128 3844 180
rect 3870 128 3922 180
rect 3952 128 4004 180
rect 856 -188 912 -132
rect 982 -188 1038 -132
rect 856 -292 912 -236
rect 982 -292 1038 -236
rect 856 -376 912 -320
rect 982 -376 1038 -320
rect 856 -462 912 -406
rect 982 -462 1038 -406
rect 856 -556 912 -500
rect 982 -556 1038 -500
rect 856 -656 912 -600
rect 982 -656 1038 -600
rect 856 -740 912 -684
rect 982 -740 1038 -684
rect 1706 -188 1762 -132
rect 1832 -188 1888 -132
rect 1706 -292 1762 -236
rect 1832 -292 1888 -236
rect 1706 -376 1762 -320
rect 1832 -376 1888 -320
rect 1706 -462 1762 -406
rect 1832 -462 1888 -406
rect 1706 -556 1762 -500
rect 1832 -556 1888 -500
rect 1706 -656 1762 -600
rect 1832 -656 1888 -600
rect 1706 -740 1762 -684
rect 1832 -740 1888 -684
rect 2890 -188 2946 -132
rect 3016 -188 3072 -132
rect 2890 -292 2946 -236
rect 3016 -292 3072 -236
rect 2890 -376 2946 -320
rect 3016 -376 3072 -320
rect 2890 -462 2946 -406
rect 3016 -462 3072 -406
rect 2890 -556 2946 -500
rect 3016 -556 3072 -500
rect 2890 -656 2946 -600
rect 3016 -656 3072 -600
rect 2890 -740 2946 -684
rect 3016 -740 3072 -684
rect 3710 -188 3766 -132
rect 3836 -188 3892 -132
rect 3710 -292 3766 -236
rect 3836 -292 3892 -236
rect 3710 -376 3766 -320
rect 3836 -376 3892 -320
rect 3710 -462 3766 -406
rect 3836 -462 3892 -406
rect 3710 -556 3766 -500
rect 3836 -556 3892 -500
rect 3710 -656 3766 -600
rect 3836 -656 3892 -600
rect 3710 -740 3766 -684
rect 3836 -740 3892 -684
<< metal2 >>
rect 866 2660 1214 2666
rect 866 2604 876 2660
rect 932 2632 966 2660
rect 1022 2632 1056 2660
rect 1112 2632 1148 2660
rect 940 2604 966 2632
rect 866 2580 888 2604
rect 940 2580 974 2604
rect 1026 2580 1052 2632
rect 1112 2604 1134 2632
rect 1204 2604 1214 2660
rect 1104 2580 1134 2604
rect 1186 2580 1214 2604
rect 866 2572 1214 2580
rect 1570 2660 1918 2666
rect 1570 2604 1580 2660
rect 1636 2632 1670 2660
rect 1726 2632 1760 2660
rect 1816 2632 1852 2660
rect 1644 2604 1670 2632
rect 1570 2580 1592 2604
rect 1644 2580 1678 2604
rect 1730 2580 1756 2632
rect 1816 2604 1838 2632
rect 1908 2604 1918 2660
rect 1808 2580 1838 2604
rect 1890 2580 1918 2604
rect 1570 2572 1918 2580
rect 2276 2660 2624 2666
rect 2276 2604 2286 2660
rect 2342 2632 2376 2660
rect 2432 2632 2466 2660
rect 2522 2632 2558 2660
rect 2350 2604 2376 2632
rect 2276 2580 2298 2604
rect 2350 2580 2384 2604
rect 2436 2580 2462 2632
rect 2522 2604 2544 2632
rect 2614 2604 2624 2660
rect 2514 2580 2544 2604
rect 2596 2580 2624 2604
rect 2276 2572 2624 2580
rect 2980 2660 3328 2666
rect 2980 2604 2990 2660
rect 3046 2632 3080 2660
rect 3136 2632 3170 2660
rect 3226 2632 3262 2660
rect 3054 2604 3080 2632
rect 2980 2580 3002 2604
rect 3054 2580 3088 2604
rect 3140 2580 3166 2632
rect 3226 2604 3248 2632
rect 3318 2604 3328 2660
rect 3218 2580 3248 2604
rect 3300 2580 3328 2604
rect 2980 2572 3328 2580
rect 3684 2660 4032 2666
rect 3684 2604 3694 2660
rect 3750 2632 3784 2660
rect 3840 2632 3874 2660
rect 3930 2632 3966 2660
rect 3758 2604 3784 2632
rect 3684 2580 3706 2604
rect 3758 2580 3792 2604
rect 3844 2580 3870 2632
rect 3930 2604 3952 2632
rect 4022 2604 4032 2660
rect 3922 2580 3952 2604
rect 4004 2580 4032 2604
rect 3684 2572 4032 2580
rect 226 -772 450 2538
rect 842 2518 1242 2538
rect 842 2462 894 2518
rect 950 2462 974 2518
rect 1030 2462 1054 2518
rect 1110 2462 1134 2518
rect 1190 2462 1242 2518
rect 842 2438 1242 2462
rect 842 2382 894 2438
rect 950 2382 974 2438
rect 1030 2382 1054 2438
rect 1110 2382 1134 2438
rect 1190 2382 1242 2438
rect 842 2358 1242 2382
rect 842 2302 894 2358
rect 950 2302 974 2358
rect 1030 2302 1054 2358
rect 1110 2302 1134 2358
rect 1190 2302 1242 2358
rect 842 2278 1242 2302
rect 842 2222 894 2278
rect 950 2222 974 2278
rect 1030 2222 1054 2278
rect 1110 2222 1134 2278
rect 1190 2222 1242 2278
rect 842 2202 1242 2222
rect 1546 2518 1946 2538
rect 1546 2462 1598 2518
rect 1654 2462 1678 2518
rect 1734 2462 1758 2518
rect 1814 2462 1838 2518
rect 1894 2462 1946 2518
rect 1546 2438 1946 2462
rect 1546 2382 1598 2438
rect 1654 2382 1678 2438
rect 1734 2382 1758 2438
rect 1814 2382 1838 2438
rect 1894 2382 1946 2438
rect 1546 2358 1946 2382
rect 1546 2302 1598 2358
rect 1654 2302 1678 2358
rect 1734 2302 1758 2358
rect 1814 2302 1838 2358
rect 1894 2302 1946 2358
rect 1546 2278 1946 2302
rect 1546 2222 1598 2278
rect 1654 2222 1678 2278
rect 1734 2222 1758 2278
rect 1814 2222 1838 2278
rect 1894 2222 1946 2278
rect 1546 2202 1946 2222
rect 2250 2518 2650 2538
rect 2250 2462 2302 2518
rect 2358 2462 2382 2518
rect 2438 2462 2462 2518
rect 2518 2462 2542 2518
rect 2598 2462 2650 2518
rect 2250 2438 2650 2462
rect 2250 2382 2302 2438
rect 2358 2382 2382 2438
rect 2438 2382 2462 2438
rect 2518 2382 2542 2438
rect 2598 2382 2650 2438
rect 2250 2358 2650 2382
rect 2250 2302 2302 2358
rect 2358 2302 2382 2358
rect 2438 2302 2462 2358
rect 2518 2302 2542 2358
rect 2598 2302 2650 2358
rect 2250 2278 2650 2302
rect 2250 2222 2302 2278
rect 2358 2222 2382 2278
rect 2438 2222 2462 2278
rect 2518 2222 2542 2278
rect 2598 2222 2650 2278
rect 2250 2202 2650 2222
rect 2954 2518 3354 2538
rect 2954 2462 3006 2518
rect 3062 2462 3086 2518
rect 3142 2462 3166 2518
rect 3222 2462 3246 2518
rect 3302 2462 3354 2518
rect 2954 2438 3354 2462
rect 2954 2382 3006 2438
rect 3062 2382 3086 2438
rect 3142 2382 3166 2438
rect 3222 2382 3246 2438
rect 3302 2382 3354 2438
rect 2954 2358 3354 2382
rect 2954 2302 3006 2358
rect 3062 2302 3086 2358
rect 3142 2302 3166 2358
rect 3222 2302 3246 2358
rect 3302 2302 3354 2358
rect 2954 2278 3354 2302
rect 2954 2222 3006 2278
rect 3062 2222 3086 2278
rect 3142 2222 3166 2278
rect 3222 2222 3246 2278
rect 3302 2222 3354 2278
rect 2954 2202 3354 2222
rect 3658 2518 4058 2538
rect 3658 2462 3710 2518
rect 3766 2462 3790 2518
rect 3846 2462 3870 2518
rect 3926 2462 3950 2518
rect 4006 2462 4058 2518
rect 3658 2438 4058 2462
rect 3658 2382 3710 2438
rect 3766 2382 3790 2438
rect 3846 2382 3870 2438
rect 3926 2382 3950 2438
rect 4006 2382 4058 2438
rect 3658 2358 4058 2382
rect 3658 2302 3710 2358
rect 3766 2302 3790 2358
rect 3846 2302 3870 2358
rect 3926 2302 3950 2358
rect 4006 2302 4058 2358
rect 3658 2278 4058 2302
rect 3658 2222 3710 2278
rect 3766 2222 3790 2278
rect 3846 2222 3870 2278
rect 3926 2222 3950 2278
rect 4006 2222 4058 2278
rect 3658 2202 4058 2222
rect 842 1858 1242 1878
rect 842 1802 894 1858
rect 950 1802 974 1858
rect 1030 1802 1054 1858
rect 1110 1802 1134 1858
rect 1190 1802 1242 1858
rect 842 1778 1242 1802
rect 842 1722 894 1778
rect 950 1722 974 1778
rect 1030 1722 1054 1778
rect 1110 1722 1134 1778
rect 1190 1722 1242 1778
rect 842 1698 1242 1722
rect 842 1642 894 1698
rect 950 1642 974 1698
rect 1030 1642 1054 1698
rect 1110 1642 1134 1698
rect 1190 1642 1242 1698
rect 842 1618 1242 1642
rect 842 1562 894 1618
rect 950 1562 974 1618
rect 1030 1562 1054 1618
rect 1110 1562 1134 1618
rect 1190 1562 1242 1618
rect 842 1542 1242 1562
rect 1546 1858 1946 1878
rect 1546 1802 1598 1858
rect 1654 1802 1678 1858
rect 1734 1802 1758 1858
rect 1814 1802 1838 1858
rect 1894 1802 1946 1858
rect 1546 1778 1946 1802
rect 1546 1722 1598 1778
rect 1654 1722 1678 1778
rect 1734 1722 1758 1778
rect 1814 1722 1838 1778
rect 1894 1722 1946 1778
rect 1546 1698 1946 1722
rect 1546 1642 1598 1698
rect 1654 1642 1678 1698
rect 1734 1642 1758 1698
rect 1814 1642 1838 1698
rect 1894 1642 1946 1698
rect 1546 1618 1946 1642
rect 1546 1562 1598 1618
rect 1654 1562 1678 1618
rect 1734 1562 1758 1618
rect 1814 1562 1838 1618
rect 1894 1562 1946 1618
rect 1546 1542 1946 1562
rect 2250 1858 2650 1878
rect 2250 1802 2302 1858
rect 2358 1802 2382 1858
rect 2438 1802 2462 1858
rect 2518 1802 2542 1858
rect 2598 1802 2650 1858
rect 2250 1778 2650 1802
rect 2250 1722 2302 1778
rect 2358 1722 2382 1778
rect 2438 1722 2462 1778
rect 2518 1722 2542 1778
rect 2598 1722 2650 1778
rect 2250 1698 2650 1722
rect 2250 1642 2302 1698
rect 2358 1642 2382 1698
rect 2438 1642 2462 1698
rect 2518 1642 2542 1698
rect 2598 1642 2650 1698
rect 2250 1618 2650 1642
rect 2250 1562 2302 1618
rect 2358 1562 2382 1618
rect 2438 1562 2462 1618
rect 2518 1562 2542 1618
rect 2598 1562 2650 1618
rect 2250 1542 2650 1562
rect 2954 1858 3354 1878
rect 2954 1802 3006 1858
rect 3062 1802 3086 1858
rect 3142 1802 3166 1858
rect 3222 1802 3246 1858
rect 3302 1802 3354 1858
rect 2954 1778 3354 1802
rect 2954 1722 3006 1778
rect 3062 1722 3086 1778
rect 3142 1722 3166 1778
rect 3222 1722 3246 1778
rect 3302 1722 3354 1778
rect 2954 1698 3354 1722
rect 2954 1642 3006 1698
rect 3062 1642 3086 1698
rect 3142 1642 3166 1698
rect 3222 1642 3246 1698
rect 3302 1642 3354 1698
rect 2954 1618 3354 1642
rect 2954 1562 3006 1618
rect 3062 1562 3086 1618
rect 3142 1562 3166 1618
rect 3222 1562 3246 1618
rect 3302 1562 3354 1618
rect 2954 1542 3354 1562
rect 3658 1858 4058 1878
rect 3658 1802 3710 1858
rect 3766 1802 3790 1858
rect 3846 1802 3870 1858
rect 3926 1802 3950 1858
rect 4006 1802 4058 1858
rect 3658 1778 4058 1802
rect 3658 1722 3710 1778
rect 3766 1722 3790 1778
rect 3846 1722 3870 1778
rect 3926 1722 3950 1778
rect 4006 1722 4058 1778
rect 3658 1698 4058 1722
rect 3658 1642 3710 1698
rect 3766 1642 3790 1698
rect 3846 1642 3870 1698
rect 3926 1642 3950 1698
rect 4006 1642 4058 1698
rect 3658 1618 4058 1642
rect 3658 1562 3710 1618
rect 3766 1562 3790 1618
rect 3846 1562 3870 1618
rect 3926 1562 3950 1618
rect 4006 1562 4058 1618
rect 3658 1542 4058 1562
rect 868 1490 1216 1508
rect 868 1476 890 1490
rect 942 1476 976 1490
rect 868 1420 878 1476
rect 942 1438 968 1476
rect 1028 1438 1054 1490
rect 1106 1476 1136 1490
rect 1188 1476 1216 1490
rect 1114 1438 1136 1476
rect 934 1420 968 1438
rect 1024 1420 1058 1438
rect 1114 1420 1150 1438
rect 1206 1420 1216 1476
rect 868 1414 1216 1420
rect 1572 1490 1920 1508
rect 1572 1476 1594 1490
rect 1646 1476 1680 1490
rect 1572 1420 1582 1476
rect 1646 1438 1672 1476
rect 1732 1438 1758 1490
rect 1810 1476 1840 1490
rect 1892 1476 1920 1490
rect 1818 1438 1840 1476
rect 1638 1420 1672 1438
rect 1728 1420 1762 1438
rect 1818 1420 1854 1438
rect 1910 1420 1920 1476
rect 1572 1414 1920 1420
rect 2276 1490 2624 1508
rect 2276 1476 2298 1490
rect 2350 1476 2384 1490
rect 2276 1420 2286 1476
rect 2350 1438 2376 1476
rect 2436 1438 2462 1490
rect 2514 1476 2544 1490
rect 2596 1476 2624 1490
rect 2522 1438 2544 1476
rect 2342 1420 2376 1438
rect 2432 1420 2466 1438
rect 2522 1420 2558 1438
rect 2614 1420 2624 1476
rect 2276 1414 2624 1420
rect 2980 1490 3328 1508
rect 2980 1476 3002 1490
rect 3054 1476 3088 1490
rect 2980 1420 2990 1476
rect 3054 1438 3080 1476
rect 3140 1438 3166 1490
rect 3218 1476 3248 1490
rect 3300 1476 3328 1490
rect 3226 1438 3248 1476
rect 3046 1420 3080 1438
rect 3136 1420 3170 1438
rect 3226 1420 3262 1438
rect 3318 1420 3328 1476
rect 2980 1414 3328 1420
rect 3684 1490 4032 1508
rect 3684 1476 3706 1490
rect 3758 1476 3792 1490
rect 3684 1420 3694 1476
rect 3758 1438 3784 1476
rect 3844 1438 3870 1490
rect 3922 1476 3952 1490
rect 4004 1476 4032 1490
rect 3930 1438 3952 1476
rect 3750 1420 3784 1438
rect 3840 1420 3874 1438
rect 3930 1420 3966 1438
rect 4022 1420 4032 1476
rect 3684 1414 4032 1420
rect 868 1336 1216 1342
rect 868 1280 878 1336
rect 934 1324 968 1336
rect 1024 1324 1058 1336
rect 1114 1324 1150 1336
rect 942 1280 968 1324
rect 868 1272 890 1280
rect 942 1272 976 1280
rect 1028 1272 1054 1324
rect 1114 1280 1136 1324
rect 1206 1280 1216 1336
rect 1106 1272 1136 1280
rect 1188 1272 1216 1280
rect 868 1248 1216 1272
rect 1572 1336 1920 1342
rect 1572 1280 1582 1336
rect 1638 1324 1672 1336
rect 1728 1324 1762 1336
rect 1818 1324 1854 1336
rect 1646 1280 1672 1324
rect 1572 1272 1594 1280
rect 1646 1272 1680 1280
rect 1732 1272 1758 1324
rect 1818 1280 1840 1324
rect 1910 1280 1920 1336
rect 1810 1272 1840 1280
rect 1892 1272 1920 1280
rect 1572 1248 1920 1272
rect 2980 1336 3328 1342
rect 2980 1280 2990 1336
rect 3046 1324 3080 1336
rect 3136 1324 3170 1336
rect 3226 1324 3262 1336
rect 3054 1280 3080 1324
rect 2980 1272 3002 1280
rect 3054 1272 3088 1280
rect 3140 1272 3166 1324
rect 3226 1280 3248 1324
rect 3318 1280 3328 1336
rect 3218 1272 3248 1280
rect 3300 1272 3328 1280
rect 2980 1248 3328 1272
rect 3684 1336 4032 1342
rect 3684 1280 3694 1336
rect 3750 1324 3784 1336
rect 3840 1324 3874 1336
rect 3930 1324 3966 1336
rect 3758 1280 3784 1324
rect 3684 1272 3706 1280
rect 3758 1272 3792 1280
rect 3844 1272 3870 1324
rect 3930 1280 3952 1324
rect 4022 1280 4032 1336
rect 3922 1272 3952 1280
rect 4004 1272 4032 1280
rect 3684 1248 4032 1272
rect 842 1194 1242 1214
rect 842 1138 894 1194
rect 950 1138 974 1194
rect 1030 1138 1054 1194
rect 1110 1138 1134 1194
rect 1190 1138 1242 1194
rect 842 1114 1242 1138
rect 842 1058 894 1114
rect 950 1058 974 1114
rect 1030 1058 1054 1114
rect 1110 1058 1134 1114
rect 1190 1058 1242 1114
rect 842 1034 1242 1058
rect 842 978 894 1034
rect 950 978 974 1034
rect 1030 978 1054 1034
rect 1110 978 1134 1034
rect 1190 978 1242 1034
rect 842 954 1242 978
rect 842 898 894 954
rect 950 898 974 954
rect 1030 898 1054 954
rect 1110 898 1134 954
rect 1190 898 1242 954
rect 842 878 1242 898
rect 1546 1194 1946 1214
rect 1546 1138 1598 1194
rect 1654 1138 1678 1194
rect 1734 1138 1758 1194
rect 1814 1138 1838 1194
rect 1894 1138 1946 1194
rect 1546 1114 1946 1138
rect 1546 1058 1598 1114
rect 1654 1058 1678 1114
rect 1734 1058 1758 1114
rect 1814 1058 1838 1114
rect 1894 1058 1946 1114
rect 1546 1034 1946 1058
rect 1546 978 1598 1034
rect 1654 978 1678 1034
rect 1734 978 1758 1034
rect 1814 978 1838 1034
rect 1894 978 1946 1034
rect 1546 954 1946 978
rect 1546 898 1598 954
rect 1654 898 1678 954
rect 1734 898 1758 954
rect 1814 898 1838 954
rect 1894 898 1946 954
rect 1546 878 1946 898
rect 842 536 1242 556
rect 842 480 894 536
rect 950 480 974 536
rect 1030 480 1054 536
rect 1110 480 1134 536
rect 1190 480 1242 536
rect 842 456 1242 480
rect 842 400 894 456
rect 950 400 974 456
rect 1030 400 1054 456
rect 1110 400 1134 456
rect 1190 400 1242 456
rect 842 376 1242 400
rect 842 320 894 376
rect 950 320 974 376
rect 1030 320 1054 376
rect 1110 320 1134 376
rect 1190 320 1242 376
rect 842 296 1242 320
rect 842 240 894 296
rect 950 240 974 296
rect 1030 240 1054 296
rect 1110 240 1134 296
rect 1190 240 1242 296
rect 842 220 1242 240
rect 1546 536 1946 556
rect 1546 480 1598 536
rect 1654 480 1678 536
rect 1734 480 1758 536
rect 1814 480 1838 536
rect 1894 480 1946 536
rect 1546 456 1946 480
rect 1546 400 1598 456
rect 1654 400 1678 456
rect 1734 400 1758 456
rect 1814 400 1838 456
rect 1894 400 1946 456
rect 1546 376 1946 400
rect 1546 320 1598 376
rect 1654 320 1678 376
rect 1734 320 1758 376
rect 1814 320 1838 376
rect 1894 320 1946 376
rect 1546 296 1946 320
rect 1546 240 1598 296
rect 1654 240 1678 296
rect 1734 240 1758 296
rect 1814 240 1838 296
rect 1894 240 1946 296
rect 1546 220 1946 240
rect 868 180 1216 186
rect 868 154 890 180
rect 942 154 976 180
rect 868 98 878 154
rect 942 128 968 154
rect 1028 128 1054 180
rect 1106 154 1136 180
rect 1188 154 1216 180
rect 1114 128 1136 154
rect 934 98 968 128
rect 1024 98 1058 128
rect 1114 98 1150 128
rect 1206 98 1216 154
rect 868 92 1216 98
rect 1572 180 1920 186
rect 1572 154 1594 180
rect 1646 154 1680 180
rect 1572 98 1582 154
rect 1646 128 1672 154
rect 1732 128 1758 180
rect 1810 154 1840 180
rect 1892 154 1920 180
rect 1818 128 1840 154
rect 1638 98 1672 128
rect 1728 98 1762 128
rect 1818 98 1854 128
rect 1910 98 1920 154
rect 1572 92 1920 98
rect 834 -130 1058 -100
rect 834 -190 854 -130
rect 914 -190 980 -130
rect 1040 -190 1058 -130
rect 834 -234 1058 -190
rect 834 -294 854 -234
rect 914 -294 980 -234
rect 1040 -294 1058 -234
rect 834 -318 1058 -294
rect 834 -378 854 -318
rect 914 -378 980 -318
rect 1040 -378 1058 -318
rect 834 -404 1058 -378
rect 834 -464 854 -404
rect 914 -464 980 -404
rect 1040 -464 1058 -404
rect 834 -498 1058 -464
rect 834 -558 854 -498
rect 914 -558 980 -498
rect 1040 -558 1058 -498
rect 834 -598 1058 -558
rect 834 -658 854 -598
rect 914 -658 980 -598
rect 1040 -658 1058 -598
rect 834 -682 1058 -658
rect 834 -742 854 -682
rect 914 -742 980 -682
rect 1040 -742 1058 -682
rect 834 -772 1058 -742
rect 1684 -130 1908 -100
rect 1684 -190 1704 -130
rect 1764 -190 1830 -130
rect 1890 -190 1908 -130
rect 1684 -234 1908 -190
rect 1684 -294 1704 -234
rect 1764 -294 1830 -234
rect 1890 -294 1908 -234
rect 1684 -318 1908 -294
rect 1684 -378 1704 -318
rect 1764 -378 1830 -318
rect 1890 -378 1908 -318
rect 1684 -404 1908 -378
rect 1684 -464 1704 -404
rect 1764 -464 1830 -404
rect 1890 -464 1908 -404
rect 1684 -498 1908 -464
rect 1684 -558 1704 -498
rect 1764 -558 1830 -498
rect 1890 -558 1908 -498
rect 1684 -598 1908 -558
rect 1684 -658 1704 -598
rect 1764 -658 1830 -598
rect 1890 -658 1908 -598
rect 1684 -682 1908 -658
rect 1684 -742 1704 -682
rect 1764 -742 1830 -682
rect 1890 -742 1908 -682
rect 1684 -772 1908 -742
rect 2354 -130 2578 1216
rect 2954 1194 3354 1214
rect 2954 1138 3006 1194
rect 3062 1138 3086 1194
rect 3142 1138 3166 1194
rect 3222 1138 3246 1194
rect 3302 1138 3354 1194
rect 2954 1114 3354 1138
rect 2954 1058 3006 1114
rect 3062 1058 3086 1114
rect 3142 1058 3166 1114
rect 3222 1058 3246 1114
rect 3302 1058 3354 1114
rect 2954 1034 3354 1058
rect 2954 978 3006 1034
rect 3062 978 3086 1034
rect 3142 978 3166 1034
rect 3222 978 3246 1034
rect 3302 978 3354 1034
rect 2954 954 3354 978
rect 2954 898 3006 954
rect 3062 898 3086 954
rect 3142 898 3166 954
rect 3222 898 3246 954
rect 3302 898 3354 954
rect 2954 878 3354 898
rect 3658 1194 4058 1214
rect 3658 1138 3710 1194
rect 3766 1138 3790 1194
rect 3846 1138 3870 1194
rect 3926 1138 3950 1194
rect 4006 1138 4058 1194
rect 3658 1114 4058 1138
rect 3658 1058 3710 1114
rect 3766 1058 3790 1114
rect 3846 1058 3870 1114
rect 3926 1058 3950 1114
rect 4006 1058 4058 1114
rect 3658 1034 4058 1058
rect 3658 978 3710 1034
rect 3766 978 3790 1034
rect 3846 978 3870 1034
rect 3926 978 3950 1034
rect 4006 978 4058 1034
rect 3658 954 4058 978
rect 3658 898 3710 954
rect 3766 898 3790 954
rect 3846 898 3870 954
rect 3926 898 3950 954
rect 4006 898 4058 954
rect 3658 878 4058 898
rect 2954 536 3354 556
rect 2954 480 3006 536
rect 3062 480 3086 536
rect 3142 480 3166 536
rect 3222 480 3246 536
rect 3302 480 3354 536
rect 2954 456 3354 480
rect 2954 400 3006 456
rect 3062 400 3086 456
rect 3142 400 3166 456
rect 3222 400 3246 456
rect 3302 400 3354 456
rect 2954 376 3354 400
rect 2954 320 3006 376
rect 3062 320 3086 376
rect 3142 320 3166 376
rect 3222 320 3246 376
rect 3302 320 3354 376
rect 2954 296 3354 320
rect 2954 240 3006 296
rect 3062 240 3086 296
rect 3142 240 3166 296
rect 3222 240 3246 296
rect 3302 240 3354 296
rect 2954 220 3354 240
rect 3658 536 4058 556
rect 3658 480 3710 536
rect 3766 480 3790 536
rect 3846 480 3870 536
rect 3926 480 3950 536
rect 4006 480 4058 536
rect 3658 456 4058 480
rect 3658 400 3710 456
rect 3766 400 3790 456
rect 3846 400 3870 456
rect 3926 400 3950 456
rect 4006 400 4058 456
rect 3658 376 4058 400
rect 3658 320 3710 376
rect 3766 320 3790 376
rect 3846 320 3870 376
rect 3926 320 3950 376
rect 4006 320 4058 376
rect 3658 296 4058 320
rect 3658 240 3710 296
rect 3766 240 3790 296
rect 3846 240 3870 296
rect 3926 240 3950 296
rect 4006 240 4058 296
rect 3658 220 4058 240
rect 2980 180 3328 186
rect 2980 154 3002 180
rect 3054 154 3088 180
rect 2980 98 2990 154
rect 3054 128 3080 154
rect 3140 128 3166 180
rect 3218 154 3248 180
rect 3300 154 3328 180
rect 3226 128 3248 154
rect 3046 98 3080 128
rect 3136 98 3170 128
rect 3226 98 3262 128
rect 3318 98 3328 154
rect 2980 92 3328 98
rect 3684 180 4032 186
rect 3684 154 3706 180
rect 3758 154 3792 180
rect 3684 98 3694 154
rect 3758 128 3784 154
rect 3844 128 3870 180
rect 3922 154 3952 180
rect 4004 154 4032 180
rect 3930 128 3952 154
rect 3750 98 3784 128
rect 3840 98 3874 128
rect 3930 98 3966 128
rect 4022 98 4032 154
rect 3684 92 4032 98
rect 2354 -190 2374 -130
rect 2434 -190 2500 -130
rect 2560 -190 2578 -130
rect 2354 -234 2578 -190
rect 2354 -294 2374 -234
rect 2434 -294 2500 -234
rect 2560 -294 2578 -234
rect 2354 -318 2578 -294
rect 2354 -378 2374 -318
rect 2434 -378 2500 -318
rect 2560 -378 2578 -318
rect 2354 -404 2578 -378
rect 2354 -464 2374 -404
rect 2434 -464 2500 -404
rect 2560 -464 2578 -404
rect 2354 -498 2578 -464
rect 2354 -558 2374 -498
rect 2434 -558 2500 -498
rect 2560 -558 2578 -498
rect 2354 -598 2578 -558
rect 2354 -658 2374 -598
rect 2434 -658 2500 -598
rect 2560 -658 2578 -598
rect 2354 -682 2578 -658
rect 2354 -742 2374 -682
rect 2434 -742 2500 -682
rect 2560 -742 2578 -682
rect 2354 -770 2578 -742
rect 2868 -130 3092 -100
rect 2868 -190 2888 -130
rect 2948 -190 3014 -130
rect 3074 -190 3092 -130
rect 2868 -234 3092 -190
rect 2868 -294 2888 -234
rect 2948 -294 3014 -234
rect 3074 -294 3092 -234
rect 2868 -318 3092 -294
rect 2868 -378 2888 -318
rect 2948 -378 3014 -318
rect 3074 -378 3092 -318
rect 2868 -404 3092 -378
rect 2868 -464 2888 -404
rect 2948 -464 3014 -404
rect 3074 -464 3092 -404
rect 2868 -498 3092 -464
rect 2868 -558 2888 -498
rect 2948 -558 3014 -498
rect 3074 -558 3092 -498
rect 2868 -598 3092 -558
rect 2868 -658 2888 -598
rect 2948 -658 3014 -598
rect 3074 -658 3092 -598
rect 2868 -682 3092 -658
rect 2868 -742 2888 -682
rect 2948 -742 3014 -682
rect 3074 -742 3092 -682
rect 2868 -772 3092 -742
rect 3688 -130 3912 -100
rect 3688 -190 3708 -130
rect 3768 -190 3834 -130
rect 3894 -190 3912 -130
rect 3688 -234 3912 -190
rect 3688 -294 3708 -234
rect 3768 -294 3834 -234
rect 3894 -294 3912 -234
rect 3688 -318 3912 -294
rect 3688 -378 3708 -318
rect 3768 -378 3834 -318
rect 3894 -378 3912 -318
rect 3688 -404 3912 -378
rect 3688 -464 3708 -404
rect 3768 -464 3834 -404
rect 3894 -464 3912 -404
rect 3688 -498 3912 -464
rect 3688 -558 3708 -498
rect 3768 -558 3834 -498
rect 3894 -558 3912 -498
rect 3688 -598 3912 -558
rect 3688 -658 3708 -598
rect 3768 -658 3834 -598
rect 3894 -658 3912 -598
rect 3688 -682 3912 -658
rect 3688 -742 3708 -682
rect 3768 -742 3834 -682
rect 3894 -742 3912 -682
rect 3688 -772 3912 -742
rect 4446 -772 4670 2540
<< via2 >>
rect 876 2632 932 2660
rect 966 2632 1022 2660
rect 1056 2632 1112 2660
rect 1148 2632 1204 2660
rect 876 2604 888 2632
rect 888 2604 932 2632
rect 966 2604 974 2632
rect 974 2604 1022 2632
rect 1056 2604 1104 2632
rect 1104 2604 1112 2632
rect 1148 2604 1186 2632
rect 1186 2604 1204 2632
rect 1580 2632 1636 2660
rect 1670 2632 1726 2660
rect 1760 2632 1816 2660
rect 1852 2632 1908 2660
rect 1580 2604 1592 2632
rect 1592 2604 1636 2632
rect 1670 2604 1678 2632
rect 1678 2604 1726 2632
rect 1760 2604 1808 2632
rect 1808 2604 1816 2632
rect 1852 2604 1890 2632
rect 1890 2604 1908 2632
rect 2286 2632 2342 2660
rect 2376 2632 2432 2660
rect 2466 2632 2522 2660
rect 2558 2632 2614 2660
rect 2286 2604 2298 2632
rect 2298 2604 2342 2632
rect 2376 2604 2384 2632
rect 2384 2604 2432 2632
rect 2466 2604 2514 2632
rect 2514 2604 2522 2632
rect 2558 2604 2596 2632
rect 2596 2604 2614 2632
rect 2990 2632 3046 2660
rect 3080 2632 3136 2660
rect 3170 2632 3226 2660
rect 3262 2632 3318 2660
rect 2990 2604 3002 2632
rect 3002 2604 3046 2632
rect 3080 2604 3088 2632
rect 3088 2604 3136 2632
rect 3170 2604 3218 2632
rect 3218 2604 3226 2632
rect 3262 2604 3300 2632
rect 3300 2604 3318 2632
rect 3694 2632 3750 2660
rect 3784 2632 3840 2660
rect 3874 2632 3930 2660
rect 3966 2632 4022 2660
rect 3694 2604 3706 2632
rect 3706 2604 3750 2632
rect 3784 2604 3792 2632
rect 3792 2604 3840 2632
rect 3874 2604 3922 2632
rect 3922 2604 3930 2632
rect 3966 2604 4004 2632
rect 4004 2604 4022 2632
rect 894 2462 950 2518
rect 974 2462 1030 2518
rect 1054 2462 1110 2518
rect 1134 2462 1190 2518
rect 894 2382 950 2438
rect 974 2382 1030 2438
rect 1054 2382 1110 2438
rect 1134 2382 1190 2438
rect 894 2302 950 2358
rect 974 2302 1030 2358
rect 1054 2302 1110 2358
rect 1134 2302 1190 2358
rect 894 2222 950 2278
rect 974 2222 1030 2278
rect 1054 2222 1110 2278
rect 1134 2222 1190 2278
rect 1598 2462 1654 2518
rect 1678 2462 1734 2518
rect 1758 2462 1814 2518
rect 1838 2462 1894 2518
rect 1598 2382 1654 2438
rect 1678 2382 1734 2438
rect 1758 2382 1814 2438
rect 1838 2382 1894 2438
rect 1598 2302 1654 2358
rect 1678 2302 1734 2358
rect 1758 2302 1814 2358
rect 1838 2302 1894 2358
rect 1598 2222 1654 2278
rect 1678 2222 1734 2278
rect 1758 2222 1814 2278
rect 1838 2222 1894 2278
rect 2302 2462 2358 2518
rect 2382 2462 2438 2518
rect 2462 2462 2518 2518
rect 2542 2462 2598 2518
rect 2302 2382 2358 2438
rect 2382 2382 2438 2438
rect 2462 2382 2518 2438
rect 2542 2382 2598 2438
rect 2302 2302 2358 2358
rect 2382 2302 2438 2358
rect 2462 2302 2518 2358
rect 2542 2302 2598 2358
rect 2302 2222 2358 2278
rect 2382 2222 2438 2278
rect 2462 2222 2518 2278
rect 2542 2222 2598 2278
rect 3006 2462 3062 2518
rect 3086 2462 3142 2518
rect 3166 2462 3222 2518
rect 3246 2462 3302 2518
rect 3006 2382 3062 2438
rect 3086 2382 3142 2438
rect 3166 2382 3222 2438
rect 3246 2382 3302 2438
rect 3006 2302 3062 2358
rect 3086 2302 3142 2358
rect 3166 2302 3222 2358
rect 3246 2302 3302 2358
rect 3006 2222 3062 2278
rect 3086 2222 3142 2278
rect 3166 2222 3222 2278
rect 3246 2222 3302 2278
rect 3710 2462 3766 2518
rect 3790 2462 3846 2518
rect 3870 2462 3926 2518
rect 3950 2462 4006 2518
rect 3710 2382 3766 2438
rect 3790 2382 3846 2438
rect 3870 2382 3926 2438
rect 3950 2382 4006 2438
rect 3710 2302 3766 2358
rect 3790 2302 3846 2358
rect 3870 2302 3926 2358
rect 3950 2302 4006 2358
rect 3710 2222 3766 2278
rect 3790 2222 3846 2278
rect 3870 2222 3926 2278
rect 3950 2222 4006 2278
rect 894 1802 950 1858
rect 974 1802 1030 1858
rect 1054 1802 1110 1858
rect 1134 1802 1190 1858
rect 894 1722 950 1778
rect 974 1722 1030 1778
rect 1054 1722 1110 1778
rect 1134 1722 1190 1778
rect 894 1642 950 1698
rect 974 1642 1030 1698
rect 1054 1642 1110 1698
rect 1134 1642 1190 1698
rect 894 1562 950 1618
rect 974 1562 1030 1618
rect 1054 1562 1110 1618
rect 1134 1562 1190 1618
rect 1598 1802 1654 1858
rect 1678 1802 1734 1858
rect 1758 1802 1814 1858
rect 1838 1802 1894 1858
rect 1598 1722 1654 1778
rect 1678 1722 1734 1778
rect 1758 1722 1814 1778
rect 1838 1722 1894 1778
rect 1598 1642 1654 1698
rect 1678 1642 1734 1698
rect 1758 1642 1814 1698
rect 1838 1642 1894 1698
rect 1598 1562 1654 1618
rect 1678 1562 1734 1618
rect 1758 1562 1814 1618
rect 1838 1562 1894 1618
rect 2302 1802 2358 1858
rect 2382 1802 2438 1858
rect 2462 1802 2518 1858
rect 2542 1802 2598 1858
rect 2302 1722 2358 1778
rect 2382 1722 2438 1778
rect 2462 1722 2518 1778
rect 2542 1722 2598 1778
rect 2302 1642 2358 1698
rect 2382 1642 2438 1698
rect 2462 1642 2518 1698
rect 2542 1642 2598 1698
rect 2302 1562 2358 1618
rect 2382 1562 2438 1618
rect 2462 1562 2518 1618
rect 2542 1562 2598 1618
rect 3006 1802 3062 1858
rect 3086 1802 3142 1858
rect 3166 1802 3222 1858
rect 3246 1802 3302 1858
rect 3006 1722 3062 1778
rect 3086 1722 3142 1778
rect 3166 1722 3222 1778
rect 3246 1722 3302 1778
rect 3006 1642 3062 1698
rect 3086 1642 3142 1698
rect 3166 1642 3222 1698
rect 3246 1642 3302 1698
rect 3006 1562 3062 1618
rect 3086 1562 3142 1618
rect 3166 1562 3222 1618
rect 3246 1562 3302 1618
rect 3710 1802 3766 1858
rect 3790 1802 3846 1858
rect 3870 1802 3926 1858
rect 3950 1802 4006 1858
rect 3710 1722 3766 1778
rect 3790 1722 3846 1778
rect 3870 1722 3926 1778
rect 3950 1722 4006 1778
rect 3710 1642 3766 1698
rect 3790 1642 3846 1698
rect 3870 1642 3926 1698
rect 3950 1642 4006 1698
rect 3710 1562 3766 1618
rect 3790 1562 3846 1618
rect 3870 1562 3926 1618
rect 3950 1562 4006 1618
rect 878 1438 890 1476
rect 890 1438 934 1476
rect 968 1438 976 1476
rect 976 1438 1024 1476
rect 1058 1438 1106 1476
rect 1106 1438 1114 1476
rect 1150 1438 1188 1476
rect 1188 1438 1206 1476
rect 878 1420 934 1438
rect 968 1420 1024 1438
rect 1058 1420 1114 1438
rect 1150 1420 1206 1438
rect 1582 1438 1594 1476
rect 1594 1438 1638 1476
rect 1672 1438 1680 1476
rect 1680 1438 1728 1476
rect 1762 1438 1810 1476
rect 1810 1438 1818 1476
rect 1854 1438 1892 1476
rect 1892 1438 1910 1476
rect 1582 1420 1638 1438
rect 1672 1420 1728 1438
rect 1762 1420 1818 1438
rect 1854 1420 1910 1438
rect 2286 1438 2298 1476
rect 2298 1438 2342 1476
rect 2376 1438 2384 1476
rect 2384 1438 2432 1476
rect 2466 1438 2514 1476
rect 2514 1438 2522 1476
rect 2558 1438 2596 1476
rect 2596 1438 2614 1476
rect 2286 1420 2342 1438
rect 2376 1420 2432 1438
rect 2466 1420 2522 1438
rect 2558 1420 2614 1438
rect 2990 1438 3002 1476
rect 3002 1438 3046 1476
rect 3080 1438 3088 1476
rect 3088 1438 3136 1476
rect 3170 1438 3218 1476
rect 3218 1438 3226 1476
rect 3262 1438 3300 1476
rect 3300 1438 3318 1476
rect 2990 1420 3046 1438
rect 3080 1420 3136 1438
rect 3170 1420 3226 1438
rect 3262 1420 3318 1438
rect 3694 1438 3706 1476
rect 3706 1438 3750 1476
rect 3784 1438 3792 1476
rect 3792 1438 3840 1476
rect 3874 1438 3922 1476
rect 3922 1438 3930 1476
rect 3966 1438 4004 1476
rect 4004 1438 4022 1476
rect 3694 1420 3750 1438
rect 3784 1420 3840 1438
rect 3874 1420 3930 1438
rect 3966 1420 4022 1438
rect 878 1324 934 1336
rect 968 1324 1024 1336
rect 1058 1324 1114 1336
rect 1150 1324 1206 1336
rect 878 1280 890 1324
rect 890 1280 934 1324
rect 968 1280 976 1324
rect 976 1280 1024 1324
rect 1058 1280 1106 1324
rect 1106 1280 1114 1324
rect 1150 1280 1188 1324
rect 1188 1280 1206 1324
rect 1582 1324 1638 1336
rect 1672 1324 1728 1336
rect 1762 1324 1818 1336
rect 1854 1324 1910 1336
rect 1582 1280 1594 1324
rect 1594 1280 1638 1324
rect 1672 1280 1680 1324
rect 1680 1280 1728 1324
rect 1762 1280 1810 1324
rect 1810 1280 1818 1324
rect 1854 1280 1892 1324
rect 1892 1280 1910 1324
rect 2990 1324 3046 1336
rect 3080 1324 3136 1336
rect 3170 1324 3226 1336
rect 3262 1324 3318 1336
rect 2990 1280 3002 1324
rect 3002 1280 3046 1324
rect 3080 1280 3088 1324
rect 3088 1280 3136 1324
rect 3170 1280 3218 1324
rect 3218 1280 3226 1324
rect 3262 1280 3300 1324
rect 3300 1280 3318 1324
rect 3694 1324 3750 1336
rect 3784 1324 3840 1336
rect 3874 1324 3930 1336
rect 3966 1324 4022 1336
rect 3694 1280 3706 1324
rect 3706 1280 3750 1324
rect 3784 1280 3792 1324
rect 3792 1280 3840 1324
rect 3874 1280 3922 1324
rect 3922 1280 3930 1324
rect 3966 1280 4004 1324
rect 4004 1280 4022 1324
rect 894 1138 950 1194
rect 974 1138 1030 1194
rect 1054 1138 1110 1194
rect 1134 1138 1190 1194
rect 894 1058 950 1114
rect 974 1058 1030 1114
rect 1054 1058 1110 1114
rect 1134 1058 1190 1114
rect 894 978 950 1034
rect 974 978 1030 1034
rect 1054 978 1110 1034
rect 1134 978 1190 1034
rect 894 898 950 954
rect 974 898 1030 954
rect 1054 898 1110 954
rect 1134 898 1190 954
rect 1598 1138 1654 1194
rect 1678 1138 1734 1194
rect 1758 1138 1814 1194
rect 1838 1138 1894 1194
rect 1598 1058 1654 1114
rect 1678 1058 1734 1114
rect 1758 1058 1814 1114
rect 1838 1058 1894 1114
rect 1598 978 1654 1034
rect 1678 978 1734 1034
rect 1758 978 1814 1034
rect 1838 978 1894 1034
rect 1598 898 1654 954
rect 1678 898 1734 954
rect 1758 898 1814 954
rect 1838 898 1894 954
rect 894 480 950 536
rect 974 480 1030 536
rect 1054 480 1110 536
rect 1134 480 1190 536
rect 894 400 950 456
rect 974 400 1030 456
rect 1054 400 1110 456
rect 1134 400 1190 456
rect 894 320 950 376
rect 974 320 1030 376
rect 1054 320 1110 376
rect 1134 320 1190 376
rect 894 240 950 296
rect 974 240 1030 296
rect 1054 240 1110 296
rect 1134 240 1190 296
rect 1598 480 1654 536
rect 1678 480 1734 536
rect 1758 480 1814 536
rect 1838 480 1894 536
rect 1598 400 1654 456
rect 1678 400 1734 456
rect 1758 400 1814 456
rect 1838 400 1894 456
rect 1598 320 1654 376
rect 1678 320 1734 376
rect 1758 320 1814 376
rect 1838 320 1894 376
rect 1598 240 1654 296
rect 1678 240 1734 296
rect 1758 240 1814 296
rect 1838 240 1894 296
rect 878 128 890 154
rect 890 128 934 154
rect 968 128 976 154
rect 976 128 1024 154
rect 1058 128 1106 154
rect 1106 128 1114 154
rect 1150 128 1188 154
rect 1188 128 1206 154
rect 878 98 934 128
rect 968 98 1024 128
rect 1058 98 1114 128
rect 1150 98 1206 128
rect 1582 128 1594 154
rect 1594 128 1638 154
rect 1672 128 1680 154
rect 1680 128 1728 154
rect 1762 128 1810 154
rect 1810 128 1818 154
rect 1854 128 1892 154
rect 1892 128 1910 154
rect 1582 98 1638 128
rect 1672 98 1728 128
rect 1762 98 1818 128
rect 1854 98 1910 128
rect 854 -132 914 -130
rect 854 -188 856 -132
rect 856 -188 912 -132
rect 912 -188 914 -132
rect 854 -190 914 -188
rect 980 -132 1040 -130
rect 980 -188 982 -132
rect 982 -188 1038 -132
rect 1038 -188 1040 -132
rect 980 -190 1040 -188
rect 854 -236 914 -234
rect 854 -292 856 -236
rect 856 -292 912 -236
rect 912 -292 914 -236
rect 854 -294 914 -292
rect 980 -236 1040 -234
rect 980 -292 982 -236
rect 982 -292 1038 -236
rect 1038 -292 1040 -236
rect 980 -294 1040 -292
rect 854 -320 914 -318
rect 854 -376 856 -320
rect 856 -376 912 -320
rect 912 -376 914 -320
rect 854 -378 914 -376
rect 980 -320 1040 -318
rect 980 -376 982 -320
rect 982 -376 1038 -320
rect 1038 -376 1040 -320
rect 980 -378 1040 -376
rect 854 -406 914 -404
rect 854 -462 856 -406
rect 856 -462 912 -406
rect 912 -462 914 -406
rect 854 -464 914 -462
rect 980 -406 1040 -404
rect 980 -462 982 -406
rect 982 -462 1038 -406
rect 1038 -462 1040 -406
rect 980 -464 1040 -462
rect 854 -500 914 -498
rect 854 -556 856 -500
rect 856 -556 912 -500
rect 912 -556 914 -500
rect 854 -558 914 -556
rect 980 -500 1040 -498
rect 980 -556 982 -500
rect 982 -556 1038 -500
rect 1038 -556 1040 -500
rect 980 -558 1040 -556
rect 854 -600 914 -598
rect 854 -656 856 -600
rect 856 -656 912 -600
rect 912 -656 914 -600
rect 854 -658 914 -656
rect 980 -600 1040 -598
rect 980 -656 982 -600
rect 982 -656 1038 -600
rect 1038 -656 1040 -600
rect 980 -658 1040 -656
rect 854 -684 914 -682
rect 854 -740 856 -684
rect 856 -740 912 -684
rect 912 -740 914 -684
rect 854 -742 914 -740
rect 980 -684 1040 -682
rect 980 -740 982 -684
rect 982 -740 1038 -684
rect 1038 -740 1040 -684
rect 980 -742 1040 -740
rect 1704 -132 1764 -130
rect 1704 -188 1706 -132
rect 1706 -188 1762 -132
rect 1762 -188 1764 -132
rect 1704 -190 1764 -188
rect 1830 -132 1890 -130
rect 1830 -188 1832 -132
rect 1832 -188 1888 -132
rect 1888 -188 1890 -132
rect 1830 -190 1890 -188
rect 1704 -236 1764 -234
rect 1704 -292 1706 -236
rect 1706 -292 1762 -236
rect 1762 -292 1764 -236
rect 1704 -294 1764 -292
rect 1830 -236 1890 -234
rect 1830 -292 1832 -236
rect 1832 -292 1888 -236
rect 1888 -292 1890 -236
rect 1830 -294 1890 -292
rect 1704 -320 1764 -318
rect 1704 -376 1706 -320
rect 1706 -376 1762 -320
rect 1762 -376 1764 -320
rect 1704 -378 1764 -376
rect 1830 -320 1890 -318
rect 1830 -376 1832 -320
rect 1832 -376 1888 -320
rect 1888 -376 1890 -320
rect 1830 -378 1890 -376
rect 1704 -406 1764 -404
rect 1704 -462 1706 -406
rect 1706 -462 1762 -406
rect 1762 -462 1764 -406
rect 1704 -464 1764 -462
rect 1830 -406 1890 -404
rect 1830 -462 1832 -406
rect 1832 -462 1888 -406
rect 1888 -462 1890 -406
rect 1830 -464 1890 -462
rect 1704 -500 1764 -498
rect 1704 -556 1706 -500
rect 1706 -556 1762 -500
rect 1762 -556 1764 -500
rect 1704 -558 1764 -556
rect 1830 -500 1890 -498
rect 1830 -556 1832 -500
rect 1832 -556 1888 -500
rect 1888 -556 1890 -500
rect 1830 -558 1890 -556
rect 1704 -600 1764 -598
rect 1704 -656 1706 -600
rect 1706 -656 1762 -600
rect 1762 -656 1764 -600
rect 1704 -658 1764 -656
rect 1830 -600 1890 -598
rect 1830 -656 1832 -600
rect 1832 -656 1888 -600
rect 1888 -656 1890 -600
rect 1830 -658 1890 -656
rect 1704 -684 1764 -682
rect 1704 -740 1706 -684
rect 1706 -740 1762 -684
rect 1762 -740 1764 -684
rect 1704 -742 1764 -740
rect 1830 -684 1890 -682
rect 1830 -740 1832 -684
rect 1832 -740 1888 -684
rect 1888 -740 1890 -684
rect 1830 -742 1890 -740
rect 3006 1138 3062 1194
rect 3086 1138 3142 1194
rect 3166 1138 3222 1194
rect 3246 1138 3302 1194
rect 3006 1058 3062 1114
rect 3086 1058 3142 1114
rect 3166 1058 3222 1114
rect 3246 1058 3302 1114
rect 3006 978 3062 1034
rect 3086 978 3142 1034
rect 3166 978 3222 1034
rect 3246 978 3302 1034
rect 3006 898 3062 954
rect 3086 898 3142 954
rect 3166 898 3222 954
rect 3246 898 3302 954
rect 3710 1138 3766 1194
rect 3790 1138 3846 1194
rect 3870 1138 3926 1194
rect 3950 1138 4006 1194
rect 3710 1058 3766 1114
rect 3790 1058 3846 1114
rect 3870 1058 3926 1114
rect 3950 1058 4006 1114
rect 3710 978 3766 1034
rect 3790 978 3846 1034
rect 3870 978 3926 1034
rect 3950 978 4006 1034
rect 3710 898 3766 954
rect 3790 898 3846 954
rect 3870 898 3926 954
rect 3950 898 4006 954
rect 3006 480 3062 536
rect 3086 480 3142 536
rect 3166 480 3222 536
rect 3246 480 3302 536
rect 3006 400 3062 456
rect 3086 400 3142 456
rect 3166 400 3222 456
rect 3246 400 3302 456
rect 3006 320 3062 376
rect 3086 320 3142 376
rect 3166 320 3222 376
rect 3246 320 3302 376
rect 3006 240 3062 296
rect 3086 240 3142 296
rect 3166 240 3222 296
rect 3246 240 3302 296
rect 3710 480 3766 536
rect 3790 480 3846 536
rect 3870 480 3926 536
rect 3950 480 4006 536
rect 3710 400 3766 456
rect 3790 400 3846 456
rect 3870 400 3926 456
rect 3950 400 4006 456
rect 3710 320 3766 376
rect 3790 320 3846 376
rect 3870 320 3926 376
rect 3950 320 4006 376
rect 3710 240 3766 296
rect 3790 240 3846 296
rect 3870 240 3926 296
rect 3950 240 4006 296
rect 2990 128 3002 154
rect 3002 128 3046 154
rect 3080 128 3088 154
rect 3088 128 3136 154
rect 3170 128 3218 154
rect 3218 128 3226 154
rect 3262 128 3300 154
rect 3300 128 3318 154
rect 2990 98 3046 128
rect 3080 98 3136 128
rect 3170 98 3226 128
rect 3262 98 3318 128
rect 3694 128 3706 154
rect 3706 128 3750 154
rect 3784 128 3792 154
rect 3792 128 3840 154
rect 3874 128 3922 154
rect 3922 128 3930 154
rect 3966 128 4004 154
rect 4004 128 4022 154
rect 3694 98 3750 128
rect 3784 98 3840 128
rect 3874 98 3930 128
rect 3966 98 4022 128
rect 2374 -190 2434 -130
rect 2500 -190 2560 -130
rect 2374 -294 2434 -234
rect 2500 -294 2560 -234
rect 2374 -378 2434 -318
rect 2500 -378 2560 -318
rect 2374 -464 2434 -404
rect 2500 -464 2560 -404
rect 2374 -558 2434 -498
rect 2500 -558 2560 -498
rect 2374 -658 2434 -598
rect 2500 -658 2560 -598
rect 2374 -742 2434 -682
rect 2500 -742 2560 -682
rect 2888 -132 2948 -130
rect 2888 -188 2890 -132
rect 2890 -188 2946 -132
rect 2946 -188 2948 -132
rect 2888 -190 2948 -188
rect 3014 -132 3074 -130
rect 3014 -188 3016 -132
rect 3016 -188 3072 -132
rect 3072 -188 3074 -132
rect 3014 -190 3074 -188
rect 2888 -236 2948 -234
rect 2888 -292 2890 -236
rect 2890 -292 2946 -236
rect 2946 -292 2948 -236
rect 2888 -294 2948 -292
rect 3014 -236 3074 -234
rect 3014 -292 3016 -236
rect 3016 -292 3072 -236
rect 3072 -292 3074 -236
rect 3014 -294 3074 -292
rect 2888 -320 2948 -318
rect 2888 -376 2890 -320
rect 2890 -376 2946 -320
rect 2946 -376 2948 -320
rect 2888 -378 2948 -376
rect 3014 -320 3074 -318
rect 3014 -376 3016 -320
rect 3016 -376 3072 -320
rect 3072 -376 3074 -320
rect 3014 -378 3074 -376
rect 2888 -406 2948 -404
rect 2888 -462 2890 -406
rect 2890 -462 2946 -406
rect 2946 -462 2948 -406
rect 2888 -464 2948 -462
rect 3014 -406 3074 -404
rect 3014 -462 3016 -406
rect 3016 -462 3072 -406
rect 3072 -462 3074 -406
rect 3014 -464 3074 -462
rect 2888 -500 2948 -498
rect 2888 -556 2890 -500
rect 2890 -556 2946 -500
rect 2946 -556 2948 -500
rect 2888 -558 2948 -556
rect 3014 -500 3074 -498
rect 3014 -556 3016 -500
rect 3016 -556 3072 -500
rect 3072 -556 3074 -500
rect 3014 -558 3074 -556
rect 2888 -600 2948 -598
rect 2888 -656 2890 -600
rect 2890 -656 2946 -600
rect 2946 -656 2948 -600
rect 2888 -658 2948 -656
rect 3014 -600 3074 -598
rect 3014 -656 3016 -600
rect 3016 -656 3072 -600
rect 3072 -656 3074 -600
rect 3014 -658 3074 -656
rect 2888 -684 2948 -682
rect 2888 -740 2890 -684
rect 2890 -740 2946 -684
rect 2946 -740 2948 -684
rect 2888 -742 2948 -740
rect 3014 -684 3074 -682
rect 3014 -740 3016 -684
rect 3016 -740 3072 -684
rect 3072 -740 3074 -684
rect 3014 -742 3074 -740
rect 3708 -132 3768 -130
rect 3708 -188 3710 -132
rect 3710 -188 3766 -132
rect 3766 -188 3768 -132
rect 3708 -190 3768 -188
rect 3834 -132 3894 -130
rect 3834 -188 3836 -132
rect 3836 -188 3892 -132
rect 3892 -188 3894 -132
rect 3834 -190 3894 -188
rect 3708 -236 3768 -234
rect 3708 -292 3710 -236
rect 3710 -292 3766 -236
rect 3766 -292 3768 -236
rect 3708 -294 3768 -292
rect 3834 -236 3894 -234
rect 3834 -292 3836 -236
rect 3836 -292 3892 -236
rect 3892 -292 3894 -236
rect 3834 -294 3894 -292
rect 3708 -320 3768 -318
rect 3708 -376 3710 -320
rect 3710 -376 3766 -320
rect 3766 -376 3768 -320
rect 3708 -378 3768 -376
rect 3834 -320 3894 -318
rect 3834 -376 3836 -320
rect 3836 -376 3892 -320
rect 3892 -376 3894 -320
rect 3834 -378 3894 -376
rect 3708 -406 3768 -404
rect 3708 -462 3710 -406
rect 3710 -462 3766 -406
rect 3766 -462 3768 -406
rect 3708 -464 3768 -462
rect 3834 -406 3894 -404
rect 3834 -462 3836 -406
rect 3836 -462 3892 -406
rect 3892 -462 3894 -406
rect 3834 -464 3894 -462
rect 3708 -500 3768 -498
rect 3708 -556 3710 -500
rect 3710 -556 3766 -500
rect 3766 -556 3768 -500
rect 3708 -558 3768 -556
rect 3834 -500 3894 -498
rect 3834 -556 3836 -500
rect 3836 -556 3892 -500
rect 3892 -556 3894 -500
rect 3834 -558 3894 -556
rect 3708 -600 3768 -598
rect 3708 -656 3710 -600
rect 3710 -656 3766 -600
rect 3766 -656 3768 -600
rect 3708 -658 3768 -656
rect 3834 -600 3894 -598
rect 3834 -656 3836 -600
rect 3836 -656 3892 -600
rect 3892 -656 3894 -600
rect 3834 -658 3894 -656
rect 3708 -684 3768 -682
rect 3708 -740 3710 -684
rect 3710 -740 3766 -684
rect 3766 -740 3768 -684
rect 3708 -742 3768 -740
rect 3834 -684 3894 -682
rect 3834 -740 3836 -684
rect 3836 -740 3892 -684
rect 3892 -740 3894 -684
rect 3834 -742 3894 -740
<< metal3 >>
rect 658 2736 738 2744
rect 658 2672 666 2736
rect 730 2672 738 2736
rect 658 2664 738 2672
rect 866 2664 1214 2666
rect 1570 2664 1918 2666
rect 2276 2664 2624 2666
rect 2980 2664 3328 2666
rect 3684 2664 4032 2666
rect 658 2660 4032 2664
rect 658 2656 876 2660
rect 658 2592 666 2656
rect 730 2604 876 2656
rect 932 2604 966 2660
rect 1022 2604 1056 2660
rect 1112 2604 1148 2660
rect 1204 2604 1580 2660
rect 1636 2604 1670 2660
rect 1726 2604 1760 2660
rect 1816 2604 1852 2660
rect 1908 2604 2286 2660
rect 2342 2604 2376 2660
rect 2432 2604 2466 2660
rect 2522 2604 2558 2660
rect 2614 2604 2990 2660
rect 3046 2604 3080 2660
rect 3136 2604 3170 2660
rect 3226 2604 3262 2660
rect 3318 2604 3694 2660
rect 3750 2604 3784 2660
rect 3840 2604 3874 2660
rect 3930 2604 3966 2660
rect 4022 2604 4032 2660
rect 730 2598 4032 2604
rect 730 2592 738 2598
rect 658 2584 738 2592
rect 842 2522 1242 2538
rect 842 2458 890 2522
rect 954 2458 970 2522
rect 1034 2458 1050 2522
rect 1114 2458 1130 2522
rect 1194 2458 1242 2522
rect 842 2442 1242 2458
rect 842 2378 890 2442
rect 954 2378 970 2442
rect 1034 2378 1050 2442
rect 1114 2378 1130 2442
rect 1194 2378 1242 2442
rect 842 2362 1242 2378
rect 842 2298 890 2362
rect 954 2298 970 2362
rect 1034 2298 1050 2362
rect 1114 2298 1130 2362
rect 1194 2298 1242 2362
rect 842 2282 1242 2298
rect 842 2218 890 2282
rect 954 2218 970 2282
rect 1034 2218 1050 2282
rect 1114 2218 1130 2282
rect 1194 2218 1242 2282
rect 842 2202 1242 2218
rect 1546 2522 1946 2538
rect 1546 2458 1594 2522
rect 1658 2458 1674 2522
rect 1738 2458 1754 2522
rect 1818 2458 1834 2522
rect 1898 2458 1946 2522
rect 1546 2442 1946 2458
rect 1546 2378 1594 2442
rect 1658 2378 1674 2442
rect 1738 2378 1754 2442
rect 1818 2378 1834 2442
rect 1898 2378 1946 2442
rect 1546 2362 1946 2378
rect 1546 2298 1594 2362
rect 1658 2298 1674 2362
rect 1738 2298 1754 2362
rect 1818 2298 1834 2362
rect 1898 2298 1946 2362
rect 1546 2282 1946 2298
rect 1546 2218 1594 2282
rect 1658 2218 1674 2282
rect 1738 2218 1754 2282
rect 1818 2218 1834 2282
rect 1898 2218 1946 2282
rect 1546 2202 1946 2218
rect 2250 2522 2650 2538
rect 2250 2458 2298 2522
rect 2362 2458 2378 2522
rect 2442 2458 2458 2522
rect 2522 2458 2538 2522
rect 2602 2458 2650 2522
rect 2250 2442 2650 2458
rect 2250 2378 2298 2442
rect 2362 2378 2378 2442
rect 2442 2378 2458 2442
rect 2522 2378 2538 2442
rect 2602 2378 2650 2442
rect 2250 2362 2650 2378
rect 2250 2298 2298 2362
rect 2362 2298 2378 2362
rect 2442 2298 2458 2362
rect 2522 2298 2538 2362
rect 2602 2298 2650 2362
rect 2250 2282 2650 2298
rect 2250 2218 2298 2282
rect 2362 2218 2378 2282
rect 2442 2218 2458 2282
rect 2522 2218 2538 2282
rect 2602 2218 2650 2282
rect 2250 2202 2650 2218
rect 2954 2522 3354 2538
rect 2954 2458 3002 2522
rect 3066 2458 3082 2522
rect 3146 2458 3162 2522
rect 3226 2458 3242 2522
rect 3306 2458 3354 2522
rect 2954 2442 3354 2458
rect 2954 2378 3002 2442
rect 3066 2378 3082 2442
rect 3146 2378 3162 2442
rect 3226 2378 3242 2442
rect 3306 2378 3354 2442
rect 2954 2362 3354 2378
rect 2954 2298 3002 2362
rect 3066 2298 3082 2362
rect 3146 2298 3162 2362
rect 3226 2298 3242 2362
rect 3306 2298 3354 2362
rect 2954 2282 3354 2298
rect 2954 2218 3002 2282
rect 3066 2218 3082 2282
rect 3146 2218 3162 2282
rect 3226 2218 3242 2282
rect 3306 2218 3354 2282
rect 2954 2202 3354 2218
rect 3658 2522 4058 2538
rect 3658 2458 3706 2522
rect 3770 2458 3786 2522
rect 3850 2458 3866 2522
rect 3930 2458 3946 2522
rect 4010 2458 4058 2522
rect 3658 2442 4058 2458
rect 3658 2378 3706 2442
rect 3770 2378 3786 2442
rect 3850 2378 3866 2442
rect 3930 2378 3946 2442
rect 4010 2378 4058 2442
rect 3658 2362 4058 2378
rect 3658 2298 3706 2362
rect 3770 2298 3786 2362
rect 3850 2298 3866 2362
rect 3930 2298 3946 2362
rect 4010 2298 4058 2362
rect 3658 2282 4058 2298
rect 3658 2218 3706 2282
rect 3770 2218 3786 2282
rect 3850 2218 3866 2282
rect 3930 2218 3946 2282
rect 4010 2218 4058 2282
rect 3658 2202 4058 2218
rect 844 1878 1244 1880
rect 842 1862 1244 1878
rect 842 1798 890 1862
rect 954 1798 970 1862
rect 1034 1798 1050 1862
rect 1114 1798 1130 1862
rect 1194 1798 1244 1862
rect 842 1782 1244 1798
rect 842 1718 890 1782
rect 954 1718 970 1782
rect 1034 1718 1050 1782
rect 1114 1718 1130 1782
rect 1194 1718 1244 1782
rect 842 1702 1244 1718
rect 842 1638 890 1702
rect 954 1638 970 1702
rect 1034 1638 1050 1702
rect 1114 1638 1130 1702
rect 1194 1638 1244 1702
rect 842 1622 1244 1638
rect 658 1572 738 1580
rect 658 1508 666 1572
rect 730 1508 738 1572
rect 842 1558 890 1622
rect 954 1558 970 1622
rect 1034 1558 1050 1622
rect 1114 1558 1130 1622
rect 1194 1558 1244 1622
rect 842 1544 1244 1558
rect 1546 1862 1948 1878
rect 1546 1798 1594 1862
rect 1658 1798 1674 1862
rect 1738 1798 1754 1862
rect 1818 1798 1834 1862
rect 1898 1798 1948 1862
rect 1546 1782 1948 1798
rect 1546 1718 1594 1782
rect 1658 1718 1674 1782
rect 1738 1718 1754 1782
rect 1818 1718 1834 1782
rect 1898 1718 1948 1782
rect 1546 1702 1948 1718
rect 1546 1638 1594 1702
rect 1658 1638 1674 1702
rect 1738 1638 1754 1702
rect 1818 1638 1834 1702
rect 1898 1638 1948 1702
rect 1546 1622 1948 1638
rect 1546 1558 1594 1622
rect 1658 1558 1674 1622
rect 1738 1558 1754 1622
rect 1818 1558 1834 1622
rect 1898 1558 1948 1622
rect 842 1542 1242 1544
rect 1546 1542 1948 1558
rect 2250 1862 2652 1878
rect 2250 1798 2298 1862
rect 2362 1798 2378 1862
rect 2442 1798 2458 1862
rect 2522 1798 2538 1862
rect 2602 1798 2652 1862
rect 2250 1782 2652 1798
rect 2250 1718 2298 1782
rect 2362 1718 2378 1782
rect 2442 1718 2458 1782
rect 2522 1718 2538 1782
rect 2602 1718 2652 1782
rect 2250 1702 2652 1718
rect 2250 1638 2298 1702
rect 2362 1638 2378 1702
rect 2442 1638 2458 1702
rect 2522 1638 2538 1702
rect 2602 1638 2652 1702
rect 2250 1622 2652 1638
rect 2250 1558 2298 1622
rect 2362 1558 2378 1622
rect 2442 1558 2458 1622
rect 2522 1558 2538 1622
rect 2602 1558 2652 1622
rect 2250 1542 2652 1558
rect 2954 1862 3356 1878
rect 2954 1798 3002 1862
rect 3066 1798 3082 1862
rect 3146 1798 3162 1862
rect 3226 1798 3242 1862
rect 3306 1798 3356 1862
rect 2954 1782 3356 1798
rect 2954 1718 3002 1782
rect 3066 1718 3082 1782
rect 3146 1718 3162 1782
rect 3226 1718 3242 1782
rect 3306 1718 3356 1782
rect 2954 1702 3356 1718
rect 2954 1638 3002 1702
rect 3066 1638 3082 1702
rect 3146 1638 3162 1702
rect 3226 1638 3242 1702
rect 3306 1638 3356 1702
rect 2954 1622 3356 1638
rect 2954 1558 3002 1622
rect 3066 1558 3082 1622
rect 3146 1558 3162 1622
rect 3226 1558 3242 1622
rect 3306 1558 3356 1622
rect 2954 1542 3356 1558
rect 3658 1862 4060 1878
rect 3658 1798 3706 1862
rect 3770 1798 3786 1862
rect 3850 1798 3866 1862
rect 3930 1798 3946 1862
rect 4010 1798 4060 1862
rect 3658 1782 4060 1798
rect 3658 1718 3706 1782
rect 3770 1718 3786 1782
rect 3850 1718 3866 1782
rect 3930 1718 3946 1782
rect 4010 1718 4060 1782
rect 3658 1702 4060 1718
rect 3658 1638 3706 1702
rect 3770 1638 3786 1702
rect 3850 1638 3866 1702
rect 3930 1638 3946 1702
rect 4010 1638 4060 1702
rect 3658 1622 4060 1638
rect 3658 1558 3706 1622
rect 3770 1558 3786 1622
rect 3850 1558 3866 1622
rect 3930 1558 3946 1622
rect 4010 1558 4060 1622
rect 3658 1542 4060 1558
rect 658 1492 738 1508
rect 658 1428 666 1492
rect 730 1482 738 1492
rect 730 1476 4032 1482
rect 730 1428 878 1476
rect 658 1420 878 1428
rect 934 1420 968 1476
rect 1024 1420 1058 1476
rect 1114 1420 1150 1476
rect 1206 1420 1582 1476
rect 1638 1420 1672 1476
rect 1728 1420 1762 1476
rect 1818 1420 1854 1476
rect 1910 1420 2286 1476
rect 2342 1420 2376 1476
rect 2432 1420 2466 1476
rect 2522 1420 2558 1476
rect 2614 1420 2990 1476
rect 3046 1420 3080 1476
rect 3136 1420 3170 1476
rect 3226 1420 3262 1476
rect 3318 1420 3694 1476
rect 3750 1420 3784 1476
rect 3840 1420 3874 1476
rect 3930 1420 3966 1476
rect 4022 1420 4032 1476
rect 868 1414 1216 1420
rect 1572 1414 1920 1420
rect 2276 1414 2624 1420
rect 2980 1414 3328 1420
rect 3684 1414 4032 1420
rect 868 1340 1216 1342
rect 1572 1340 1920 1342
rect 2980 1340 3328 1342
rect 3684 1340 4032 1342
rect 658 1336 4032 1340
rect 658 1332 878 1336
rect 658 1268 666 1332
rect 730 1280 878 1332
rect 934 1280 968 1336
rect 1024 1280 1058 1336
rect 1114 1280 1150 1336
rect 1206 1280 1582 1336
rect 1638 1280 1672 1336
rect 1728 1280 1762 1336
rect 1818 1280 1854 1336
rect 1910 1280 2990 1336
rect 3046 1280 3080 1336
rect 3136 1280 3170 1336
rect 3226 1280 3262 1336
rect 3318 1280 3694 1336
rect 3750 1280 3784 1336
rect 3840 1280 3874 1336
rect 3930 1280 3966 1336
rect 4022 1280 4032 1336
rect 730 1274 4032 1280
rect 730 1268 738 1274
rect 658 1252 738 1268
rect 658 1188 666 1252
rect 730 1188 738 1252
rect 658 1182 738 1188
rect 842 1198 1242 1214
rect 842 1134 890 1198
rect 954 1134 970 1198
rect 1034 1134 1050 1198
rect 1114 1134 1130 1198
rect 1194 1134 1242 1198
rect 842 1118 1242 1134
rect 842 1054 890 1118
rect 954 1054 970 1118
rect 1034 1054 1050 1118
rect 1114 1054 1130 1118
rect 1194 1054 1242 1118
rect 842 1038 1242 1054
rect 842 974 890 1038
rect 954 974 970 1038
rect 1034 974 1050 1038
rect 1114 974 1130 1038
rect 1194 974 1242 1038
rect 842 958 1242 974
rect 842 894 890 958
rect 954 894 970 958
rect 1034 894 1050 958
rect 1114 894 1130 958
rect 1194 894 1242 958
rect 842 878 1242 894
rect 1546 1198 1946 1214
rect 1546 1134 1594 1198
rect 1658 1134 1674 1198
rect 1738 1134 1754 1198
rect 1818 1134 1834 1198
rect 1898 1134 1946 1198
rect 1546 1118 1946 1134
rect 1546 1054 1594 1118
rect 1658 1054 1674 1118
rect 1738 1054 1754 1118
rect 1818 1054 1834 1118
rect 1898 1054 1946 1118
rect 1546 1038 1946 1054
rect 1546 974 1594 1038
rect 1658 974 1674 1038
rect 1738 974 1754 1038
rect 1818 974 1834 1038
rect 1898 974 1946 1038
rect 1546 958 1946 974
rect 1546 894 1594 958
rect 1658 894 1674 958
rect 1738 894 1754 958
rect 1818 894 1834 958
rect 1898 894 1946 958
rect 1546 878 1946 894
rect 2954 1198 3354 1214
rect 2954 1134 3002 1198
rect 3066 1134 3082 1198
rect 3146 1134 3162 1198
rect 3226 1134 3242 1198
rect 3306 1134 3354 1198
rect 2954 1118 3354 1134
rect 2954 1054 3002 1118
rect 3066 1054 3082 1118
rect 3146 1054 3162 1118
rect 3226 1054 3242 1118
rect 3306 1054 3354 1118
rect 2954 1038 3354 1054
rect 2954 974 3002 1038
rect 3066 974 3082 1038
rect 3146 974 3162 1038
rect 3226 974 3242 1038
rect 3306 974 3354 1038
rect 2954 958 3354 974
rect 2954 894 3002 958
rect 3066 894 3082 958
rect 3146 894 3162 958
rect 3226 894 3242 958
rect 3306 894 3354 958
rect 2954 878 3354 894
rect 3658 1198 4058 1214
rect 3658 1134 3706 1198
rect 3770 1134 3786 1198
rect 3850 1134 3866 1198
rect 3930 1134 3946 1198
rect 4010 1134 4058 1198
rect 3658 1118 4058 1134
rect 3658 1054 3706 1118
rect 3770 1054 3786 1118
rect 3850 1054 3866 1118
rect 3930 1054 3946 1118
rect 4010 1054 4058 1118
rect 3658 1038 4058 1054
rect 3658 974 3706 1038
rect 3770 974 3786 1038
rect 3850 974 3866 1038
rect 3930 974 3946 1038
rect 4010 974 4058 1038
rect 3658 958 4058 974
rect 3658 894 3706 958
rect 3770 894 3786 958
rect 3850 894 3866 958
rect 3930 894 3946 958
rect 4010 894 4058 958
rect 3658 878 4058 894
rect 842 540 1244 556
rect 842 476 890 540
rect 954 476 970 540
rect 1034 476 1050 540
rect 1114 476 1130 540
rect 1194 476 1244 540
rect 842 460 1244 476
rect 842 396 890 460
rect 954 396 970 460
rect 1034 396 1050 460
rect 1114 396 1130 460
rect 1194 396 1244 460
rect 842 380 1244 396
rect 842 316 890 380
rect 954 316 970 380
rect 1034 316 1050 380
rect 1114 316 1130 380
rect 1194 316 1244 380
rect 842 300 1244 316
rect 658 246 738 254
rect 658 182 666 246
rect 730 182 738 246
rect 842 236 890 300
rect 954 236 970 300
rect 1034 236 1050 300
rect 1114 236 1130 300
rect 1194 236 1244 300
rect 842 220 1244 236
rect 1546 540 1948 556
rect 1546 476 1594 540
rect 1658 476 1674 540
rect 1738 476 1754 540
rect 1818 476 1834 540
rect 1898 476 1948 540
rect 1546 460 1948 476
rect 1546 396 1594 460
rect 1658 396 1674 460
rect 1738 396 1754 460
rect 1818 396 1834 460
rect 1898 396 1948 460
rect 1546 380 1948 396
rect 1546 316 1594 380
rect 1658 316 1674 380
rect 1738 316 1754 380
rect 1818 316 1834 380
rect 1898 316 1948 380
rect 1546 300 1948 316
rect 1546 236 1594 300
rect 1658 236 1674 300
rect 1738 236 1754 300
rect 1818 236 1834 300
rect 1898 236 1948 300
rect 1546 220 1948 236
rect 2954 540 3356 556
rect 2954 476 3002 540
rect 3066 476 3082 540
rect 3146 476 3162 540
rect 3226 476 3242 540
rect 3306 476 3356 540
rect 2954 460 3356 476
rect 2954 396 3002 460
rect 3066 396 3082 460
rect 3146 396 3162 460
rect 3226 396 3242 460
rect 3306 396 3356 460
rect 2954 380 3356 396
rect 2954 316 3002 380
rect 3066 316 3082 380
rect 3146 316 3162 380
rect 3226 316 3242 380
rect 3306 316 3356 380
rect 2954 300 3356 316
rect 2954 236 3002 300
rect 3066 236 3082 300
rect 3146 236 3162 300
rect 3226 236 3242 300
rect 3306 236 3356 300
rect 2954 220 3356 236
rect 3604 540 4058 556
rect 3604 476 3706 540
rect 3770 476 3786 540
rect 3850 476 3866 540
rect 3930 476 3946 540
rect 4010 476 4058 540
rect 3604 460 4058 476
rect 3604 396 3706 460
rect 3770 396 3786 460
rect 3850 396 3866 460
rect 3930 396 3946 460
rect 4010 396 4058 460
rect 3604 380 4058 396
rect 3604 316 3706 380
rect 3770 316 3786 380
rect 3850 316 3866 380
rect 3930 316 3946 380
rect 4010 316 4058 380
rect 3604 300 4058 316
rect 3604 236 3706 300
rect 3770 236 3786 300
rect 3850 236 3866 300
rect 3930 236 3946 300
rect 4010 236 4058 300
rect 3604 220 4058 236
rect 658 166 738 182
rect 658 102 666 166
rect 730 160 738 166
rect 730 154 4032 160
rect 730 102 878 154
rect 658 98 878 102
rect 934 98 968 154
rect 1024 98 1058 154
rect 1114 98 1150 154
rect 1206 98 1582 154
rect 1638 98 1672 154
rect 1728 98 1762 154
rect 1818 98 1854 154
rect 1910 98 2990 154
rect 3046 98 3080 154
rect 3136 98 3170 154
rect 3226 98 3262 154
rect 3318 98 3694 154
rect 3750 98 3784 154
rect 3840 98 3874 154
rect 3930 98 3966 154
rect 4022 98 4032 154
rect 658 94 4032 98
rect 868 92 1216 94
rect 1572 92 1920 94
rect 2980 92 3328 94
rect 3684 92 4032 94
rect 226 -128 450 -100
rect 226 -192 244 -128
rect 308 -192 370 -128
rect 434 -192 450 -128
rect 226 -232 450 -192
rect 226 -296 244 -232
rect 308 -296 370 -232
rect 434 -296 450 -232
rect 226 -316 450 -296
rect 226 -380 244 -316
rect 308 -380 370 -316
rect 434 -380 450 -316
rect 226 -402 450 -380
rect 226 -466 244 -402
rect 308 -466 370 -402
rect 434 -466 450 -402
rect 226 -496 450 -466
rect 226 -560 244 -496
rect 308 -560 370 -496
rect 434 -560 450 -496
rect 226 -596 450 -560
rect 226 -660 244 -596
rect 308 -660 370 -596
rect 434 -660 450 -596
rect 226 -680 450 -660
rect 226 -744 244 -680
rect 308 -744 370 -680
rect 434 -744 450 -680
rect 226 -772 450 -744
rect 834 -128 1058 -100
rect 834 -192 852 -128
rect 916 -192 978 -128
rect 1042 -192 1058 -128
rect 834 -232 1058 -192
rect 834 -296 852 -232
rect 916 -296 978 -232
rect 1042 -296 1058 -232
rect 834 -316 1058 -296
rect 834 -380 852 -316
rect 916 -380 978 -316
rect 1042 -380 1058 -316
rect 834 -402 1058 -380
rect 834 -466 852 -402
rect 916 -466 978 -402
rect 1042 -466 1058 -402
rect 834 -496 1058 -466
rect 834 -560 852 -496
rect 916 -560 978 -496
rect 1042 -560 1058 -496
rect 834 -596 1058 -560
rect 834 -660 852 -596
rect 916 -660 978 -596
rect 1042 -660 1058 -596
rect 834 -680 1058 -660
rect 834 -744 852 -680
rect 916 -744 978 -680
rect 1042 -744 1058 -680
rect 834 -772 1058 -744
rect 1684 -128 1908 -100
rect 1684 -192 1702 -128
rect 1766 -192 1828 -128
rect 1892 -192 1908 -128
rect 1684 -232 1908 -192
rect 1684 -296 1702 -232
rect 1766 -296 1828 -232
rect 1892 -296 1908 -232
rect 1684 -316 1908 -296
rect 1684 -380 1702 -316
rect 1766 -380 1828 -316
rect 1892 -380 1908 -316
rect 1684 -402 1908 -380
rect 1684 -466 1702 -402
rect 1766 -466 1828 -402
rect 1892 -466 1908 -402
rect 1684 -496 1908 -466
rect 1684 -560 1702 -496
rect 1766 -560 1828 -496
rect 1892 -560 1908 -496
rect 1684 -596 1908 -560
rect 1684 -660 1702 -596
rect 1766 -660 1828 -596
rect 1892 -660 1908 -596
rect 1684 -680 1908 -660
rect 1684 -744 1702 -680
rect 1766 -744 1828 -680
rect 1892 -744 1908 -680
rect 1684 -772 1908 -744
rect 2354 -128 2578 -100
rect 2354 -192 2372 -128
rect 2436 -192 2498 -128
rect 2562 -192 2578 -128
rect 2354 -232 2578 -192
rect 2354 -296 2372 -232
rect 2436 -296 2498 -232
rect 2562 -296 2578 -232
rect 2354 -316 2578 -296
rect 2354 -380 2372 -316
rect 2436 -380 2498 -316
rect 2562 -380 2578 -316
rect 2354 -402 2578 -380
rect 2354 -466 2372 -402
rect 2436 -466 2498 -402
rect 2562 -466 2578 -402
rect 2354 -496 2578 -466
rect 2354 -560 2372 -496
rect 2436 -560 2498 -496
rect 2562 -560 2578 -496
rect 2354 -596 2578 -560
rect 2354 -660 2372 -596
rect 2436 -660 2498 -596
rect 2562 -660 2578 -596
rect 2354 -680 2578 -660
rect 2354 -744 2372 -680
rect 2436 -744 2498 -680
rect 2562 -744 2578 -680
rect 2354 -772 2578 -744
rect 2868 -128 3092 -100
rect 2868 -192 2886 -128
rect 2950 -192 3012 -128
rect 3076 -192 3092 -128
rect 2868 -232 3092 -192
rect 2868 -296 2886 -232
rect 2950 -296 3012 -232
rect 3076 -296 3092 -232
rect 2868 -316 3092 -296
rect 2868 -380 2886 -316
rect 2950 -380 3012 -316
rect 3076 -380 3092 -316
rect 2868 -402 3092 -380
rect 2868 -466 2886 -402
rect 2950 -466 3012 -402
rect 3076 -466 3092 -402
rect 2868 -496 3092 -466
rect 2868 -560 2886 -496
rect 2950 -560 3012 -496
rect 3076 -560 3092 -496
rect 2868 -596 3092 -560
rect 2868 -660 2886 -596
rect 2950 -660 3012 -596
rect 3076 -660 3092 -596
rect 2868 -680 3092 -660
rect 2868 -744 2886 -680
rect 2950 -744 3012 -680
rect 3076 -744 3092 -680
rect 2868 -772 3092 -744
rect 3688 -128 3912 -100
rect 3688 -192 3706 -128
rect 3770 -192 3832 -128
rect 3896 -192 3912 -128
rect 3688 -232 3912 -192
rect 3688 -296 3706 -232
rect 3770 -296 3832 -232
rect 3896 -296 3912 -232
rect 3688 -316 3912 -296
rect 3688 -380 3706 -316
rect 3770 -380 3832 -316
rect 3896 -380 3912 -316
rect 3688 -402 3912 -380
rect 3688 -466 3706 -402
rect 3770 -466 3832 -402
rect 3896 -466 3912 -402
rect 3688 -496 3912 -466
rect 3688 -560 3706 -496
rect 3770 -560 3832 -496
rect 3896 -560 3912 -496
rect 3688 -596 3912 -560
rect 3688 -660 3706 -596
rect 3770 -660 3832 -596
rect 3896 -660 3912 -596
rect 3688 -680 3912 -660
rect 3688 -744 3706 -680
rect 3770 -744 3832 -680
rect 3896 -744 3912 -680
rect 3688 -772 3912 -744
rect 4446 -128 4670 -100
rect 4446 -192 4464 -128
rect 4528 -192 4590 -128
rect 4654 -192 4670 -128
rect 4446 -232 4670 -192
rect 4446 -296 4464 -232
rect 4528 -296 4590 -232
rect 4654 -296 4670 -232
rect 4446 -316 4670 -296
rect 4446 -380 4464 -316
rect 4528 -380 4590 -316
rect 4654 -380 4670 -316
rect 4446 -402 4670 -380
rect 4446 -466 4464 -402
rect 4528 -466 4590 -402
rect 4654 -466 4670 -402
rect 4446 -496 4670 -466
rect 4446 -560 4464 -496
rect 4528 -560 4590 -496
rect 4654 -560 4670 -496
rect 4446 -596 4670 -560
rect 4446 -660 4464 -596
rect 4528 -660 4590 -596
rect 4654 -660 4670 -596
rect 4446 -680 4670 -660
rect 4446 -744 4464 -680
rect 4528 -744 4590 -680
rect 4654 -744 4670 -680
rect 4446 -772 4670 -744
<< via3 >>
rect 666 2672 730 2736
rect 666 2592 730 2656
rect 890 2518 954 2522
rect 890 2462 894 2518
rect 894 2462 950 2518
rect 950 2462 954 2518
rect 890 2458 954 2462
rect 970 2518 1034 2522
rect 970 2462 974 2518
rect 974 2462 1030 2518
rect 1030 2462 1034 2518
rect 970 2458 1034 2462
rect 1050 2518 1114 2522
rect 1050 2462 1054 2518
rect 1054 2462 1110 2518
rect 1110 2462 1114 2518
rect 1050 2458 1114 2462
rect 1130 2518 1194 2522
rect 1130 2462 1134 2518
rect 1134 2462 1190 2518
rect 1190 2462 1194 2518
rect 1130 2458 1194 2462
rect 890 2438 954 2442
rect 890 2382 894 2438
rect 894 2382 950 2438
rect 950 2382 954 2438
rect 890 2378 954 2382
rect 970 2438 1034 2442
rect 970 2382 974 2438
rect 974 2382 1030 2438
rect 1030 2382 1034 2438
rect 970 2378 1034 2382
rect 1050 2438 1114 2442
rect 1050 2382 1054 2438
rect 1054 2382 1110 2438
rect 1110 2382 1114 2438
rect 1050 2378 1114 2382
rect 1130 2438 1194 2442
rect 1130 2382 1134 2438
rect 1134 2382 1190 2438
rect 1190 2382 1194 2438
rect 1130 2378 1194 2382
rect 890 2358 954 2362
rect 890 2302 894 2358
rect 894 2302 950 2358
rect 950 2302 954 2358
rect 890 2298 954 2302
rect 970 2358 1034 2362
rect 970 2302 974 2358
rect 974 2302 1030 2358
rect 1030 2302 1034 2358
rect 970 2298 1034 2302
rect 1050 2358 1114 2362
rect 1050 2302 1054 2358
rect 1054 2302 1110 2358
rect 1110 2302 1114 2358
rect 1050 2298 1114 2302
rect 1130 2358 1194 2362
rect 1130 2302 1134 2358
rect 1134 2302 1190 2358
rect 1190 2302 1194 2358
rect 1130 2298 1194 2302
rect 890 2278 954 2282
rect 890 2222 894 2278
rect 894 2222 950 2278
rect 950 2222 954 2278
rect 890 2218 954 2222
rect 970 2278 1034 2282
rect 970 2222 974 2278
rect 974 2222 1030 2278
rect 1030 2222 1034 2278
rect 970 2218 1034 2222
rect 1050 2278 1114 2282
rect 1050 2222 1054 2278
rect 1054 2222 1110 2278
rect 1110 2222 1114 2278
rect 1050 2218 1114 2222
rect 1130 2278 1194 2282
rect 1130 2222 1134 2278
rect 1134 2222 1190 2278
rect 1190 2222 1194 2278
rect 1130 2218 1194 2222
rect 1594 2518 1658 2522
rect 1594 2462 1598 2518
rect 1598 2462 1654 2518
rect 1654 2462 1658 2518
rect 1594 2458 1658 2462
rect 1674 2518 1738 2522
rect 1674 2462 1678 2518
rect 1678 2462 1734 2518
rect 1734 2462 1738 2518
rect 1674 2458 1738 2462
rect 1754 2518 1818 2522
rect 1754 2462 1758 2518
rect 1758 2462 1814 2518
rect 1814 2462 1818 2518
rect 1754 2458 1818 2462
rect 1834 2518 1898 2522
rect 1834 2462 1838 2518
rect 1838 2462 1894 2518
rect 1894 2462 1898 2518
rect 1834 2458 1898 2462
rect 1594 2438 1658 2442
rect 1594 2382 1598 2438
rect 1598 2382 1654 2438
rect 1654 2382 1658 2438
rect 1594 2378 1658 2382
rect 1674 2438 1738 2442
rect 1674 2382 1678 2438
rect 1678 2382 1734 2438
rect 1734 2382 1738 2438
rect 1674 2378 1738 2382
rect 1754 2438 1818 2442
rect 1754 2382 1758 2438
rect 1758 2382 1814 2438
rect 1814 2382 1818 2438
rect 1754 2378 1818 2382
rect 1834 2438 1898 2442
rect 1834 2382 1838 2438
rect 1838 2382 1894 2438
rect 1894 2382 1898 2438
rect 1834 2378 1898 2382
rect 1594 2358 1658 2362
rect 1594 2302 1598 2358
rect 1598 2302 1654 2358
rect 1654 2302 1658 2358
rect 1594 2298 1658 2302
rect 1674 2358 1738 2362
rect 1674 2302 1678 2358
rect 1678 2302 1734 2358
rect 1734 2302 1738 2358
rect 1674 2298 1738 2302
rect 1754 2358 1818 2362
rect 1754 2302 1758 2358
rect 1758 2302 1814 2358
rect 1814 2302 1818 2358
rect 1754 2298 1818 2302
rect 1834 2358 1898 2362
rect 1834 2302 1838 2358
rect 1838 2302 1894 2358
rect 1894 2302 1898 2358
rect 1834 2298 1898 2302
rect 1594 2278 1658 2282
rect 1594 2222 1598 2278
rect 1598 2222 1654 2278
rect 1654 2222 1658 2278
rect 1594 2218 1658 2222
rect 1674 2278 1738 2282
rect 1674 2222 1678 2278
rect 1678 2222 1734 2278
rect 1734 2222 1738 2278
rect 1674 2218 1738 2222
rect 1754 2278 1818 2282
rect 1754 2222 1758 2278
rect 1758 2222 1814 2278
rect 1814 2222 1818 2278
rect 1754 2218 1818 2222
rect 1834 2278 1898 2282
rect 1834 2222 1838 2278
rect 1838 2222 1894 2278
rect 1894 2222 1898 2278
rect 1834 2218 1898 2222
rect 2298 2518 2362 2522
rect 2298 2462 2302 2518
rect 2302 2462 2358 2518
rect 2358 2462 2362 2518
rect 2298 2458 2362 2462
rect 2378 2518 2442 2522
rect 2378 2462 2382 2518
rect 2382 2462 2438 2518
rect 2438 2462 2442 2518
rect 2378 2458 2442 2462
rect 2458 2518 2522 2522
rect 2458 2462 2462 2518
rect 2462 2462 2518 2518
rect 2518 2462 2522 2518
rect 2458 2458 2522 2462
rect 2538 2518 2602 2522
rect 2538 2462 2542 2518
rect 2542 2462 2598 2518
rect 2598 2462 2602 2518
rect 2538 2458 2602 2462
rect 2298 2438 2362 2442
rect 2298 2382 2302 2438
rect 2302 2382 2358 2438
rect 2358 2382 2362 2438
rect 2298 2378 2362 2382
rect 2378 2438 2442 2442
rect 2378 2382 2382 2438
rect 2382 2382 2438 2438
rect 2438 2382 2442 2438
rect 2378 2378 2442 2382
rect 2458 2438 2522 2442
rect 2458 2382 2462 2438
rect 2462 2382 2518 2438
rect 2518 2382 2522 2438
rect 2458 2378 2522 2382
rect 2538 2438 2602 2442
rect 2538 2382 2542 2438
rect 2542 2382 2598 2438
rect 2598 2382 2602 2438
rect 2538 2378 2602 2382
rect 2298 2358 2362 2362
rect 2298 2302 2302 2358
rect 2302 2302 2358 2358
rect 2358 2302 2362 2358
rect 2298 2298 2362 2302
rect 2378 2358 2442 2362
rect 2378 2302 2382 2358
rect 2382 2302 2438 2358
rect 2438 2302 2442 2358
rect 2378 2298 2442 2302
rect 2458 2358 2522 2362
rect 2458 2302 2462 2358
rect 2462 2302 2518 2358
rect 2518 2302 2522 2358
rect 2458 2298 2522 2302
rect 2538 2358 2602 2362
rect 2538 2302 2542 2358
rect 2542 2302 2598 2358
rect 2598 2302 2602 2358
rect 2538 2298 2602 2302
rect 2298 2278 2362 2282
rect 2298 2222 2302 2278
rect 2302 2222 2358 2278
rect 2358 2222 2362 2278
rect 2298 2218 2362 2222
rect 2378 2278 2442 2282
rect 2378 2222 2382 2278
rect 2382 2222 2438 2278
rect 2438 2222 2442 2278
rect 2378 2218 2442 2222
rect 2458 2278 2522 2282
rect 2458 2222 2462 2278
rect 2462 2222 2518 2278
rect 2518 2222 2522 2278
rect 2458 2218 2522 2222
rect 2538 2278 2602 2282
rect 2538 2222 2542 2278
rect 2542 2222 2598 2278
rect 2598 2222 2602 2278
rect 2538 2218 2602 2222
rect 3002 2518 3066 2522
rect 3002 2462 3006 2518
rect 3006 2462 3062 2518
rect 3062 2462 3066 2518
rect 3002 2458 3066 2462
rect 3082 2518 3146 2522
rect 3082 2462 3086 2518
rect 3086 2462 3142 2518
rect 3142 2462 3146 2518
rect 3082 2458 3146 2462
rect 3162 2518 3226 2522
rect 3162 2462 3166 2518
rect 3166 2462 3222 2518
rect 3222 2462 3226 2518
rect 3162 2458 3226 2462
rect 3242 2518 3306 2522
rect 3242 2462 3246 2518
rect 3246 2462 3302 2518
rect 3302 2462 3306 2518
rect 3242 2458 3306 2462
rect 3002 2438 3066 2442
rect 3002 2382 3006 2438
rect 3006 2382 3062 2438
rect 3062 2382 3066 2438
rect 3002 2378 3066 2382
rect 3082 2438 3146 2442
rect 3082 2382 3086 2438
rect 3086 2382 3142 2438
rect 3142 2382 3146 2438
rect 3082 2378 3146 2382
rect 3162 2438 3226 2442
rect 3162 2382 3166 2438
rect 3166 2382 3222 2438
rect 3222 2382 3226 2438
rect 3162 2378 3226 2382
rect 3242 2438 3306 2442
rect 3242 2382 3246 2438
rect 3246 2382 3302 2438
rect 3302 2382 3306 2438
rect 3242 2378 3306 2382
rect 3002 2358 3066 2362
rect 3002 2302 3006 2358
rect 3006 2302 3062 2358
rect 3062 2302 3066 2358
rect 3002 2298 3066 2302
rect 3082 2358 3146 2362
rect 3082 2302 3086 2358
rect 3086 2302 3142 2358
rect 3142 2302 3146 2358
rect 3082 2298 3146 2302
rect 3162 2358 3226 2362
rect 3162 2302 3166 2358
rect 3166 2302 3222 2358
rect 3222 2302 3226 2358
rect 3162 2298 3226 2302
rect 3242 2358 3306 2362
rect 3242 2302 3246 2358
rect 3246 2302 3302 2358
rect 3302 2302 3306 2358
rect 3242 2298 3306 2302
rect 3002 2278 3066 2282
rect 3002 2222 3006 2278
rect 3006 2222 3062 2278
rect 3062 2222 3066 2278
rect 3002 2218 3066 2222
rect 3082 2278 3146 2282
rect 3082 2222 3086 2278
rect 3086 2222 3142 2278
rect 3142 2222 3146 2278
rect 3082 2218 3146 2222
rect 3162 2278 3226 2282
rect 3162 2222 3166 2278
rect 3166 2222 3222 2278
rect 3222 2222 3226 2278
rect 3162 2218 3226 2222
rect 3242 2278 3306 2282
rect 3242 2222 3246 2278
rect 3246 2222 3302 2278
rect 3302 2222 3306 2278
rect 3242 2218 3306 2222
rect 3706 2518 3770 2522
rect 3706 2462 3710 2518
rect 3710 2462 3766 2518
rect 3766 2462 3770 2518
rect 3706 2458 3770 2462
rect 3786 2518 3850 2522
rect 3786 2462 3790 2518
rect 3790 2462 3846 2518
rect 3846 2462 3850 2518
rect 3786 2458 3850 2462
rect 3866 2518 3930 2522
rect 3866 2462 3870 2518
rect 3870 2462 3926 2518
rect 3926 2462 3930 2518
rect 3866 2458 3930 2462
rect 3946 2518 4010 2522
rect 3946 2462 3950 2518
rect 3950 2462 4006 2518
rect 4006 2462 4010 2518
rect 3946 2458 4010 2462
rect 3706 2438 3770 2442
rect 3706 2382 3710 2438
rect 3710 2382 3766 2438
rect 3766 2382 3770 2438
rect 3706 2378 3770 2382
rect 3786 2438 3850 2442
rect 3786 2382 3790 2438
rect 3790 2382 3846 2438
rect 3846 2382 3850 2438
rect 3786 2378 3850 2382
rect 3866 2438 3930 2442
rect 3866 2382 3870 2438
rect 3870 2382 3926 2438
rect 3926 2382 3930 2438
rect 3866 2378 3930 2382
rect 3946 2438 4010 2442
rect 3946 2382 3950 2438
rect 3950 2382 4006 2438
rect 4006 2382 4010 2438
rect 3946 2378 4010 2382
rect 3706 2358 3770 2362
rect 3706 2302 3710 2358
rect 3710 2302 3766 2358
rect 3766 2302 3770 2358
rect 3706 2298 3770 2302
rect 3786 2358 3850 2362
rect 3786 2302 3790 2358
rect 3790 2302 3846 2358
rect 3846 2302 3850 2358
rect 3786 2298 3850 2302
rect 3866 2358 3930 2362
rect 3866 2302 3870 2358
rect 3870 2302 3926 2358
rect 3926 2302 3930 2358
rect 3866 2298 3930 2302
rect 3946 2358 4010 2362
rect 3946 2302 3950 2358
rect 3950 2302 4006 2358
rect 4006 2302 4010 2358
rect 3946 2298 4010 2302
rect 3706 2278 3770 2282
rect 3706 2222 3710 2278
rect 3710 2222 3766 2278
rect 3766 2222 3770 2278
rect 3706 2218 3770 2222
rect 3786 2278 3850 2282
rect 3786 2222 3790 2278
rect 3790 2222 3846 2278
rect 3846 2222 3850 2278
rect 3786 2218 3850 2222
rect 3866 2278 3930 2282
rect 3866 2222 3870 2278
rect 3870 2222 3926 2278
rect 3926 2222 3930 2278
rect 3866 2218 3930 2222
rect 3946 2278 4010 2282
rect 3946 2222 3950 2278
rect 3950 2222 4006 2278
rect 4006 2222 4010 2278
rect 3946 2218 4010 2222
rect 890 1858 954 1862
rect 890 1802 894 1858
rect 894 1802 950 1858
rect 950 1802 954 1858
rect 890 1798 954 1802
rect 970 1858 1034 1862
rect 970 1802 974 1858
rect 974 1802 1030 1858
rect 1030 1802 1034 1858
rect 970 1798 1034 1802
rect 1050 1858 1114 1862
rect 1050 1802 1054 1858
rect 1054 1802 1110 1858
rect 1110 1802 1114 1858
rect 1050 1798 1114 1802
rect 1130 1858 1194 1862
rect 1130 1802 1134 1858
rect 1134 1802 1190 1858
rect 1190 1802 1194 1858
rect 1130 1798 1194 1802
rect 890 1778 954 1782
rect 890 1722 894 1778
rect 894 1722 950 1778
rect 950 1722 954 1778
rect 890 1718 954 1722
rect 970 1778 1034 1782
rect 970 1722 974 1778
rect 974 1722 1030 1778
rect 1030 1722 1034 1778
rect 970 1718 1034 1722
rect 1050 1778 1114 1782
rect 1050 1722 1054 1778
rect 1054 1722 1110 1778
rect 1110 1722 1114 1778
rect 1050 1718 1114 1722
rect 1130 1778 1194 1782
rect 1130 1722 1134 1778
rect 1134 1722 1190 1778
rect 1190 1722 1194 1778
rect 1130 1718 1194 1722
rect 890 1698 954 1702
rect 890 1642 894 1698
rect 894 1642 950 1698
rect 950 1642 954 1698
rect 890 1638 954 1642
rect 970 1698 1034 1702
rect 970 1642 974 1698
rect 974 1642 1030 1698
rect 1030 1642 1034 1698
rect 970 1638 1034 1642
rect 1050 1698 1114 1702
rect 1050 1642 1054 1698
rect 1054 1642 1110 1698
rect 1110 1642 1114 1698
rect 1050 1638 1114 1642
rect 1130 1698 1194 1702
rect 1130 1642 1134 1698
rect 1134 1642 1190 1698
rect 1190 1642 1194 1698
rect 1130 1638 1194 1642
rect 666 1508 730 1572
rect 890 1618 954 1622
rect 890 1562 894 1618
rect 894 1562 950 1618
rect 950 1562 954 1618
rect 890 1558 954 1562
rect 970 1618 1034 1622
rect 970 1562 974 1618
rect 974 1562 1030 1618
rect 1030 1562 1034 1618
rect 970 1558 1034 1562
rect 1050 1618 1114 1622
rect 1050 1562 1054 1618
rect 1054 1562 1110 1618
rect 1110 1562 1114 1618
rect 1050 1558 1114 1562
rect 1130 1618 1194 1622
rect 1130 1562 1134 1618
rect 1134 1562 1190 1618
rect 1190 1562 1194 1618
rect 1130 1558 1194 1562
rect 1594 1858 1658 1862
rect 1594 1802 1598 1858
rect 1598 1802 1654 1858
rect 1654 1802 1658 1858
rect 1594 1798 1658 1802
rect 1674 1858 1738 1862
rect 1674 1802 1678 1858
rect 1678 1802 1734 1858
rect 1734 1802 1738 1858
rect 1674 1798 1738 1802
rect 1754 1858 1818 1862
rect 1754 1802 1758 1858
rect 1758 1802 1814 1858
rect 1814 1802 1818 1858
rect 1754 1798 1818 1802
rect 1834 1858 1898 1862
rect 1834 1802 1838 1858
rect 1838 1802 1894 1858
rect 1894 1802 1898 1858
rect 1834 1798 1898 1802
rect 1594 1778 1658 1782
rect 1594 1722 1598 1778
rect 1598 1722 1654 1778
rect 1654 1722 1658 1778
rect 1594 1718 1658 1722
rect 1674 1778 1738 1782
rect 1674 1722 1678 1778
rect 1678 1722 1734 1778
rect 1734 1722 1738 1778
rect 1674 1718 1738 1722
rect 1754 1778 1818 1782
rect 1754 1722 1758 1778
rect 1758 1722 1814 1778
rect 1814 1722 1818 1778
rect 1754 1718 1818 1722
rect 1834 1778 1898 1782
rect 1834 1722 1838 1778
rect 1838 1722 1894 1778
rect 1894 1722 1898 1778
rect 1834 1718 1898 1722
rect 1594 1698 1658 1702
rect 1594 1642 1598 1698
rect 1598 1642 1654 1698
rect 1654 1642 1658 1698
rect 1594 1638 1658 1642
rect 1674 1698 1738 1702
rect 1674 1642 1678 1698
rect 1678 1642 1734 1698
rect 1734 1642 1738 1698
rect 1674 1638 1738 1642
rect 1754 1698 1818 1702
rect 1754 1642 1758 1698
rect 1758 1642 1814 1698
rect 1814 1642 1818 1698
rect 1754 1638 1818 1642
rect 1834 1698 1898 1702
rect 1834 1642 1838 1698
rect 1838 1642 1894 1698
rect 1894 1642 1898 1698
rect 1834 1638 1898 1642
rect 1594 1618 1658 1622
rect 1594 1562 1598 1618
rect 1598 1562 1654 1618
rect 1654 1562 1658 1618
rect 1594 1558 1658 1562
rect 1674 1618 1738 1622
rect 1674 1562 1678 1618
rect 1678 1562 1734 1618
rect 1734 1562 1738 1618
rect 1674 1558 1738 1562
rect 1754 1618 1818 1622
rect 1754 1562 1758 1618
rect 1758 1562 1814 1618
rect 1814 1562 1818 1618
rect 1754 1558 1818 1562
rect 1834 1618 1898 1622
rect 1834 1562 1838 1618
rect 1838 1562 1894 1618
rect 1894 1562 1898 1618
rect 1834 1558 1898 1562
rect 2298 1858 2362 1862
rect 2298 1802 2302 1858
rect 2302 1802 2358 1858
rect 2358 1802 2362 1858
rect 2298 1798 2362 1802
rect 2378 1858 2442 1862
rect 2378 1802 2382 1858
rect 2382 1802 2438 1858
rect 2438 1802 2442 1858
rect 2378 1798 2442 1802
rect 2458 1858 2522 1862
rect 2458 1802 2462 1858
rect 2462 1802 2518 1858
rect 2518 1802 2522 1858
rect 2458 1798 2522 1802
rect 2538 1858 2602 1862
rect 2538 1802 2542 1858
rect 2542 1802 2598 1858
rect 2598 1802 2602 1858
rect 2538 1798 2602 1802
rect 2298 1778 2362 1782
rect 2298 1722 2302 1778
rect 2302 1722 2358 1778
rect 2358 1722 2362 1778
rect 2298 1718 2362 1722
rect 2378 1778 2442 1782
rect 2378 1722 2382 1778
rect 2382 1722 2438 1778
rect 2438 1722 2442 1778
rect 2378 1718 2442 1722
rect 2458 1778 2522 1782
rect 2458 1722 2462 1778
rect 2462 1722 2518 1778
rect 2518 1722 2522 1778
rect 2458 1718 2522 1722
rect 2538 1778 2602 1782
rect 2538 1722 2542 1778
rect 2542 1722 2598 1778
rect 2598 1722 2602 1778
rect 2538 1718 2602 1722
rect 2298 1698 2362 1702
rect 2298 1642 2302 1698
rect 2302 1642 2358 1698
rect 2358 1642 2362 1698
rect 2298 1638 2362 1642
rect 2378 1698 2442 1702
rect 2378 1642 2382 1698
rect 2382 1642 2438 1698
rect 2438 1642 2442 1698
rect 2378 1638 2442 1642
rect 2458 1698 2522 1702
rect 2458 1642 2462 1698
rect 2462 1642 2518 1698
rect 2518 1642 2522 1698
rect 2458 1638 2522 1642
rect 2538 1698 2602 1702
rect 2538 1642 2542 1698
rect 2542 1642 2598 1698
rect 2598 1642 2602 1698
rect 2538 1638 2602 1642
rect 2298 1618 2362 1622
rect 2298 1562 2302 1618
rect 2302 1562 2358 1618
rect 2358 1562 2362 1618
rect 2298 1558 2362 1562
rect 2378 1618 2442 1622
rect 2378 1562 2382 1618
rect 2382 1562 2438 1618
rect 2438 1562 2442 1618
rect 2378 1558 2442 1562
rect 2458 1618 2522 1622
rect 2458 1562 2462 1618
rect 2462 1562 2518 1618
rect 2518 1562 2522 1618
rect 2458 1558 2522 1562
rect 2538 1618 2602 1622
rect 2538 1562 2542 1618
rect 2542 1562 2598 1618
rect 2598 1562 2602 1618
rect 2538 1558 2602 1562
rect 3002 1858 3066 1862
rect 3002 1802 3006 1858
rect 3006 1802 3062 1858
rect 3062 1802 3066 1858
rect 3002 1798 3066 1802
rect 3082 1858 3146 1862
rect 3082 1802 3086 1858
rect 3086 1802 3142 1858
rect 3142 1802 3146 1858
rect 3082 1798 3146 1802
rect 3162 1858 3226 1862
rect 3162 1802 3166 1858
rect 3166 1802 3222 1858
rect 3222 1802 3226 1858
rect 3162 1798 3226 1802
rect 3242 1858 3306 1862
rect 3242 1802 3246 1858
rect 3246 1802 3302 1858
rect 3302 1802 3306 1858
rect 3242 1798 3306 1802
rect 3002 1778 3066 1782
rect 3002 1722 3006 1778
rect 3006 1722 3062 1778
rect 3062 1722 3066 1778
rect 3002 1718 3066 1722
rect 3082 1778 3146 1782
rect 3082 1722 3086 1778
rect 3086 1722 3142 1778
rect 3142 1722 3146 1778
rect 3082 1718 3146 1722
rect 3162 1778 3226 1782
rect 3162 1722 3166 1778
rect 3166 1722 3222 1778
rect 3222 1722 3226 1778
rect 3162 1718 3226 1722
rect 3242 1778 3306 1782
rect 3242 1722 3246 1778
rect 3246 1722 3302 1778
rect 3302 1722 3306 1778
rect 3242 1718 3306 1722
rect 3002 1698 3066 1702
rect 3002 1642 3006 1698
rect 3006 1642 3062 1698
rect 3062 1642 3066 1698
rect 3002 1638 3066 1642
rect 3082 1698 3146 1702
rect 3082 1642 3086 1698
rect 3086 1642 3142 1698
rect 3142 1642 3146 1698
rect 3082 1638 3146 1642
rect 3162 1698 3226 1702
rect 3162 1642 3166 1698
rect 3166 1642 3222 1698
rect 3222 1642 3226 1698
rect 3162 1638 3226 1642
rect 3242 1698 3306 1702
rect 3242 1642 3246 1698
rect 3246 1642 3302 1698
rect 3302 1642 3306 1698
rect 3242 1638 3306 1642
rect 3002 1618 3066 1622
rect 3002 1562 3006 1618
rect 3006 1562 3062 1618
rect 3062 1562 3066 1618
rect 3002 1558 3066 1562
rect 3082 1618 3146 1622
rect 3082 1562 3086 1618
rect 3086 1562 3142 1618
rect 3142 1562 3146 1618
rect 3082 1558 3146 1562
rect 3162 1618 3226 1622
rect 3162 1562 3166 1618
rect 3166 1562 3222 1618
rect 3222 1562 3226 1618
rect 3162 1558 3226 1562
rect 3242 1618 3306 1622
rect 3242 1562 3246 1618
rect 3246 1562 3302 1618
rect 3302 1562 3306 1618
rect 3242 1558 3306 1562
rect 3706 1858 3770 1862
rect 3706 1802 3710 1858
rect 3710 1802 3766 1858
rect 3766 1802 3770 1858
rect 3706 1798 3770 1802
rect 3786 1858 3850 1862
rect 3786 1802 3790 1858
rect 3790 1802 3846 1858
rect 3846 1802 3850 1858
rect 3786 1798 3850 1802
rect 3866 1858 3930 1862
rect 3866 1802 3870 1858
rect 3870 1802 3926 1858
rect 3926 1802 3930 1858
rect 3866 1798 3930 1802
rect 3946 1858 4010 1862
rect 3946 1802 3950 1858
rect 3950 1802 4006 1858
rect 4006 1802 4010 1858
rect 3946 1798 4010 1802
rect 3706 1778 3770 1782
rect 3706 1722 3710 1778
rect 3710 1722 3766 1778
rect 3766 1722 3770 1778
rect 3706 1718 3770 1722
rect 3786 1778 3850 1782
rect 3786 1722 3790 1778
rect 3790 1722 3846 1778
rect 3846 1722 3850 1778
rect 3786 1718 3850 1722
rect 3866 1778 3930 1782
rect 3866 1722 3870 1778
rect 3870 1722 3926 1778
rect 3926 1722 3930 1778
rect 3866 1718 3930 1722
rect 3946 1778 4010 1782
rect 3946 1722 3950 1778
rect 3950 1722 4006 1778
rect 4006 1722 4010 1778
rect 3946 1718 4010 1722
rect 3706 1698 3770 1702
rect 3706 1642 3710 1698
rect 3710 1642 3766 1698
rect 3766 1642 3770 1698
rect 3706 1638 3770 1642
rect 3786 1698 3850 1702
rect 3786 1642 3790 1698
rect 3790 1642 3846 1698
rect 3846 1642 3850 1698
rect 3786 1638 3850 1642
rect 3866 1698 3930 1702
rect 3866 1642 3870 1698
rect 3870 1642 3926 1698
rect 3926 1642 3930 1698
rect 3866 1638 3930 1642
rect 3946 1698 4010 1702
rect 3946 1642 3950 1698
rect 3950 1642 4006 1698
rect 4006 1642 4010 1698
rect 3946 1638 4010 1642
rect 3706 1618 3770 1622
rect 3706 1562 3710 1618
rect 3710 1562 3766 1618
rect 3766 1562 3770 1618
rect 3706 1558 3770 1562
rect 3786 1618 3850 1622
rect 3786 1562 3790 1618
rect 3790 1562 3846 1618
rect 3846 1562 3850 1618
rect 3786 1558 3850 1562
rect 3866 1618 3930 1622
rect 3866 1562 3870 1618
rect 3870 1562 3926 1618
rect 3926 1562 3930 1618
rect 3866 1558 3930 1562
rect 3946 1618 4010 1622
rect 3946 1562 3950 1618
rect 3950 1562 4006 1618
rect 4006 1562 4010 1618
rect 3946 1558 4010 1562
rect 666 1428 730 1492
rect 666 1268 730 1332
rect 666 1188 730 1252
rect 890 1194 954 1198
rect 890 1138 894 1194
rect 894 1138 950 1194
rect 950 1138 954 1194
rect 890 1134 954 1138
rect 970 1194 1034 1198
rect 970 1138 974 1194
rect 974 1138 1030 1194
rect 1030 1138 1034 1194
rect 970 1134 1034 1138
rect 1050 1194 1114 1198
rect 1050 1138 1054 1194
rect 1054 1138 1110 1194
rect 1110 1138 1114 1194
rect 1050 1134 1114 1138
rect 1130 1194 1194 1198
rect 1130 1138 1134 1194
rect 1134 1138 1190 1194
rect 1190 1138 1194 1194
rect 1130 1134 1194 1138
rect 890 1114 954 1118
rect 890 1058 894 1114
rect 894 1058 950 1114
rect 950 1058 954 1114
rect 890 1054 954 1058
rect 970 1114 1034 1118
rect 970 1058 974 1114
rect 974 1058 1030 1114
rect 1030 1058 1034 1114
rect 970 1054 1034 1058
rect 1050 1114 1114 1118
rect 1050 1058 1054 1114
rect 1054 1058 1110 1114
rect 1110 1058 1114 1114
rect 1050 1054 1114 1058
rect 1130 1114 1194 1118
rect 1130 1058 1134 1114
rect 1134 1058 1190 1114
rect 1190 1058 1194 1114
rect 1130 1054 1194 1058
rect 890 1034 954 1038
rect 890 978 894 1034
rect 894 978 950 1034
rect 950 978 954 1034
rect 890 974 954 978
rect 970 1034 1034 1038
rect 970 978 974 1034
rect 974 978 1030 1034
rect 1030 978 1034 1034
rect 970 974 1034 978
rect 1050 1034 1114 1038
rect 1050 978 1054 1034
rect 1054 978 1110 1034
rect 1110 978 1114 1034
rect 1050 974 1114 978
rect 1130 1034 1194 1038
rect 1130 978 1134 1034
rect 1134 978 1190 1034
rect 1190 978 1194 1034
rect 1130 974 1194 978
rect 890 954 954 958
rect 890 898 894 954
rect 894 898 950 954
rect 950 898 954 954
rect 890 894 954 898
rect 970 954 1034 958
rect 970 898 974 954
rect 974 898 1030 954
rect 1030 898 1034 954
rect 970 894 1034 898
rect 1050 954 1114 958
rect 1050 898 1054 954
rect 1054 898 1110 954
rect 1110 898 1114 954
rect 1050 894 1114 898
rect 1130 954 1194 958
rect 1130 898 1134 954
rect 1134 898 1190 954
rect 1190 898 1194 954
rect 1130 894 1194 898
rect 1594 1194 1658 1198
rect 1594 1138 1598 1194
rect 1598 1138 1654 1194
rect 1654 1138 1658 1194
rect 1594 1134 1658 1138
rect 1674 1194 1738 1198
rect 1674 1138 1678 1194
rect 1678 1138 1734 1194
rect 1734 1138 1738 1194
rect 1674 1134 1738 1138
rect 1754 1194 1818 1198
rect 1754 1138 1758 1194
rect 1758 1138 1814 1194
rect 1814 1138 1818 1194
rect 1754 1134 1818 1138
rect 1834 1194 1898 1198
rect 1834 1138 1838 1194
rect 1838 1138 1894 1194
rect 1894 1138 1898 1194
rect 1834 1134 1898 1138
rect 1594 1114 1658 1118
rect 1594 1058 1598 1114
rect 1598 1058 1654 1114
rect 1654 1058 1658 1114
rect 1594 1054 1658 1058
rect 1674 1114 1738 1118
rect 1674 1058 1678 1114
rect 1678 1058 1734 1114
rect 1734 1058 1738 1114
rect 1674 1054 1738 1058
rect 1754 1114 1818 1118
rect 1754 1058 1758 1114
rect 1758 1058 1814 1114
rect 1814 1058 1818 1114
rect 1754 1054 1818 1058
rect 1834 1114 1898 1118
rect 1834 1058 1838 1114
rect 1838 1058 1894 1114
rect 1894 1058 1898 1114
rect 1834 1054 1898 1058
rect 1594 1034 1658 1038
rect 1594 978 1598 1034
rect 1598 978 1654 1034
rect 1654 978 1658 1034
rect 1594 974 1658 978
rect 1674 1034 1738 1038
rect 1674 978 1678 1034
rect 1678 978 1734 1034
rect 1734 978 1738 1034
rect 1674 974 1738 978
rect 1754 1034 1818 1038
rect 1754 978 1758 1034
rect 1758 978 1814 1034
rect 1814 978 1818 1034
rect 1754 974 1818 978
rect 1834 1034 1898 1038
rect 1834 978 1838 1034
rect 1838 978 1894 1034
rect 1894 978 1898 1034
rect 1834 974 1898 978
rect 1594 954 1658 958
rect 1594 898 1598 954
rect 1598 898 1654 954
rect 1654 898 1658 954
rect 1594 894 1658 898
rect 1674 954 1738 958
rect 1674 898 1678 954
rect 1678 898 1734 954
rect 1734 898 1738 954
rect 1674 894 1738 898
rect 1754 954 1818 958
rect 1754 898 1758 954
rect 1758 898 1814 954
rect 1814 898 1818 954
rect 1754 894 1818 898
rect 1834 954 1898 958
rect 1834 898 1838 954
rect 1838 898 1894 954
rect 1894 898 1898 954
rect 1834 894 1898 898
rect 3002 1194 3066 1198
rect 3002 1138 3006 1194
rect 3006 1138 3062 1194
rect 3062 1138 3066 1194
rect 3002 1134 3066 1138
rect 3082 1194 3146 1198
rect 3082 1138 3086 1194
rect 3086 1138 3142 1194
rect 3142 1138 3146 1194
rect 3082 1134 3146 1138
rect 3162 1194 3226 1198
rect 3162 1138 3166 1194
rect 3166 1138 3222 1194
rect 3222 1138 3226 1194
rect 3162 1134 3226 1138
rect 3242 1194 3306 1198
rect 3242 1138 3246 1194
rect 3246 1138 3302 1194
rect 3302 1138 3306 1194
rect 3242 1134 3306 1138
rect 3002 1114 3066 1118
rect 3002 1058 3006 1114
rect 3006 1058 3062 1114
rect 3062 1058 3066 1114
rect 3002 1054 3066 1058
rect 3082 1114 3146 1118
rect 3082 1058 3086 1114
rect 3086 1058 3142 1114
rect 3142 1058 3146 1114
rect 3082 1054 3146 1058
rect 3162 1114 3226 1118
rect 3162 1058 3166 1114
rect 3166 1058 3222 1114
rect 3222 1058 3226 1114
rect 3162 1054 3226 1058
rect 3242 1114 3306 1118
rect 3242 1058 3246 1114
rect 3246 1058 3302 1114
rect 3302 1058 3306 1114
rect 3242 1054 3306 1058
rect 3002 1034 3066 1038
rect 3002 978 3006 1034
rect 3006 978 3062 1034
rect 3062 978 3066 1034
rect 3002 974 3066 978
rect 3082 1034 3146 1038
rect 3082 978 3086 1034
rect 3086 978 3142 1034
rect 3142 978 3146 1034
rect 3082 974 3146 978
rect 3162 1034 3226 1038
rect 3162 978 3166 1034
rect 3166 978 3222 1034
rect 3222 978 3226 1034
rect 3162 974 3226 978
rect 3242 1034 3306 1038
rect 3242 978 3246 1034
rect 3246 978 3302 1034
rect 3302 978 3306 1034
rect 3242 974 3306 978
rect 3002 954 3066 958
rect 3002 898 3006 954
rect 3006 898 3062 954
rect 3062 898 3066 954
rect 3002 894 3066 898
rect 3082 954 3146 958
rect 3082 898 3086 954
rect 3086 898 3142 954
rect 3142 898 3146 954
rect 3082 894 3146 898
rect 3162 954 3226 958
rect 3162 898 3166 954
rect 3166 898 3222 954
rect 3222 898 3226 954
rect 3162 894 3226 898
rect 3242 954 3306 958
rect 3242 898 3246 954
rect 3246 898 3302 954
rect 3302 898 3306 954
rect 3242 894 3306 898
rect 3706 1194 3770 1198
rect 3706 1138 3710 1194
rect 3710 1138 3766 1194
rect 3766 1138 3770 1194
rect 3706 1134 3770 1138
rect 3786 1194 3850 1198
rect 3786 1138 3790 1194
rect 3790 1138 3846 1194
rect 3846 1138 3850 1194
rect 3786 1134 3850 1138
rect 3866 1194 3930 1198
rect 3866 1138 3870 1194
rect 3870 1138 3926 1194
rect 3926 1138 3930 1194
rect 3866 1134 3930 1138
rect 3946 1194 4010 1198
rect 3946 1138 3950 1194
rect 3950 1138 4006 1194
rect 4006 1138 4010 1194
rect 3946 1134 4010 1138
rect 3706 1114 3770 1118
rect 3706 1058 3710 1114
rect 3710 1058 3766 1114
rect 3766 1058 3770 1114
rect 3706 1054 3770 1058
rect 3786 1114 3850 1118
rect 3786 1058 3790 1114
rect 3790 1058 3846 1114
rect 3846 1058 3850 1114
rect 3786 1054 3850 1058
rect 3866 1114 3930 1118
rect 3866 1058 3870 1114
rect 3870 1058 3926 1114
rect 3926 1058 3930 1114
rect 3866 1054 3930 1058
rect 3946 1114 4010 1118
rect 3946 1058 3950 1114
rect 3950 1058 4006 1114
rect 4006 1058 4010 1114
rect 3946 1054 4010 1058
rect 3706 1034 3770 1038
rect 3706 978 3710 1034
rect 3710 978 3766 1034
rect 3766 978 3770 1034
rect 3706 974 3770 978
rect 3786 1034 3850 1038
rect 3786 978 3790 1034
rect 3790 978 3846 1034
rect 3846 978 3850 1034
rect 3786 974 3850 978
rect 3866 1034 3930 1038
rect 3866 978 3870 1034
rect 3870 978 3926 1034
rect 3926 978 3930 1034
rect 3866 974 3930 978
rect 3946 1034 4010 1038
rect 3946 978 3950 1034
rect 3950 978 4006 1034
rect 4006 978 4010 1034
rect 3946 974 4010 978
rect 3706 954 3770 958
rect 3706 898 3710 954
rect 3710 898 3766 954
rect 3766 898 3770 954
rect 3706 894 3770 898
rect 3786 954 3850 958
rect 3786 898 3790 954
rect 3790 898 3846 954
rect 3846 898 3850 954
rect 3786 894 3850 898
rect 3866 954 3930 958
rect 3866 898 3870 954
rect 3870 898 3926 954
rect 3926 898 3930 954
rect 3866 894 3930 898
rect 3946 954 4010 958
rect 3946 898 3950 954
rect 3950 898 4006 954
rect 4006 898 4010 954
rect 3946 894 4010 898
rect 890 536 954 540
rect 890 480 894 536
rect 894 480 950 536
rect 950 480 954 536
rect 890 476 954 480
rect 970 536 1034 540
rect 970 480 974 536
rect 974 480 1030 536
rect 1030 480 1034 536
rect 970 476 1034 480
rect 1050 536 1114 540
rect 1050 480 1054 536
rect 1054 480 1110 536
rect 1110 480 1114 536
rect 1050 476 1114 480
rect 1130 536 1194 540
rect 1130 480 1134 536
rect 1134 480 1190 536
rect 1190 480 1194 536
rect 1130 476 1194 480
rect 890 456 954 460
rect 890 400 894 456
rect 894 400 950 456
rect 950 400 954 456
rect 890 396 954 400
rect 970 456 1034 460
rect 970 400 974 456
rect 974 400 1030 456
rect 1030 400 1034 456
rect 970 396 1034 400
rect 1050 456 1114 460
rect 1050 400 1054 456
rect 1054 400 1110 456
rect 1110 400 1114 456
rect 1050 396 1114 400
rect 1130 456 1194 460
rect 1130 400 1134 456
rect 1134 400 1190 456
rect 1190 400 1194 456
rect 1130 396 1194 400
rect 890 376 954 380
rect 890 320 894 376
rect 894 320 950 376
rect 950 320 954 376
rect 890 316 954 320
rect 970 376 1034 380
rect 970 320 974 376
rect 974 320 1030 376
rect 1030 320 1034 376
rect 970 316 1034 320
rect 1050 376 1114 380
rect 1050 320 1054 376
rect 1054 320 1110 376
rect 1110 320 1114 376
rect 1050 316 1114 320
rect 1130 376 1194 380
rect 1130 320 1134 376
rect 1134 320 1190 376
rect 1190 320 1194 376
rect 1130 316 1194 320
rect 666 182 730 246
rect 890 296 954 300
rect 890 240 894 296
rect 894 240 950 296
rect 950 240 954 296
rect 890 236 954 240
rect 970 296 1034 300
rect 970 240 974 296
rect 974 240 1030 296
rect 1030 240 1034 296
rect 970 236 1034 240
rect 1050 296 1114 300
rect 1050 240 1054 296
rect 1054 240 1110 296
rect 1110 240 1114 296
rect 1050 236 1114 240
rect 1130 296 1194 300
rect 1130 240 1134 296
rect 1134 240 1190 296
rect 1190 240 1194 296
rect 1130 236 1194 240
rect 1594 536 1658 540
rect 1594 480 1598 536
rect 1598 480 1654 536
rect 1654 480 1658 536
rect 1594 476 1658 480
rect 1674 536 1738 540
rect 1674 480 1678 536
rect 1678 480 1734 536
rect 1734 480 1738 536
rect 1674 476 1738 480
rect 1754 536 1818 540
rect 1754 480 1758 536
rect 1758 480 1814 536
rect 1814 480 1818 536
rect 1754 476 1818 480
rect 1834 536 1898 540
rect 1834 480 1838 536
rect 1838 480 1894 536
rect 1894 480 1898 536
rect 1834 476 1898 480
rect 1594 456 1658 460
rect 1594 400 1598 456
rect 1598 400 1654 456
rect 1654 400 1658 456
rect 1594 396 1658 400
rect 1674 456 1738 460
rect 1674 400 1678 456
rect 1678 400 1734 456
rect 1734 400 1738 456
rect 1674 396 1738 400
rect 1754 456 1818 460
rect 1754 400 1758 456
rect 1758 400 1814 456
rect 1814 400 1818 456
rect 1754 396 1818 400
rect 1834 456 1898 460
rect 1834 400 1838 456
rect 1838 400 1894 456
rect 1894 400 1898 456
rect 1834 396 1898 400
rect 1594 376 1658 380
rect 1594 320 1598 376
rect 1598 320 1654 376
rect 1654 320 1658 376
rect 1594 316 1658 320
rect 1674 376 1738 380
rect 1674 320 1678 376
rect 1678 320 1734 376
rect 1734 320 1738 376
rect 1674 316 1738 320
rect 1754 376 1818 380
rect 1754 320 1758 376
rect 1758 320 1814 376
rect 1814 320 1818 376
rect 1754 316 1818 320
rect 1834 376 1898 380
rect 1834 320 1838 376
rect 1838 320 1894 376
rect 1894 320 1898 376
rect 1834 316 1898 320
rect 1594 296 1658 300
rect 1594 240 1598 296
rect 1598 240 1654 296
rect 1654 240 1658 296
rect 1594 236 1658 240
rect 1674 296 1738 300
rect 1674 240 1678 296
rect 1678 240 1734 296
rect 1734 240 1738 296
rect 1674 236 1738 240
rect 1754 296 1818 300
rect 1754 240 1758 296
rect 1758 240 1814 296
rect 1814 240 1818 296
rect 1754 236 1818 240
rect 1834 296 1898 300
rect 1834 240 1838 296
rect 1838 240 1894 296
rect 1894 240 1898 296
rect 1834 236 1898 240
rect 3002 536 3066 540
rect 3002 480 3006 536
rect 3006 480 3062 536
rect 3062 480 3066 536
rect 3002 476 3066 480
rect 3082 536 3146 540
rect 3082 480 3086 536
rect 3086 480 3142 536
rect 3142 480 3146 536
rect 3082 476 3146 480
rect 3162 536 3226 540
rect 3162 480 3166 536
rect 3166 480 3222 536
rect 3222 480 3226 536
rect 3162 476 3226 480
rect 3242 536 3306 540
rect 3242 480 3246 536
rect 3246 480 3302 536
rect 3302 480 3306 536
rect 3242 476 3306 480
rect 3002 456 3066 460
rect 3002 400 3006 456
rect 3006 400 3062 456
rect 3062 400 3066 456
rect 3002 396 3066 400
rect 3082 456 3146 460
rect 3082 400 3086 456
rect 3086 400 3142 456
rect 3142 400 3146 456
rect 3082 396 3146 400
rect 3162 456 3226 460
rect 3162 400 3166 456
rect 3166 400 3222 456
rect 3222 400 3226 456
rect 3162 396 3226 400
rect 3242 456 3306 460
rect 3242 400 3246 456
rect 3246 400 3302 456
rect 3302 400 3306 456
rect 3242 396 3306 400
rect 3002 376 3066 380
rect 3002 320 3006 376
rect 3006 320 3062 376
rect 3062 320 3066 376
rect 3002 316 3066 320
rect 3082 376 3146 380
rect 3082 320 3086 376
rect 3086 320 3142 376
rect 3142 320 3146 376
rect 3082 316 3146 320
rect 3162 376 3226 380
rect 3162 320 3166 376
rect 3166 320 3222 376
rect 3222 320 3226 376
rect 3162 316 3226 320
rect 3242 376 3306 380
rect 3242 320 3246 376
rect 3246 320 3302 376
rect 3302 320 3306 376
rect 3242 316 3306 320
rect 3002 296 3066 300
rect 3002 240 3006 296
rect 3006 240 3062 296
rect 3062 240 3066 296
rect 3002 236 3066 240
rect 3082 296 3146 300
rect 3082 240 3086 296
rect 3086 240 3142 296
rect 3142 240 3146 296
rect 3082 236 3146 240
rect 3162 296 3226 300
rect 3162 240 3166 296
rect 3166 240 3222 296
rect 3222 240 3226 296
rect 3162 236 3226 240
rect 3242 296 3306 300
rect 3242 240 3246 296
rect 3246 240 3302 296
rect 3302 240 3306 296
rect 3242 236 3306 240
rect 3706 536 3770 540
rect 3706 480 3710 536
rect 3710 480 3766 536
rect 3766 480 3770 536
rect 3706 476 3770 480
rect 3786 536 3850 540
rect 3786 480 3790 536
rect 3790 480 3846 536
rect 3846 480 3850 536
rect 3786 476 3850 480
rect 3866 536 3930 540
rect 3866 480 3870 536
rect 3870 480 3926 536
rect 3926 480 3930 536
rect 3866 476 3930 480
rect 3946 536 4010 540
rect 3946 480 3950 536
rect 3950 480 4006 536
rect 4006 480 4010 536
rect 3946 476 4010 480
rect 3706 456 3770 460
rect 3706 400 3710 456
rect 3710 400 3766 456
rect 3766 400 3770 456
rect 3706 396 3770 400
rect 3786 456 3850 460
rect 3786 400 3790 456
rect 3790 400 3846 456
rect 3846 400 3850 456
rect 3786 396 3850 400
rect 3866 456 3930 460
rect 3866 400 3870 456
rect 3870 400 3926 456
rect 3926 400 3930 456
rect 3866 396 3930 400
rect 3946 456 4010 460
rect 3946 400 3950 456
rect 3950 400 4006 456
rect 4006 400 4010 456
rect 3946 396 4010 400
rect 3706 376 3770 380
rect 3706 320 3710 376
rect 3710 320 3766 376
rect 3766 320 3770 376
rect 3706 316 3770 320
rect 3786 376 3850 380
rect 3786 320 3790 376
rect 3790 320 3846 376
rect 3846 320 3850 376
rect 3786 316 3850 320
rect 3866 376 3930 380
rect 3866 320 3870 376
rect 3870 320 3926 376
rect 3926 320 3930 376
rect 3866 316 3930 320
rect 3946 376 4010 380
rect 3946 320 3950 376
rect 3950 320 4006 376
rect 4006 320 4010 376
rect 3946 316 4010 320
rect 3706 296 3770 300
rect 3706 240 3710 296
rect 3710 240 3766 296
rect 3766 240 3770 296
rect 3706 236 3770 240
rect 3786 296 3850 300
rect 3786 240 3790 296
rect 3790 240 3846 296
rect 3846 240 3850 296
rect 3786 236 3850 240
rect 3866 296 3930 300
rect 3866 240 3870 296
rect 3870 240 3926 296
rect 3926 240 3930 296
rect 3866 236 3930 240
rect 3946 296 4010 300
rect 3946 240 3950 296
rect 3950 240 4006 296
rect 4006 240 4010 296
rect 3946 236 4010 240
rect 666 102 730 166
rect 244 -192 308 -128
rect 370 -192 434 -128
rect 244 -296 308 -232
rect 370 -296 434 -232
rect 244 -380 308 -316
rect 370 -380 434 -316
rect 244 -466 308 -402
rect 370 -466 434 -402
rect 244 -560 308 -496
rect 370 -560 434 -496
rect 244 -660 308 -596
rect 370 -660 434 -596
rect 244 -744 308 -680
rect 370 -744 434 -680
rect 852 -130 916 -128
rect 852 -190 854 -130
rect 854 -190 914 -130
rect 914 -190 916 -130
rect 852 -192 916 -190
rect 978 -130 1042 -128
rect 978 -190 980 -130
rect 980 -190 1040 -130
rect 1040 -190 1042 -130
rect 978 -192 1042 -190
rect 852 -234 916 -232
rect 852 -294 854 -234
rect 854 -294 914 -234
rect 914 -294 916 -234
rect 852 -296 916 -294
rect 978 -234 1042 -232
rect 978 -294 980 -234
rect 980 -294 1040 -234
rect 1040 -294 1042 -234
rect 978 -296 1042 -294
rect 852 -318 916 -316
rect 852 -378 854 -318
rect 854 -378 914 -318
rect 914 -378 916 -318
rect 852 -380 916 -378
rect 978 -318 1042 -316
rect 978 -378 980 -318
rect 980 -378 1040 -318
rect 1040 -378 1042 -318
rect 978 -380 1042 -378
rect 852 -404 916 -402
rect 852 -464 854 -404
rect 854 -464 914 -404
rect 914 -464 916 -404
rect 852 -466 916 -464
rect 978 -404 1042 -402
rect 978 -464 980 -404
rect 980 -464 1040 -404
rect 1040 -464 1042 -404
rect 978 -466 1042 -464
rect 852 -498 916 -496
rect 852 -558 854 -498
rect 854 -558 914 -498
rect 914 -558 916 -498
rect 852 -560 916 -558
rect 978 -498 1042 -496
rect 978 -558 980 -498
rect 980 -558 1040 -498
rect 1040 -558 1042 -498
rect 978 -560 1042 -558
rect 852 -598 916 -596
rect 852 -658 854 -598
rect 854 -658 914 -598
rect 914 -658 916 -598
rect 852 -660 916 -658
rect 978 -598 1042 -596
rect 978 -658 980 -598
rect 980 -658 1040 -598
rect 1040 -658 1042 -598
rect 978 -660 1042 -658
rect 852 -682 916 -680
rect 852 -742 854 -682
rect 854 -742 914 -682
rect 914 -742 916 -682
rect 852 -744 916 -742
rect 978 -682 1042 -680
rect 978 -742 980 -682
rect 980 -742 1040 -682
rect 1040 -742 1042 -682
rect 978 -744 1042 -742
rect 1702 -130 1766 -128
rect 1702 -190 1704 -130
rect 1704 -190 1764 -130
rect 1764 -190 1766 -130
rect 1702 -192 1766 -190
rect 1828 -130 1892 -128
rect 1828 -190 1830 -130
rect 1830 -190 1890 -130
rect 1890 -190 1892 -130
rect 1828 -192 1892 -190
rect 1702 -234 1766 -232
rect 1702 -294 1704 -234
rect 1704 -294 1764 -234
rect 1764 -294 1766 -234
rect 1702 -296 1766 -294
rect 1828 -234 1892 -232
rect 1828 -294 1830 -234
rect 1830 -294 1890 -234
rect 1890 -294 1892 -234
rect 1828 -296 1892 -294
rect 1702 -318 1766 -316
rect 1702 -378 1704 -318
rect 1704 -378 1764 -318
rect 1764 -378 1766 -318
rect 1702 -380 1766 -378
rect 1828 -318 1892 -316
rect 1828 -378 1830 -318
rect 1830 -378 1890 -318
rect 1890 -378 1892 -318
rect 1828 -380 1892 -378
rect 1702 -404 1766 -402
rect 1702 -464 1704 -404
rect 1704 -464 1764 -404
rect 1764 -464 1766 -404
rect 1702 -466 1766 -464
rect 1828 -404 1892 -402
rect 1828 -464 1830 -404
rect 1830 -464 1890 -404
rect 1890 -464 1892 -404
rect 1828 -466 1892 -464
rect 1702 -498 1766 -496
rect 1702 -558 1704 -498
rect 1704 -558 1764 -498
rect 1764 -558 1766 -498
rect 1702 -560 1766 -558
rect 1828 -498 1892 -496
rect 1828 -558 1830 -498
rect 1830 -558 1890 -498
rect 1890 -558 1892 -498
rect 1828 -560 1892 -558
rect 1702 -598 1766 -596
rect 1702 -658 1704 -598
rect 1704 -658 1764 -598
rect 1764 -658 1766 -598
rect 1702 -660 1766 -658
rect 1828 -598 1892 -596
rect 1828 -658 1830 -598
rect 1830 -658 1890 -598
rect 1890 -658 1892 -598
rect 1828 -660 1892 -658
rect 1702 -682 1766 -680
rect 1702 -742 1704 -682
rect 1704 -742 1764 -682
rect 1764 -742 1766 -682
rect 1702 -744 1766 -742
rect 1828 -682 1892 -680
rect 1828 -742 1830 -682
rect 1830 -742 1890 -682
rect 1890 -742 1892 -682
rect 1828 -744 1892 -742
rect 2372 -130 2436 -128
rect 2372 -190 2374 -130
rect 2374 -190 2434 -130
rect 2434 -190 2436 -130
rect 2372 -192 2436 -190
rect 2498 -130 2562 -128
rect 2498 -190 2500 -130
rect 2500 -190 2560 -130
rect 2560 -190 2562 -130
rect 2498 -192 2562 -190
rect 2372 -234 2436 -232
rect 2372 -294 2374 -234
rect 2374 -294 2434 -234
rect 2434 -294 2436 -234
rect 2372 -296 2436 -294
rect 2498 -234 2562 -232
rect 2498 -294 2500 -234
rect 2500 -294 2560 -234
rect 2560 -294 2562 -234
rect 2498 -296 2562 -294
rect 2372 -318 2436 -316
rect 2372 -378 2374 -318
rect 2374 -378 2434 -318
rect 2434 -378 2436 -318
rect 2372 -380 2436 -378
rect 2498 -318 2562 -316
rect 2498 -378 2500 -318
rect 2500 -378 2560 -318
rect 2560 -378 2562 -318
rect 2498 -380 2562 -378
rect 2372 -404 2436 -402
rect 2372 -464 2374 -404
rect 2374 -464 2434 -404
rect 2434 -464 2436 -404
rect 2372 -466 2436 -464
rect 2498 -404 2562 -402
rect 2498 -464 2500 -404
rect 2500 -464 2560 -404
rect 2560 -464 2562 -404
rect 2498 -466 2562 -464
rect 2372 -498 2436 -496
rect 2372 -558 2374 -498
rect 2374 -558 2434 -498
rect 2434 -558 2436 -498
rect 2372 -560 2436 -558
rect 2498 -498 2562 -496
rect 2498 -558 2500 -498
rect 2500 -558 2560 -498
rect 2560 -558 2562 -498
rect 2498 -560 2562 -558
rect 2372 -598 2436 -596
rect 2372 -658 2374 -598
rect 2374 -658 2434 -598
rect 2434 -658 2436 -598
rect 2372 -660 2436 -658
rect 2498 -598 2562 -596
rect 2498 -658 2500 -598
rect 2500 -658 2560 -598
rect 2560 -658 2562 -598
rect 2498 -660 2562 -658
rect 2372 -682 2436 -680
rect 2372 -742 2374 -682
rect 2374 -742 2434 -682
rect 2434 -742 2436 -682
rect 2372 -744 2436 -742
rect 2498 -682 2562 -680
rect 2498 -742 2500 -682
rect 2500 -742 2560 -682
rect 2560 -742 2562 -682
rect 2498 -744 2562 -742
rect 2886 -130 2950 -128
rect 2886 -190 2888 -130
rect 2888 -190 2948 -130
rect 2948 -190 2950 -130
rect 2886 -192 2950 -190
rect 3012 -130 3076 -128
rect 3012 -190 3014 -130
rect 3014 -190 3074 -130
rect 3074 -190 3076 -130
rect 3012 -192 3076 -190
rect 2886 -234 2950 -232
rect 2886 -294 2888 -234
rect 2888 -294 2948 -234
rect 2948 -294 2950 -234
rect 2886 -296 2950 -294
rect 3012 -234 3076 -232
rect 3012 -294 3014 -234
rect 3014 -294 3074 -234
rect 3074 -294 3076 -234
rect 3012 -296 3076 -294
rect 2886 -318 2950 -316
rect 2886 -378 2888 -318
rect 2888 -378 2948 -318
rect 2948 -378 2950 -318
rect 2886 -380 2950 -378
rect 3012 -318 3076 -316
rect 3012 -378 3014 -318
rect 3014 -378 3074 -318
rect 3074 -378 3076 -318
rect 3012 -380 3076 -378
rect 2886 -404 2950 -402
rect 2886 -464 2888 -404
rect 2888 -464 2948 -404
rect 2948 -464 2950 -404
rect 2886 -466 2950 -464
rect 3012 -404 3076 -402
rect 3012 -464 3014 -404
rect 3014 -464 3074 -404
rect 3074 -464 3076 -404
rect 3012 -466 3076 -464
rect 2886 -498 2950 -496
rect 2886 -558 2888 -498
rect 2888 -558 2948 -498
rect 2948 -558 2950 -498
rect 2886 -560 2950 -558
rect 3012 -498 3076 -496
rect 3012 -558 3014 -498
rect 3014 -558 3074 -498
rect 3074 -558 3076 -498
rect 3012 -560 3076 -558
rect 2886 -598 2950 -596
rect 2886 -658 2888 -598
rect 2888 -658 2948 -598
rect 2948 -658 2950 -598
rect 2886 -660 2950 -658
rect 3012 -598 3076 -596
rect 3012 -658 3014 -598
rect 3014 -658 3074 -598
rect 3074 -658 3076 -598
rect 3012 -660 3076 -658
rect 2886 -682 2950 -680
rect 2886 -742 2888 -682
rect 2888 -742 2948 -682
rect 2948 -742 2950 -682
rect 2886 -744 2950 -742
rect 3012 -682 3076 -680
rect 3012 -742 3014 -682
rect 3014 -742 3074 -682
rect 3074 -742 3076 -682
rect 3012 -744 3076 -742
rect 3706 -130 3770 -128
rect 3706 -190 3708 -130
rect 3708 -190 3768 -130
rect 3768 -190 3770 -130
rect 3706 -192 3770 -190
rect 3832 -130 3896 -128
rect 3832 -190 3834 -130
rect 3834 -190 3894 -130
rect 3894 -190 3896 -130
rect 3832 -192 3896 -190
rect 3706 -234 3770 -232
rect 3706 -294 3708 -234
rect 3708 -294 3768 -234
rect 3768 -294 3770 -234
rect 3706 -296 3770 -294
rect 3832 -234 3896 -232
rect 3832 -294 3834 -234
rect 3834 -294 3894 -234
rect 3894 -294 3896 -234
rect 3832 -296 3896 -294
rect 3706 -318 3770 -316
rect 3706 -378 3708 -318
rect 3708 -378 3768 -318
rect 3768 -378 3770 -318
rect 3706 -380 3770 -378
rect 3832 -318 3896 -316
rect 3832 -378 3834 -318
rect 3834 -378 3894 -318
rect 3894 -378 3896 -318
rect 3832 -380 3896 -378
rect 3706 -404 3770 -402
rect 3706 -464 3708 -404
rect 3708 -464 3768 -404
rect 3768 -464 3770 -404
rect 3706 -466 3770 -464
rect 3832 -404 3896 -402
rect 3832 -464 3834 -404
rect 3834 -464 3894 -404
rect 3894 -464 3896 -404
rect 3832 -466 3896 -464
rect 3706 -498 3770 -496
rect 3706 -558 3708 -498
rect 3708 -558 3768 -498
rect 3768 -558 3770 -498
rect 3706 -560 3770 -558
rect 3832 -498 3896 -496
rect 3832 -558 3834 -498
rect 3834 -558 3894 -498
rect 3894 -558 3896 -498
rect 3832 -560 3896 -558
rect 3706 -598 3770 -596
rect 3706 -658 3708 -598
rect 3708 -658 3768 -598
rect 3768 -658 3770 -598
rect 3706 -660 3770 -658
rect 3832 -598 3896 -596
rect 3832 -658 3834 -598
rect 3834 -658 3894 -598
rect 3894 -658 3896 -598
rect 3832 -660 3896 -658
rect 3706 -682 3770 -680
rect 3706 -742 3708 -682
rect 3708 -742 3768 -682
rect 3768 -742 3770 -682
rect 3706 -744 3770 -742
rect 3832 -682 3896 -680
rect 3832 -742 3834 -682
rect 3834 -742 3894 -682
rect 3894 -742 3896 -682
rect 3832 -744 3896 -742
rect 4464 -192 4528 -128
rect 4590 -192 4654 -128
rect 4464 -296 4528 -232
rect 4590 -296 4654 -232
rect 4464 -380 4528 -316
rect 4590 -380 4654 -316
rect 4464 -466 4528 -402
rect 4590 -466 4654 -402
rect 4464 -560 4528 -496
rect 4590 -560 4654 -496
rect 4464 -660 4528 -596
rect 4590 -660 4654 -596
rect 4464 -744 4528 -680
rect 4590 -744 4654 -680
<< metal4 >>
rect 526 3142 860 3192
rect 526 2906 574 3142
rect 810 2906 860 3142
rect 526 2858 860 2906
rect 2014 3144 2704 3194
rect 2014 2908 2088 3144
rect 2324 2908 2418 3144
rect 2654 2908 2704 3144
rect 2014 2858 2704 2908
rect 658 2744 724 2858
rect 658 2736 738 2744
rect 658 2672 666 2736
rect 730 2672 738 2736
rect 658 2656 738 2672
rect 658 2592 666 2656
rect 730 2592 738 2656
rect 658 2584 738 2592
rect 0 1832 334 1878
rect 0 1596 48 1832
rect 284 1596 334 1832
rect 0 1488 334 1596
rect 0 1252 46 1488
rect 282 1252 334 1488
rect 0 522 334 1252
rect 0 286 52 522
rect 288 286 334 522
rect 0 180 334 286
rect 0 76 46 180
rect -2 -56 46 76
rect 282 -56 334 180
rect 658 1580 724 2584
rect 842 2522 1242 2538
rect 842 2458 890 2522
rect 954 2484 970 2522
rect 1034 2484 1050 2522
rect 1114 2484 1130 2522
rect 1194 2458 1242 2522
rect 842 2442 896 2458
rect 1188 2442 1242 2458
rect 842 2378 890 2442
rect 1194 2378 1242 2442
rect 842 2362 896 2378
rect 1188 2362 1242 2378
rect 842 2298 890 2362
rect 1194 2298 1242 2362
rect 842 2282 896 2298
rect 1188 2282 1242 2298
rect 842 2218 890 2282
rect 954 2218 970 2228
rect 1034 2218 1050 2228
rect 1114 2218 1130 2228
rect 1194 2218 1242 2282
rect 842 2202 1242 2218
rect 1546 2522 1946 2538
rect 1546 2458 1594 2522
rect 1658 2484 1674 2522
rect 1738 2484 1754 2522
rect 1818 2484 1834 2522
rect 1898 2458 1946 2522
rect 1546 2442 1600 2458
rect 1892 2442 1946 2458
rect 1546 2378 1594 2442
rect 1898 2378 1946 2442
rect 1546 2362 1600 2378
rect 1892 2362 1946 2378
rect 1546 2298 1594 2362
rect 1898 2298 1946 2362
rect 1546 2282 1600 2298
rect 1892 2282 1946 2298
rect 1546 2218 1594 2282
rect 1658 2218 1674 2228
rect 1738 2218 1754 2228
rect 1818 2218 1834 2228
rect 1898 2218 1946 2282
rect 1546 2202 1946 2218
rect 2196 2522 2704 2858
rect 4566 2820 4900 2874
rect 4566 2584 4612 2820
rect 4848 2584 4900 2820
rect 2196 2458 2298 2522
rect 2362 2458 2378 2522
rect 2442 2458 2458 2522
rect 2522 2458 2538 2522
rect 2602 2458 2704 2522
rect 2196 2442 2704 2458
rect 2196 2378 2298 2442
rect 2362 2378 2378 2442
rect 2442 2378 2458 2442
rect 2522 2378 2538 2442
rect 2602 2378 2704 2442
rect 2196 2362 2704 2378
rect 2196 2298 2298 2362
rect 2362 2298 2378 2362
rect 2442 2298 2458 2362
rect 2522 2298 2538 2362
rect 2602 2298 2704 2362
rect 2196 2282 2704 2298
rect 2196 2218 2298 2282
rect 2362 2218 2378 2282
rect 2442 2218 2458 2282
rect 2522 2218 2538 2282
rect 2602 2218 2704 2282
rect 2196 2066 2704 2218
rect 2954 2522 3354 2538
rect 2954 2458 3002 2522
rect 3066 2484 3082 2522
rect 3146 2484 3162 2522
rect 3226 2484 3242 2522
rect 3306 2458 3354 2522
rect 2954 2442 3008 2458
rect 3300 2442 3354 2458
rect 2954 2378 3002 2442
rect 3306 2378 3354 2442
rect 2954 2362 3008 2378
rect 3300 2362 3354 2378
rect 2954 2298 3002 2362
rect 3306 2298 3354 2362
rect 2954 2282 3008 2298
rect 3300 2282 3354 2298
rect 2954 2218 3002 2282
rect 3066 2218 3082 2228
rect 3146 2218 3162 2228
rect 3226 2218 3242 2228
rect 3306 2218 3354 2282
rect 2954 2202 3354 2218
rect 3658 2522 4058 2538
rect 3658 2458 3706 2522
rect 3770 2484 3786 2522
rect 3850 2484 3866 2522
rect 3930 2484 3946 2522
rect 4010 2458 4058 2522
rect 3658 2442 3712 2458
rect 4004 2442 4058 2458
rect 3658 2378 3706 2442
rect 4010 2378 4058 2442
rect 3658 2362 3712 2378
rect 4004 2362 4058 2378
rect 3658 2298 3706 2362
rect 4010 2298 4058 2362
rect 3658 2282 3712 2298
rect 4004 2282 4058 2298
rect 3658 2218 3706 2282
rect 3770 2218 3786 2228
rect 3850 2218 3866 2228
rect 3930 2218 3946 2228
rect 4010 2218 4058 2282
rect 3658 2202 4058 2218
rect 4566 2492 4900 2584
rect 4566 2256 4620 2492
rect 4856 2256 4900 2492
rect 844 1878 1244 1880
rect 820 1862 1268 1878
rect 820 1798 890 1862
rect 954 1854 970 1862
rect 1034 1854 1050 1862
rect 1114 1854 1130 1862
rect 1194 1798 1268 1862
rect 820 1782 896 1798
rect 1188 1782 1268 1798
rect 820 1718 890 1782
rect 1194 1718 1268 1782
rect 820 1702 896 1718
rect 1188 1702 1268 1718
rect 820 1638 890 1702
rect 1194 1638 1268 1702
rect 820 1622 896 1638
rect 1188 1622 1268 1638
rect 658 1572 738 1580
rect 658 1508 666 1572
rect 730 1508 738 1572
rect 820 1558 890 1622
rect 954 1558 970 1598
rect 1034 1558 1050 1598
rect 1114 1558 1130 1598
rect 1194 1558 1268 1622
rect 820 1542 1268 1558
rect 1546 1862 1948 1878
rect 1546 1798 1594 1862
rect 1658 1854 1674 1862
rect 1738 1854 1754 1862
rect 1818 1854 1834 1862
rect 1898 1798 1948 1862
rect 1546 1782 1600 1798
rect 1892 1782 1948 1798
rect 1546 1718 1594 1782
rect 1898 1718 1948 1782
rect 1546 1702 1600 1718
rect 1892 1702 1948 1718
rect 1546 1638 1594 1702
rect 1898 1638 1948 1702
rect 1546 1622 1600 1638
rect 1892 1622 1948 1638
rect 1546 1558 1594 1622
rect 1658 1558 1674 1598
rect 1738 1558 1754 1598
rect 1818 1558 1834 1598
rect 1898 1558 1948 1622
rect 1546 1542 1948 1558
rect 2250 1862 2652 1878
rect 2250 1798 2298 1862
rect 2362 1854 2378 1862
rect 2442 1854 2458 1862
rect 2522 1854 2538 1862
rect 2602 1798 2652 1862
rect 2250 1782 2304 1798
rect 2596 1782 2652 1798
rect 2250 1718 2298 1782
rect 2602 1718 2652 1782
rect 2250 1702 2304 1718
rect 2596 1702 2652 1718
rect 2250 1638 2298 1702
rect 2602 1638 2652 1702
rect 2250 1622 2304 1638
rect 2596 1622 2652 1638
rect 2250 1558 2298 1622
rect 2362 1558 2378 1598
rect 2442 1558 2458 1598
rect 2522 1558 2538 1598
rect 2602 1558 2652 1622
rect 2250 1542 2652 1558
rect 2954 1862 3356 1878
rect 2954 1798 3002 1862
rect 3066 1854 3082 1862
rect 3146 1854 3162 1862
rect 3226 1854 3242 1862
rect 3306 1798 3356 1862
rect 2954 1782 3008 1798
rect 3300 1782 3356 1798
rect 2954 1718 3002 1782
rect 3306 1718 3356 1782
rect 2954 1702 3008 1718
rect 3300 1702 3356 1718
rect 2954 1638 3002 1702
rect 3306 1638 3356 1702
rect 2954 1622 3008 1638
rect 3300 1622 3356 1638
rect 2954 1558 3002 1622
rect 3066 1558 3082 1598
rect 3146 1558 3162 1598
rect 3226 1558 3242 1598
rect 3306 1558 3356 1622
rect 2954 1542 3356 1558
rect 3658 1862 4058 1878
rect 3658 1798 3706 1862
rect 3770 1854 3786 1862
rect 3850 1854 3866 1862
rect 3930 1854 3946 1862
rect 4010 1798 4058 1862
rect 3658 1782 3712 1798
rect 4004 1782 4058 1798
rect 3658 1718 3706 1782
rect 4010 1718 4058 1782
rect 3658 1702 3712 1718
rect 4004 1702 4058 1718
rect 3658 1638 3706 1702
rect 4010 1638 4058 1702
rect 3658 1622 3712 1638
rect 4004 1622 4058 1638
rect 3658 1558 3706 1622
rect 3770 1558 3786 1598
rect 3850 1558 3866 1598
rect 3930 1558 3946 1598
rect 4010 1558 4058 1622
rect 3658 1542 4058 1558
rect 658 1492 738 1508
rect 658 1428 666 1492
rect 730 1428 738 1492
rect 658 1420 738 1428
rect 4566 1496 4900 2256
rect 658 1340 724 1420
rect 658 1332 738 1340
rect 658 1268 666 1332
rect 730 1268 738 1332
rect 658 1252 738 1268
rect 658 1188 666 1252
rect 730 1188 738 1252
rect 4566 1260 4612 1496
rect 4848 1260 4900 1496
rect 658 1182 738 1188
rect 842 1198 1242 1214
rect 658 254 724 1182
rect 842 1134 890 1198
rect 954 1160 970 1198
rect 1034 1160 1050 1198
rect 1114 1160 1130 1198
rect 1194 1134 1242 1198
rect 842 1118 896 1134
rect 1188 1118 1242 1134
rect 842 1054 890 1118
rect 1194 1054 1242 1118
rect 842 1038 896 1054
rect 1188 1038 1242 1054
rect 842 974 890 1038
rect 1194 974 1242 1038
rect 842 958 896 974
rect 1188 958 1242 974
rect 842 894 890 958
rect 954 894 970 904
rect 1034 894 1050 904
rect 1114 894 1130 904
rect 1194 894 1242 958
rect 842 878 1242 894
rect 1546 1198 1946 1214
rect 1546 1134 1594 1198
rect 1658 1160 1674 1198
rect 1738 1160 1754 1198
rect 1818 1160 1834 1198
rect 1898 1134 1946 1198
rect 1546 1118 1600 1134
rect 1892 1118 1946 1134
rect 1546 1054 1594 1118
rect 1898 1054 1946 1118
rect 1546 1038 1600 1054
rect 1892 1038 1946 1054
rect 1546 974 1594 1038
rect 1898 974 1946 1038
rect 1546 958 1600 974
rect 1892 958 1946 974
rect 1546 894 1594 958
rect 1658 894 1674 904
rect 1738 894 1754 904
rect 1818 894 1834 904
rect 1898 894 1946 958
rect 1546 878 1946 894
rect 2954 1198 3354 1214
rect 2954 1134 3002 1198
rect 3066 1160 3082 1198
rect 3146 1160 3162 1198
rect 3226 1160 3242 1198
rect 3306 1134 3354 1198
rect 2954 1118 3008 1134
rect 3300 1118 3354 1134
rect 2954 1054 3002 1118
rect 3306 1054 3354 1118
rect 2954 1038 3008 1054
rect 3300 1038 3354 1054
rect 2954 974 3002 1038
rect 3306 974 3354 1038
rect 2954 958 3008 974
rect 3300 958 3354 974
rect 2954 894 3002 958
rect 3066 894 3082 904
rect 3146 894 3162 904
rect 3226 894 3242 904
rect 3306 894 3354 958
rect 2954 878 3354 894
rect 3658 1198 4058 1214
rect 3658 1134 3706 1198
rect 3770 1160 3786 1198
rect 3850 1160 3866 1198
rect 3930 1160 3946 1198
rect 4010 1134 4058 1198
rect 3658 1118 3712 1134
rect 4004 1118 4058 1134
rect 3658 1054 3706 1118
rect 4010 1054 4058 1118
rect 3658 1038 3712 1054
rect 4004 1038 4058 1054
rect 3658 974 3706 1038
rect 4010 974 4058 1038
rect 3658 958 3712 974
rect 4004 958 4058 974
rect 3658 894 3706 958
rect 3770 894 3786 904
rect 3850 894 3866 904
rect 3930 894 3946 904
rect 4010 894 4058 958
rect 3658 878 4058 894
rect 4566 1176 4900 1260
rect 4566 940 4606 1176
rect 4842 940 4900 1176
rect 4566 878 4900 940
rect 842 540 1244 556
rect 842 476 890 540
rect 954 530 970 540
rect 1034 530 1050 540
rect 1114 530 1130 540
rect 1194 476 1244 540
rect 842 460 896 476
rect 1188 460 1244 476
rect 842 396 890 460
rect 1194 396 1244 460
rect 842 380 896 396
rect 1188 380 1244 396
rect 842 316 890 380
rect 1194 316 1244 380
rect 842 300 896 316
rect 1188 300 1244 316
rect 658 246 738 254
rect 658 182 666 246
rect 730 182 738 246
rect 842 236 890 300
rect 954 236 970 274
rect 1034 236 1050 274
rect 1114 236 1130 274
rect 1194 236 1244 300
rect 842 220 1244 236
rect 1546 540 1948 556
rect 1546 476 1594 540
rect 1658 530 1674 540
rect 1738 530 1754 540
rect 1818 530 1834 540
rect 1898 476 1948 540
rect 1546 460 1600 476
rect 1892 460 1948 476
rect 1546 396 1594 460
rect 1898 396 1948 460
rect 1546 380 1600 396
rect 1892 380 1948 396
rect 1546 316 1594 380
rect 1898 316 1948 380
rect 1546 300 1600 316
rect 1892 300 1948 316
rect 1546 236 1594 300
rect 1658 236 1674 274
rect 1738 236 1754 274
rect 1818 236 1834 274
rect 1898 236 1948 300
rect 1546 220 1948 236
rect 2954 540 3356 556
rect 2954 476 3002 540
rect 3066 530 3082 540
rect 3146 530 3162 540
rect 3226 530 3242 540
rect 3306 476 3356 540
rect 2954 460 3008 476
rect 3300 460 3356 476
rect 2954 396 3002 460
rect 3306 396 3356 460
rect 2954 380 3008 396
rect 3300 380 3356 396
rect 2954 316 3002 380
rect 3306 316 3356 380
rect 2954 300 3008 316
rect 3300 300 3356 316
rect 2954 236 3002 300
rect 3066 236 3082 274
rect 3146 236 3162 274
rect 3226 236 3242 274
rect 3306 236 3356 300
rect 2954 220 3356 236
rect 3604 540 4058 556
rect 3604 476 3706 540
rect 3770 530 3786 540
rect 3850 530 3866 540
rect 3930 530 3946 540
rect 4010 476 4058 540
rect 3604 460 3712 476
rect 4004 460 4058 476
rect 3604 396 3706 460
rect 4010 396 4058 460
rect 3604 380 3712 396
rect 4004 380 4058 396
rect 3604 316 3706 380
rect 4010 316 4058 380
rect 3604 300 3712 316
rect 4004 300 4058 316
rect 3604 236 3706 300
rect 3770 236 3786 274
rect 3850 236 3866 274
rect 3930 236 3946 274
rect 4010 236 4058 300
rect 3604 220 4058 236
rect 658 166 738 182
rect 658 102 666 166
rect 730 102 738 166
rect 658 94 738 102
rect -2 -100 334 -56
rect -2 -128 512 -100
rect -2 -158 244 -128
rect 308 -158 370 -128
rect 434 -158 512 -128
rect -2 -394 56 -158
rect 456 -394 512 -158
rect -2 -402 512 -394
rect -2 -466 244 -402
rect 308 -466 370 -402
rect 434 -466 512 -402
rect -2 -480 512 -466
rect -2 -716 54 -480
rect 454 -716 512 -480
rect -2 -744 244 -716
rect 308 -744 370 -716
rect 434 -744 512 -716
rect -2 -772 512 -744
rect 800 -128 1098 -100
rect 800 -158 852 -128
rect 916 -158 978 -128
rect 1042 -158 1098 -128
rect 800 -394 828 -158
rect 1064 -394 1098 -158
rect 800 -402 1098 -394
rect 800 -466 852 -402
rect 916 -466 978 -402
rect 1042 -466 1098 -402
rect 800 -480 1098 -466
rect 800 -716 826 -480
rect 1062 -716 1098 -480
rect 800 -744 852 -716
rect 916 -744 978 -716
rect 1042 -744 1098 -716
rect 800 -772 1098 -744
rect 1650 -128 1948 -100
rect 1650 -158 1702 -128
rect 1766 -158 1828 -128
rect 1892 -158 1948 -128
rect 1650 -394 1678 -158
rect 1914 -394 1948 -158
rect 1650 -402 1948 -394
rect 1650 -466 1702 -402
rect 1766 -466 1828 -402
rect 1892 -466 1948 -402
rect 1650 -480 1948 -466
rect 1650 -716 1676 -480
rect 1912 -716 1948 -480
rect 1650 -744 1702 -716
rect 1766 -744 1828 -716
rect 1892 -744 1948 -716
rect 1650 -772 1948 -744
rect 2294 -128 2640 -100
rect 2294 -158 2372 -128
rect 2436 -158 2498 -128
rect 2562 -158 2640 -128
rect 2294 -394 2348 -158
rect 2584 -394 2640 -158
rect 2294 -402 2640 -394
rect 2294 -466 2372 -402
rect 2436 -466 2498 -402
rect 2562 -466 2640 -402
rect 2294 -480 2640 -466
rect 2294 -716 2346 -480
rect 2582 -716 2640 -480
rect 2294 -744 2372 -716
rect 2436 -744 2498 -716
rect 2562 -744 2640 -716
rect 2294 -772 2640 -744
rect 2834 -128 3132 -100
rect 2834 -158 2886 -128
rect 2950 -158 3012 -128
rect 3076 -158 3132 -128
rect 2834 -394 2862 -158
rect 3098 -394 3132 -158
rect 2834 -402 3132 -394
rect 2834 -466 2886 -402
rect 2950 -466 3012 -402
rect 3076 -466 3132 -402
rect 2834 -480 3132 -466
rect 2834 -716 2860 -480
rect 3096 -716 3132 -480
rect 2834 -744 2886 -716
rect 2950 -744 3012 -716
rect 3076 -744 3132 -716
rect 2834 -772 3132 -744
rect 3654 -128 3952 -100
rect 3654 -158 3706 -128
rect 3770 -158 3832 -128
rect 3896 -158 3952 -128
rect 3654 -394 3682 -158
rect 3918 -394 3952 -158
rect 3654 -402 3952 -394
rect 3654 -466 3706 -402
rect 3770 -466 3832 -402
rect 3896 -466 3952 -402
rect 3654 -480 3952 -466
rect 3654 -716 3680 -480
rect 3916 -716 3952 -480
rect 3654 -744 3706 -716
rect 3770 -744 3832 -716
rect 3896 -744 3952 -716
rect 3654 -772 3952 -744
rect 4386 -128 4732 -100
rect 4386 -158 4464 -128
rect 4528 -158 4590 -128
rect 4654 -158 4732 -128
rect 4386 -394 4440 -158
rect 4676 -394 4732 -158
rect 4386 -402 4732 -394
rect 4386 -466 4464 -402
rect 4528 -466 4590 -402
rect 4654 -466 4732 -402
rect 4386 -480 4732 -466
rect 4386 -716 4438 -480
rect 4674 -716 4732 -480
rect 4386 -744 4464 -716
rect 4528 -744 4590 -716
rect 4654 -744 4732 -716
rect 4386 -772 4732 -744
<< via4 >>
rect 574 2906 810 3142
rect 2088 2908 2324 3144
rect 2418 2908 2654 3144
rect 48 1596 284 1832
rect 46 1252 282 1488
rect 52 286 288 522
rect 46 -56 282 180
rect 896 2458 954 2484
rect 954 2458 970 2484
rect 970 2458 1034 2484
rect 1034 2458 1050 2484
rect 1050 2458 1114 2484
rect 1114 2458 1130 2484
rect 1130 2458 1188 2484
rect 896 2442 1188 2458
rect 896 2378 954 2442
rect 954 2378 970 2442
rect 970 2378 1034 2442
rect 1034 2378 1050 2442
rect 1050 2378 1114 2442
rect 1114 2378 1130 2442
rect 1130 2378 1188 2442
rect 896 2362 1188 2378
rect 896 2298 954 2362
rect 954 2298 970 2362
rect 970 2298 1034 2362
rect 1034 2298 1050 2362
rect 1050 2298 1114 2362
rect 1114 2298 1130 2362
rect 1130 2298 1188 2362
rect 896 2282 1188 2298
rect 896 2228 954 2282
rect 954 2228 970 2282
rect 970 2228 1034 2282
rect 1034 2228 1050 2282
rect 1050 2228 1114 2282
rect 1114 2228 1130 2282
rect 1130 2228 1188 2282
rect 1600 2458 1658 2484
rect 1658 2458 1674 2484
rect 1674 2458 1738 2484
rect 1738 2458 1754 2484
rect 1754 2458 1818 2484
rect 1818 2458 1834 2484
rect 1834 2458 1892 2484
rect 1600 2442 1892 2458
rect 1600 2378 1658 2442
rect 1658 2378 1674 2442
rect 1674 2378 1738 2442
rect 1738 2378 1754 2442
rect 1754 2378 1818 2442
rect 1818 2378 1834 2442
rect 1834 2378 1892 2442
rect 1600 2362 1892 2378
rect 1600 2298 1658 2362
rect 1658 2298 1674 2362
rect 1674 2298 1738 2362
rect 1738 2298 1754 2362
rect 1754 2298 1818 2362
rect 1818 2298 1834 2362
rect 1834 2298 1892 2362
rect 1600 2282 1892 2298
rect 1600 2228 1658 2282
rect 1658 2228 1674 2282
rect 1674 2228 1738 2282
rect 1738 2228 1754 2282
rect 1754 2228 1818 2282
rect 1818 2228 1834 2282
rect 1834 2228 1892 2282
rect 4612 2584 4848 2820
rect 3008 2458 3066 2484
rect 3066 2458 3082 2484
rect 3082 2458 3146 2484
rect 3146 2458 3162 2484
rect 3162 2458 3226 2484
rect 3226 2458 3242 2484
rect 3242 2458 3300 2484
rect 3008 2442 3300 2458
rect 3008 2378 3066 2442
rect 3066 2378 3082 2442
rect 3082 2378 3146 2442
rect 3146 2378 3162 2442
rect 3162 2378 3226 2442
rect 3226 2378 3242 2442
rect 3242 2378 3300 2442
rect 3008 2362 3300 2378
rect 3008 2298 3066 2362
rect 3066 2298 3082 2362
rect 3082 2298 3146 2362
rect 3146 2298 3162 2362
rect 3162 2298 3226 2362
rect 3226 2298 3242 2362
rect 3242 2298 3300 2362
rect 3008 2282 3300 2298
rect 3008 2228 3066 2282
rect 3066 2228 3082 2282
rect 3082 2228 3146 2282
rect 3146 2228 3162 2282
rect 3162 2228 3226 2282
rect 3226 2228 3242 2282
rect 3242 2228 3300 2282
rect 3712 2458 3770 2484
rect 3770 2458 3786 2484
rect 3786 2458 3850 2484
rect 3850 2458 3866 2484
rect 3866 2458 3930 2484
rect 3930 2458 3946 2484
rect 3946 2458 4004 2484
rect 3712 2442 4004 2458
rect 3712 2378 3770 2442
rect 3770 2378 3786 2442
rect 3786 2378 3850 2442
rect 3850 2378 3866 2442
rect 3866 2378 3930 2442
rect 3930 2378 3946 2442
rect 3946 2378 4004 2442
rect 3712 2362 4004 2378
rect 3712 2298 3770 2362
rect 3770 2298 3786 2362
rect 3786 2298 3850 2362
rect 3850 2298 3866 2362
rect 3866 2298 3930 2362
rect 3930 2298 3946 2362
rect 3946 2298 4004 2362
rect 3712 2282 4004 2298
rect 3712 2228 3770 2282
rect 3770 2228 3786 2282
rect 3786 2228 3850 2282
rect 3850 2228 3866 2282
rect 3866 2228 3930 2282
rect 3930 2228 3946 2282
rect 3946 2228 4004 2282
rect 4620 2256 4856 2492
rect 896 1798 954 1854
rect 954 1798 970 1854
rect 970 1798 1034 1854
rect 1034 1798 1050 1854
rect 1050 1798 1114 1854
rect 1114 1798 1130 1854
rect 1130 1798 1188 1854
rect 896 1782 1188 1798
rect 896 1718 954 1782
rect 954 1718 970 1782
rect 970 1718 1034 1782
rect 1034 1718 1050 1782
rect 1050 1718 1114 1782
rect 1114 1718 1130 1782
rect 1130 1718 1188 1782
rect 896 1702 1188 1718
rect 896 1638 954 1702
rect 954 1638 970 1702
rect 970 1638 1034 1702
rect 1034 1638 1050 1702
rect 1050 1638 1114 1702
rect 1114 1638 1130 1702
rect 1130 1638 1188 1702
rect 896 1622 1188 1638
rect 896 1598 954 1622
rect 954 1598 970 1622
rect 970 1598 1034 1622
rect 1034 1598 1050 1622
rect 1050 1598 1114 1622
rect 1114 1598 1130 1622
rect 1130 1598 1188 1622
rect 1600 1798 1658 1854
rect 1658 1798 1674 1854
rect 1674 1798 1738 1854
rect 1738 1798 1754 1854
rect 1754 1798 1818 1854
rect 1818 1798 1834 1854
rect 1834 1798 1892 1854
rect 1600 1782 1892 1798
rect 1600 1718 1658 1782
rect 1658 1718 1674 1782
rect 1674 1718 1738 1782
rect 1738 1718 1754 1782
rect 1754 1718 1818 1782
rect 1818 1718 1834 1782
rect 1834 1718 1892 1782
rect 1600 1702 1892 1718
rect 1600 1638 1658 1702
rect 1658 1638 1674 1702
rect 1674 1638 1738 1702
rect 1738 1638 1754 1702
rect 1754 1638 1818 1702
rect 1818 1638 1834 1702
rect 1834 1638 1892 1702
rect 1600 1622 1892 1638
rect 1600 1598 1658 1622
rect 1658 1598 1674 1622
rect 1674 1598 1738 1622
rect 1738 1598 1754 1622
rect 1754 1598 1818 1622
rect 1818 1598 1834 1622
rect 1834 1598 1892 1622
rect 2304 1798 2362 1854
rect 2362 1798 2378 1854
rect 2378 1798 2442 1854
rect 2442 1798 2458 1854
rect 2458 1798 2522 1854
rect 2522 1798 2538 1854
rect 2538 1798 2596 1854
rect 2304 1782 2596 1798
rect 2304 1718 2362 1782
rect 2362 1718 2378 1782
rect 2378 1718 2442 1782
rect 2442 1718 2458 1782
rect 2458 1718 2522 1782
rect 2522 1718 2538 1782
rect 2538 1718 2596 1782
rect 2304 1702 2596 1718
rect 2304 1638 2362 1702
rect 2362 1638 2378 1702
rect 2378 1638 2442 1702
rect 2442 1638 2458 1702
rect 2458 1638 2522 1702
rect 2522 1638 2538 1702
rect 2538 1638 2596 1702
rect 2304 1622 2596 1638
rect 2304 1598 2362 1622
rect 2362 1598 2378 1622
rect 2378 1598 2442 1622
rect 2442 1598 2458 1622
rect 2458 1598 2522 1622
rect 2522 1598 2538 1622
rect 2538 1598 2596 1622
rect 3008 1798 3066 1854
rect 3066 1798 3082 1854
rect 3082 1798 3146 1854
rect 3146 1798 3162 1854
rect 3162 1798 3226 1854
rect 3226 1798 3242 1854
rect 3242 1798 3300 1854
rect 3008 1782 3300 1798
rect 3008 1718 3066 1782
rect 3066 1718 3082 1782
rect 3082 1718 3146 1782
rect 3146 1718 3162 1782
rect 3162 1718 3226 1782
rect 3226 1718 3242 1782
rect 3242 1718 3300 1782
rect 3008 1702 3300 1718
rect 3008 1638 3066 1702
rect 3066 1638 3082 1702
rect 3082 1638 3146 1702
rect 3146 1638 3162 1702
rect 3162 1638 3226 1702
rect 3226 1638 3242 1702
rect 3242 1638 3300 1702
rect 3008 1622 3300 1638
rect 3008 1598 3066 1622
rect 3066 1598 3082 1622
rect 3082 1598 3146 1622
rect 3146 1598 3162 1622
rect 3162 1598 3226 1622
rect 3226 1598 3242 1622
rect 3242 1598 3300 1622
rect 3712 1798 3770 1854
rect 3770 1798 3786 1854
rect 3786 1798 3850 1854
rect 3850 1798 3866 1854
rect 3866 1798 3930 1854
rect 3930 1798 3946 1854
rect 3946 1798 4004 1854
rect 3712 1782 4004 1798
rect 3712 1718 3770 1782
rect 3770 1718 3786 1782
rect 3786 1718 3850 1782
rect 3850 1718 3866 1782
rect 3866 1718 3930 1782
rect 3930 1718 3946 1782
rect 3946 1718 4004 1782
rect 3712 1702 4004 1718
rect 3712 1638 3770 1702
rect 3770 1638 3786 1702
rect 3786 1638 3850 1702
rect 3850 1638 3866 1702
rect 3866 1638 3930 1702
rect 3930 1638 3946 1702
rect 3946 1638 4004 1702
rect 3712 1622 4004 1638
rect 3712 1598 3770 1622
rect 3770 1598 3786 1622
rect 3786 1598 3850 1622
rect 3850 1598 3866 1622
rect 3866 1598 3930 1622
rect 3930 1598 3946 1622
rect 3946 1598 4004 1622
rect 4612 1260 4848 1496
rect 896 1134 954 1160
rect 954 1134 970 1160
rect 970 1134 1034 1160
rect 1034 1134 1050 1160
rect 1050 1134 1114 1160
rect 1114 1134 1130 1160
rect 1130 1134 1188 1160
rect 896 1118 1188 1134
rect 896 1054 954 1118
rect 954 1054 970 1118
rect 970 1054 1034 1118
rect 1034 1054 1050 1118
rect 1050 1054 1114 1118
rect 1114 1054 1130 1118
rect 1130 1054 1188 1118
rect 896 1038 1188 1054
rect 896 974 954 1038
rect 954 974 970 1038
rect 970 974 1034 1038
rect 1034 974 1050 1038
rect 1050 974 1114 1038
rect 1114 974 1130 1038
rect 1130 974 1188 1038
rect 896 958 1188 974
rect 896 904 954 958
rect 954 904 970 958
rect 970 904 1034 958
rect 1034 904 1050 958
rect 1050 904 1114 958
rect 1114 904 1130 958
rect 1130 904 1188 958
rect 1600 1134 1658 1160
rect 1658 1134 1674 1160
rect 1674 1134 1738 1160
rect 1738 1134 1754 1160
rect 1754 1134 1818 1160
rect 1818 1134 1834 1160
rect 1834 1134 1892 1160
rect 1600 1118 1892 1134
rect 1600 1054 1658 1118
rect 1658 1054 1674 1118
rect 1674 1054 1738 1118
rect 1738 1054 1754 1118
rect 1754 1054 1818 1118
rect 1818 1054 1834 1118
rect 1834 1054 1892 1118
rect 1600 1038 1892 1054
rect 1600 974 1658 1038
rect 1658 974 1674 1038
rect 1674 974 1738 1038
rect 1738 974 1754 1038
rect 1754 974 1818 1038
rect 1818 974 1834 1038
rect 1834 974 1892 1038
rect 1600 958 1892 974
rect 1600 904 1658 958
rect 1658 904 1674 958
rect 1674 904 1738 958
rect 1738 904 1754 958
rect 1754 904 1818 958
rect 1818 904 1834 958
rect 1834 904 1892 958
rect 3008 1134 3066 1160
rect 3066 1134 3082 1160
rect 3082 1134 3146 1160
rect 3146 1134 3162 1160
rect 3162 1134 3226 1160
rect 3226 1134 3242 1160
rect 3242 1134 3300 1160
rect 3008 1118 3300 1134
rect 3008 1054 3066 1118
rect 3066 1054 3082 1118
rect 3082 1054 3146 1118
rect 3146 1054 3162 1118
rect 3162 1054 3226 1118
rect 3226 1054 3242 1118
rect 3242 1054 3300 1118
rect 3008 1038 3300 1054
rect 3008 974 3066 1038
rect 3066 974 3082 1038
rect 3082 974 3146 1038
rect 3146 974 3162 1038
rect 3162 974 3226 1038
rect 3226 974 3242 1038
rect 3242 974 3300 1038
rect 3008 958 3300 974
rect 3008 904 3066 958
rect 3066 904 3082 958
rect 3082 904 3146 958
rect 3146 904 3162 958
rect 3162 904 3226 958
rect 3226 904 3242 958
rect 3242 904 3300 958
rect 3712 1134 3770 1160
rect 3770 1134 3786 1160
rect 3786 1134 3850 1160
rect 3850 1134 3866 1160
rect 3866 1134 3930 1160
rect 3930 1134 3946 1160
rect 3946 1134 4004 1160
rect 3712 1118 4004 1134
rect 3712 1054 3770 1118
rect 3770 1054 3786 1118
rect 3786 1054 3850 1118
rect 3850 1054 3866 1118
rect 3866 1054 3930 1118
rect 3930 1054 3946 1118
rect 3946 1054 4004 1118
rect 3712 1038 4004 1054
rect 3712 974 3770 1038
rect 3770 974 3786 1038
rect 3786 974 3850 1038
rect 3850 974 3866 1038
rect 3866 974 3930 1038
rect 3930 974 3946 1038
rect 3946 974 4004 1038
rect 3712 958 4004 974
rect 3712 904 3770 958
rect 3770 904 3786 958
rect 3786 904 3850 958
rect 3850 904 3866 958
rect 3866 904 3930 958
rect 3930 904 3946 958
rect 3946 904 4004 958
rect 4606 940 4842 1176
rect 896 476 954 530
rect 954 476 970 530
rect 970 476 1034 530
rect 1034 476 1050 530
rect 1050 476 1114 530
rect 1114 476 1130 530
rect 1130 476 1188 530
rect 896 460 1188 476
rect 896 396 954 460
rect 954 396 970 460
rect 970 396 1034 460
rect 1034 396 1050 460
rect 1050 396 1114 460
rect 1114 396 1130 460
rect 1130 396 1188 460
rect 896 380 1188 396
rect 896 316 954 380
rect 954 316 970 380
rect 970 316 1034 380
rect 1034 316 1050 380
rect 1050 316 1114 380
rect 1114 316 1130 380
rect 1130 316 1188 380
rect 896 300 1188 316
rect 896 274 954 300
rect 954 274 970 300
rect 970 274 1034 300
rect 1034 274 1050 300
rect 1050 274 1114 300
rect 1114 274 1130 300
rect 1130 274 1188 300
rect 1600 476 1658 530
rect 1658 476 1674 530
rect 1674 476 1738 530
rect 1738 476 1754 530
rect 1754 476 1818 530
rect 1818 476 1834 530
rect 1834 476 1892 530
rect 1600 460 1892 476
rect 1600 396 1658 460
rect 1658 396 1674 460
rect 1674 396 1738 460
rect 1738 396 1754 460
rect 1754 396 1818 460
rect 1818 396 1834 460
rect 1834 396 1892 460
rect 1600 380 1892 396
rect 1600 316 1658 380
rect 1658 316 1674 380
rect 1674 316 1738 380
rect 1738 316 1754 380
rect 1754 316 1818 380
rect 1818 316 1834 380
rect 1834 316 1892 380
rect 1600 300 1892 316
rect 1600 274 1658 300
rect 1658 274 1674 300
rect 1674 274 1738 300
rect 1738 274 1754 300
rect 1754 274 1818 300
rect 1818 274 1834 300
rect 1834 274 1892 300
rect 3008 476 3066 530
rect 3066 476 3082 530
rect 3082 476 3146 530
rect 3146 476 3162 530
rect 3162 476 3226 530
rect 3226 476 3242 530
rect 3242 476 3300 530
rect 3008 460 3300 476
rect 3008 396 3066 460
rect 3066 396 3082 460
rect 3082 396 3146 460
rect 3146 396 3162 460
rect 3162 396 3226 460
rect 3226 396 3242 460
rect 3242 396 3300 460
rect 3008 380 3300 396
rect 3008 316 3066 380
rect 3066 316 3082 380
rect 3082 316 3146 380
rect 3146 316 3162 380
rect 3162 316 3226 380
rect 3226 316 3242 380
rect 3242 316 3300 380
rect 3008 300 3300 316
rect 3008 274 3066 300
rect 3066 274 3082 300
rect 3082 274 3146 300
rect 3146 274 3162 300
rect 3162 274 3226 300
rect 3226 274 3242 300
rect 3242 274 3300 300
rect 3712 476 3770 530
rect 3770 476 3786 530
rect 3786 476 3850 530
rect 3850 476 3866 530
rect 3866 476 3930 530
rect 3930 476 3946 530
rect 3946 476 4004 530
rect 3712 460 4004 476
rect 3712 396 3770 460
rect 3770 396 3786 460
rect 3786 396 3850 460
rect 3850 396 3866 460
rect 3866 396 3930 460
rect 3930 396 3946 460
rect 3946 396 4004 460
rect 3712 380 4004 396
rect 3712 316 3770 380
rect 3770 316 3786 380
rect 3786 316 3850 380
rect 3850 316 3866 380
rect 3866 316 3930 380
rect 3930 316 3946 380
rect 3946 316 4004 380
rect 3712 300 4004 316
rect 3712 274 3770 300
rect 3770 274 3786 300
rect 3786 274 3850 300
rect 3850 274 3866 300
rect 3866 274 3930 300
rect 3930 274 3946 300
rect 3946 274 4004 300
rect 56 -192 244 -158
rect 244 -192 308 -158
rect 308 -192 370 -158
rect 370 -192 434 -158
rect 434 -192 456 -158
rect 56 -232 456 -192
rect 56 -296 244 -232
rect 244 -296 308 -232
rect 308 -296 370 -232
rect 370 -296 434 -232
rect 434 -296 456 -232
rect 56 -316 456 -296
rect 56 -380 244 -316
rect 244 -380 308 -316
rect 308 -380 370 -316
rect 370 -380 434 -316
rect 434 -380 456 -316
rect 56 -394 456 -380
rect 54 -496 454 -480
rect 54 -560 244 -496
rect 244 -560 308 -496
rect 308 -560 370 -496
rect 370 -560 434 -496
rect 434 -560 454 -496
rect 54 -596 454 -560
rect 54 -660 244 -596
rect 244 -660 308 -596
rect 308 -660 370 -596
rect 370 -660 434 -596
rect 434 -660 454 -596
rect 54 -680 454 -660
rect 54 -716 244 -680
rect 244 -716 308 -680
rect 308 -716 370 -680
rect 370 -716 434 -680
rect 434 -716 454 -680
rect 828 -192 852 -158
rect 852 -192 916 -158
rect 916 -192 978 -158
rect 978 -192 1042 -158
rect 1042 -192 1064 -158
rect 828 -232 1064 -192
rect 828 -296 852 -232
rect 852 -296 916 -232
rect 916 -296 978 -232
rect 978 -296 1042 -232
rect 1042 -296 1064 -232
rect 828 -316 1064 -296
rect 828 -380 852 -316
rect 852 -380 916 -316
rect 916 -380 978 -316
rect 978 -380 1042 -316
rect 1042 -380 1064 -316
rect 828 -394 1064 -380
rect 826 -496 1062 -480
rect 826 -560 852 -496
rect 852 -560 916 -496
rect 916 -560 978 -496
rect 978 -560 1042 -496
rect 1042 -560 1062 -496
rect 826 -596 1062 -560
rect 826 -660 852 -596
rect 852 -660 916 -596
rect 916 -660 978 -596
rect 978 -660 1042 -596
rect 1042 -660 1062 -596
rect 826 -680 1062 -660
rect 826 -716 852 -680
rect 852 -716 916 -680
rect 916 -716 978 -680
rect 978 -716 1042 -680
rect 1042 -716 1062 -680
rect 1678 -192 1702 -158
rect 1702 -192 1766 -158
rect 1766 -192 1828 -158
rect 1828 -192 1892 -158
rect 1892 -192 1914 -158
rect 1678 -232 1914 -192
rect 1678 -296 1702 -232
rect 1702 -296 1766 -232
rect 1766 -296 1828 -232
rect 1828 -296 1892 -232
rect 1892 -296 1914 -232
rect 1678 -316 1914 -296
rect 1678 -380 1702 -316
rect 1702 -380 1766 -316
rect 1766 -380 1828 -316
rect 1828 -380 1892 -316
rect 1892 -380 1914 -316
rect 1678 -394 1914 -380
rect 1676 -496 1912 -480
rect 1676 -560 1702 -496
rect 1702 -560 1766 -496
rect 1766 -560 1828 -496
rect 1828 -560 1892 -496
rect 1892 -560 1912 -496
rect 1676 -596 1912 -560
rect 1676 -660 1702 -596
rect 1702 -660 1766 -596
rect 1766 -660 1828 -596
rect 1828 -660 1892 -596
rect 1892 -660 1912 -596
rect 1676 -680 1912 -660
rect 1676 -716 1702 -680
rect 1702 -716 1766 -680
rect 1766 -716 1828 -680
rect 1828 -716 1892 -680
rect 1892 -716 1912 -680
rect 2348 -192 2372 -158
rect 2372 -192 2436 -158
rect 2436 -192 2498 -158
rect 2498 -192 2562 -158
rect 2562 -192 2584 -158
rect 2348 -232 2584 -192
rect 2348 -296 2372 -232
rect 2372 -296 2436 -232
rect 2436 -296 2498 -232
rect 2498 -296 2562 -232
rect 2562 -296 2584 -232
rect 2348 -316 2584 -296
rect 2348 -380 2372 -316
rect 2372 -380 2436 -316
rect 2436 -380 2498 -316
rect 2498 -380 2562 -316
rect 2562 -380 2584 -316
rect 2348 -394 2584 -380
rect 2346 -496 2582 -480
rect 2346 -560 2372 -496
rect 2372 -560 2436 -496
rect 2436 -560 2498 -496
rect 2498 -560 2562 -496
rect 2562 -560 2582 -496
rect 2346 -596 2582 -560
rect 2346 -660 2372 -596
rect 2372 -660 2436 -596
rect 2436 -660 2498 -596
rect 2498 -660 2562 -596
rect 2562 -660 2582 -596
rect 2346 -680 2582 -660
rect 2346 -716 2372 -680
rect 2372 -716 2436 -680
rect 2436 -716 2498 -680
rect 2498 -716 2562 -680
rect 2562 -716 2582 -680
rect 2862 -192 2886 -158
rect 2886 -192 2950 -158
rect 2950 -192 3012 -158
rect 3012 -192 3076 -158
rect 3076 -192 3098 -158
rect 2862 -232 3098 -192
rect 2862 -296 2886 -232
rect 2886 -296 2950 -232
rect 2950 -296 3012 -232
rect 3012 -296 3076 -232
rect 3076 -296 3098 -232
rect 2862 -316 3098 -296
rect 2862 -380 2886 -316
rect 2886 -380 2950 -316
rect 2950 -380 3012 -316
rect 3012 -380 3076 -316
rect 3076 -380 3098 -316
rect 2862 -394 3098 -380
rect 2860 -496 3096 -480
rect 2860 -560 2886 -496
rect 2886 -560 2950 -496
rect 2950 -560 3012 -496
rect 3012 -560 3076 -496
rect 3076 -560 3096 -496
rect 2860 -596 3096 -560
rect 2860 -660 2886 -596
rect 2886 -660 2950 -596
rect 2950 -660 3012 -596
rect 3012 -660 3076 -596
rect 3076 -660 3096 -596
rect 2860 -680 3096 -660
rect 2860 -716 2886 -680
rect 2886 -716 2950 -680
rect 2950 -716 3012 -680
rect 3012 -716 3076 -680
rect 3076 -716 3096 -680
rect 3682 -192 3706 -158
rect 3706 -192 3770 -158
rect 3770 -192 3832 -158
rect 3832 -192 3896 -158
rect 3896 -192 3918 -158
rect 3682 -232 3918 -192
rect 3682 -296 3706 -232
rect 3706 -296 3770 -232
rect 3770 -296 3832 -232
rect 3832 -296 3896 -232
rect 3896 -296 3918 -232
rect 3682 -316 3918 -296
rect 3682 -380 3706 -316
rect 3706 -380 3770 -316
rect 3770 -380 3832 -316
rect 3832 -380 3896 -316
rect 3896 -380 3918 -316
rect 3682 -394 3918 -380
rect 3680 -496 3916 -480
rect 3680 -560 3706 -496
rect 3706 -560 3770 -496
rect 3770 -560 3832 -496
rect 3832 -560 3896 -496
rect 3896 -560 3916 -496
rect 3680 -596 3916 -560
rect 3680 -660 3706 -596
rect 3706 -660 3770 -596
rect 3770 -660 3832 -596
rect 3832 -660 3896 -596
rect 3896 -660 3916 -596
rect 3680 -680 3916 -660
rect 3680 -716 3706 -680
rect 3706 -716 3770 -680
rect 3770 -716 3832 -680
rect 3832 -716 3896 -680
rect 3896 -716 3916 -680
rect 4440 -192 4464 -158
rect 4464 -192 4528 -158
rect 4528 -192 4590 -158
rect 4590 -192 4654 -158
rect 4654 -192 4676 -158
rect 4440 -232 4676 -192
rect 4440 -296 4464 -232
rect 4464 -296 4528 -232
rect 4528 -296 4590 -232
rect 4590 -296 4654 -232
rect 4654 -296 4676 -232
rect 4440 -316 4676 -296
rect 4440 -380 4464 -316
rect 4464 -380 4528 -316
rect 4528 -380 4590 -316
rect 4590 -380 4654 -316
rect 4654 -380 4676 -316
rect 4440 -394 4676 -380
rect 4438 -496 4674 -480
rect 4438 -560 4464 -496
rect 4464 -560 4528 -496
rect 4528 -560 4590 -496
rect 4590 -560 4654 -496
rect 4654 -560 4674 -496
rect 4438 -596 4674 -560
rect 4438 -660 4464 -596
rect 4464 -660 4528 -596
rect 4528 -660 4590 -596
rect 4590 -660 4654 -596
rect 4654 -660 4674 -596
rect 4438 -680 4674 -660
rect 4438 -716 4464 -680
rect 4464 -716 4528 -680
rect 4528 -716 4590 -680
rect 4590 -716 4654 -680
rect 4654 -716 4674 -680
<< metal5 >>
rect 0 3144 2704 3194
rect 0 3142 2088 3144
rect 0 2906 574 3142
rect 810 2908 2088 3142
rect 2324 2908 2418 3144
rect 2654 2908 2704 3144
rect 810 2906 2704 2908
rect 0 2858 2704 2906
rect 4566 2820 4900 2874
rect 4566 2584 4612 2820
rect 4848 2584 4900 2820
rect 4566 2538 4900 2584
rect 704 2492 4900 2538
rect 704 2484 4620 2492
rect 704 2228 896 2484
rect 1188 2228 1600 2484
rect 1892 2228 3008 2484
rect 3300 2228 3712 2484
rect 4004 2256 4620 2484
rect 4856 2256 4900 2492
rect 4004 2228 4900 2256
rect 704 2202 4900 2228
rect 0 1854 4196 1878
rect 0 1832 896 1854
rect 0 1596 48 1832
rect 284 1598 896 1832
rect 1188 1598 1600 1854
rect 1892 1598 2304 1854
rect 2596 1598 3008 1854
rect 3300 1598 3712 1854
rect 4004 1598 4196 1854
rect 284 1596 4196 1598
rect 0 1544 4196 1596
rect 0 1488 334 1544
rect 704 1542 4196 1544
rect 0 1252 46 1488
rect 282 1252 334 1488
rect 0 1208 334 1252
rect 4566 1496 4900 1550
rect 4566 1260 4612 1496
rect 4848 1260 4900 1496
rect 4566 1214 4900 1260
rect 704 1176 4900 1214
rect 704 1160 4606 1176
rect 704 904 896 1160
rect 1188 904 1600 1160
rect 1892 904 3008 1160
rect 3300 904 3712 1160
rect 4004 940 4606 1160
rect 4842 940 4900 1176
rect 4004 904 4900 940
rect 704 878 4900 904
rect 2 530 4196 556
rect 2 522 896 530
rect 2 286 52 522
rect 288 286 896 522
rect 2 274 896 286
rect 1188 274 1600 530
rect 1892 274 3008 530
rect 3300 274 3712 530
rect 4004 274 4196 530
rect 2 220 4196 274
rect -2 180 334 220
rect -2 -56 46 180
rect 282 -56 334 180
rect -2 -100 334 -56
rect -2 -158 4900 -100
rect -2 -394 56 -158
rect 456 -394 828 -158
rect 1064 -394 1678 -158
rect 1914 -394 2348 -158
rect 2584 -394 2862 -158
rect 3098 -394 3682 -158
rect 3918 -394 4440 -158
rect 4676 -394 4900 -158
rect -2 -480 4900 -394
rect -2 -716 54 -480
rect 454 -716 826 -480
rect 1062 -716 1676 -480
rect 1912 -716 2346 -480
rect 2582 -716 2860 -480
rect 3096 -716 3680 -480
rect 3916 -716 4438 -480
rect 4674 -716 4900 -480
rect -2 -772 4900 -716
use buffer_mirror_base  buffer_mirror_base_0
timestamp 1654373441
transform 1 0 746 0 1 128
box -753 -8 4154 2510
<< end >>
