magic
tech sky130B
timestamp 1654639816
<< metal1 >>
rect 74 1259 176 1263
rect 74 1233 77 1259
rect 103 1233 112 1259
rect 138 1233 147 1259
rect 173 1233 176 1259
rect 74 1229 176 1233
rect 271 1259 373 1263
rect 271 1233 274 1259
rect 300 1233 309 1259
rect 335 1233 344 1259
rect 370 1233 373 1259
rect 271 1229 373 1233
rect 468 1259 570 1263
rect 468 1233 471 1259
rect 497 1233 506 1259
rect 532 1233 541 1259
rect 567 1233 570 1259
rect 468 1229 570 1233
rect 665 1259 767 1263
rect 665 1233 668 1259
rect 694 1233 703 1259
rect 729 1233 738 1259
rect 764 1233 767 1259
rect 665 1229 767 1233
rect 862 1259 964 1263
rect 862 1233 865 1259
rect 891 1233 900 1259
rect 926 1233 935 1259
rect 961 1233 964 1259
rect 862 1229 964 1233
rect 1059 1259 1161 1263
rect 1059 1233 1062 1259
rect 1088 1233 1097 1259
rect 1123 1233 1132 1259
rect 1158 1233 1161 1259
rect 1059 1229 1161 1233
rect 1256 1259 1358 1263
rect 1256 1233 1259 1259
rect 1285 1233 1294 1259
rect 1320 1233 1329 1259
rect 1355 1233 1358 1259
rect 1256 1229 1358 1233
rect 76 694 178 698
rect 76 668 80 694
rect 106 668 114 694
rect 140 668 148 694
rect 174 668 178 694
rect 76 664 178 668
rect 273 695 375 699
rect 471 698 573 699
rect 273 669 277 695
rect 303 669 311 695
rect 337 669 345 695
rect 371 669 375 695
rect 273 664 375 669
rect 469 695 573 698
rect 469 669 475 695
rect 501 669 509 695
rect 535 669 543 695
rect 569 669 573 695
rect 469 664 573 669
rect 667 695 769 699
rect 865 698 967 699
rect 667 669 671 695
rect 697 669 705 695
rect 731 669 739 695
rect 765 669 769 695
rect 667 664 769 669
rect 863 695 967 698
rect 863 669 869 695
rect 895 669 903 695
rect 929 669 937 695
rect 963 669 967 695
rect 863 664 967 669
rect 1061 695 1163 699
rect 1259 698 1361 699
rect 1061 669 1065 695
rect 1091 669 1099 695
rect 1125 669 1133 695
rect 1159 669 1163 695
rect 1061 664 1163 669
rect 1257 695 1361 698
rect 1257 669 1263 695
rect 1289 669 1297 695
rect 1323 669 1331 695
rect 1357 669 1361 695
rect 1257 664 1361 669
rect 74 595 176 599
rect 74 569 78 595
rect 104 569 112 595
rect 138 569 146 595
rect 172 569 176 595
rect 74 564 176 569
rect 273 595 375 599
rect 273 569 277 595
rect 303 569 311 595
rect 337 569 345 595
rect 371 569 375 595
rect 273 564 375 569
rect 468 595 570 599
rect 468 569 472 595
rect 498 569 506 595
rect 532 569 540 595
rect 566 569 570 595
rect 468 564 570 569
rect 667 595 769 599
rect 667 569 671 595
rect 697 569 705 595
rect 731 569 739 595
rect 765 569 769 595
rect 667 564 769 569
rect 862 595 967 599
rect 862 569 869 595
rect 895 569 903 595
rect 929 569 937 595
rect 963 569 967 595
rect 862 565 967 569
rect 865 564 967 565
rect 1061 595 1163 599
rect 1061 569 1065 595
rect 1091 569 1099 595
rect 1125 569 1133 595
rect 1159 569 1163 595
rect 1061 564 1163 569
rect 1257 595 1361 599
rect 1257 569 1263 595
rect 1289 569 1297 595
rect 1323 569 1331 595
rect 1357 569 1361 595
rect 1257 565 1361 569
rect 1259 564 1361 565
rect 74 32 176 36
rect 74 6 77 32
rect 103 6 112 32
rect 138 6 147 32
rect 173 6 176 32
rect 74 2 176 6
rect 271 32 373 36
rect 271 6 274 32
rect 300 6 309 32
rect 335 6 344 32
rect 370 6 373 32
rect 271 2 373 6
rect 468 32 570 36
rect 468 6 471 32
rect 497 6 506 32
rect 532 6 541 32
rect 567 6 570 32
rect 468 2 570 6
rect 665 32 767 36
rect 665 6 668 32
rect 694 6 703 32
rect 729 6 738 32
rect 764 6 767 32
rect 665 2 767 6
rect 862 32 964 36
rect 862 6 865 32
rect 891 6 900 32
rect 926 6 935 32
rect 961 6 964 32
rect 862 2 964 6
rect 1059 32 1161 36
rect 1059 6 1062 32
rect 1088 6 1097 32
rect 1123 6 1132 32
rect 1158 6 1161 32
rect 1059 2 1161 6
rect 1256 32 1358 36
rect 1256 6 1259 32
rect 1285 6 1294 32
rect 1320 6 1329 32
rect 1355 6 1358 32
rect 1256 2 1358 6
rect -193 -109 43 -41
rect 603 -103 829 -41
rect 593 -109 829 -103
rect 1389 -109 1617 -35
rect -193 -135 -175 -109
rect -149 -135 -135 -109
rect -109 -135 -95 -109
rect -69 -135 -55 -109
rect -29 -135 -15 -109
rect 11 -135 25 -109
rect 51 -135 65 -109
rect 91 -135 109 -109
rect -193 -149 109 -135
rect -193 -175 -175 -149
rect -149 -175 -135 -149
rect -109 -175 -95 -149
rect -69 -175 -55 -149
rect -29 -175 -15 -149
rect 11 -175 25 -149
rect 51 -175 65 -149
rect 91 -175 109 -149
rect -193 -189 109 -175
rect -193 -215 -175 -189
rect -149 -215 -135 -189
rect -109 -215 -95 -189
rect -69 -215 -55 -189
rect -29 -215 -15 -189
rect 11 -215 25 -189
rect 51 -215 65 -189
rect 91 -215 109 -189
rect -193 -229 109 -215
rect -193 -255 -175 -229
rect -149 -255 -135 -229
rect -109 -255 -95 -229
rect -69 -255 -55 -229
rect -29 -255 -15 -229
rect 11 -255 25 -229
rect 51 -255 65 -229
rect 91 -255 109 -229
rect -193 -269 109 -255
rect -193 -295 -175 -269
rect -149 -295 -135 -269
rect -109 -295 -95 -269
rect -69 -295 -55 -269
rect -29 -295 -15 -269
rect 11 -295 25 -269
rect 51 -295 65 -269
rect 91 -295 109 -269
rect -193 -309 109 -295
rect -193 -335 -175 -309
rect -149 -335 -135 -309
rect -109 -335 -95 -309
rect -69 -335 -55 -309
rect -29 -335 -15 -309
rect 11 -335 25 -309
rect 51 -335 65 -309
rect 91 -335 109 -309
rect -193 -343 109 -335
rect 565 -135 583 -109
rect 609 -135 623 -109
rect 649 -135 663 -109
rect 689 -135 703 -109
rect 729 -135 743 -109
rect 769 -135 783 -109
rect 809 -135 823 -109
rect 849 -135 867 -109
rect 565 -149 867 -135
rect 565 -175 583 -149
rect 609 -175 623 -149
rect 649 -175 663 -149
rect 689 -175 703 -149
rect 729 -175 743 -149
rect 769 -175 783 -149
rect 809 -175 823 -149
rect 849 -175 867 -149
rect 565 -189 867 -175
rect 565 -215 583 -189
rect 609 -215 623 -189
rect 649 -215 663 -189
rect 689 -215 703 -189
rect 729 -215 743 -189
rect 769 -215 783 -189
rect 809 -215 823 -189
rect 849 -215 867 -189
rect 565 -229 867 -215
rect 565 -255 583 -229
rect 609 -255 623 -229
rect 649 -255 663 -229
rect 689 -255 703 -229
rect 729 -255 743 -229
rect 769 -255 783 -229
rect 809 -255 823 -229
rect 849 -255 867 -229
rect 565 -269 867 -255
rect 565 -295 583 -269
rect 609 -295 623 -269
rect 649 -295 663 -269
rect 689 -295 703 -269
rect 729 -295 743 -269
rect 769 -295 783 -269
rect 809 -295 823 -269
rect 849 -295 867 -269
rect 565 -309 867 -295
rect 565 -335 583 -309
rect 609 -335 623 -309
rect 649 -335 663 -309
rect 689 -335 703 -309
rect 729 -335 743 -309
rect 769 -335 783 -309
rect 809 -335 823 -309
rect 849 -335 867 -309
rect 565 -343 867 -335
rect 1353 -135 1371 -109
rect 1397 -135 1411 -109
rect 1437 -135 1451 -109
rect 1477 -135 1491 -109
rect 1517 -135 1531 -109
rect 1557 -135 1571 -109
rect 1597 -135 1611 -109
rect 1637 -135 1655 -109
rect 1353 -149 1655 -135
rect 1353 -175 1371 -149
rect 1397 -175 1411 -149
rect 1437 -175 1451 -149
rect 1477 -175 1491 -149
rect 1517 -175 1531 -149
rect 1557 -175 1571 -149
rect 1597 -175 1611 -149
rect 1637 -175 1655 -149
rect 1353 -189 1655 -175
rect 1353 -215 1371 -189
rect 1397 -215 1411 -189
rect 1437 -215 1451 -189
rect 1477 -215 1491 -189
rect 1517 -215 1531 -189
rect 1557 -215 1571 -189
rect 1597 -215 1611 -189
rect 1637 -215 1655 -189
rect 1353 -229 1655 -215
rect 1353 -255 1371 -229
rect 1397 -255 1411 -229
rect 1437 -255 1451 -229
rect 1477 -255 1491 -229
rect 1517 -255 1531 -229
rect 1557 -255 1571 -229
rect 1597 -255 1611 -229
rect 1637 -255 1655 -229
rect 1353 -269 1655 -255
rect 1353 -295 1371 -269
rect 1397 -295 1411 -269
rect 1437 -295 1451 -269
rect 1477 -295 1491 -269
rect 1517 -295 1531 -269
rect 1557 -295 1571 -269
rect 1597 -295 1611 -269
rect 1637 -295 1655 -269
rect 1353 -309 1655 -295
rect 1353 -335 1371 -309
rect 1397 -335 1411 -309
rect 1437 -335 1451 -309
rect 1477 -335 1491 -309
rect 1517 -335 1531 -309
rect 1557 -335 1571 -309
rect 1597 -335 1611 -309
rect 1637 -335 1655 -309
rect 1353 -343 1655 -335
<< via1 >>
rect 77 1233 103 1259
rect 112 1233 138 1259
rect 147 1233 173 1259
rect 274 1233 300 1259
rect 309 1233 335 1259
rect 344 1233 370 1259
rect 471 1233 497 1259
rect 506 1233 532 1259
rect 541 1233 567 1259
rect 668 1233 694 1259
rect 703 1233 729 1259
rect 738 1233 764 1259
rect 865 1233 891 1259
rect 900 1233 926 1259
rect 935 1233 961 1259
rect 1062 1233 1088 1259
rect 1097 1233 1123 1259
rect 1132 1233 1158 1259
rect 1259 1233 1285 1259
rect 1294 1233 1320 1259
rect 1329 1233 1355 1259
rect 80 668 106 694
rect 114 668 140 694
rect 148 668 174 694
rect 277 669 303 695
rect 311 669 337 695
rect 345 669 371 695
rect 475 669 501 695
rect 509 669 535 695
rect 543 669 569 695
rect 671 669 697 695
rect 705 669 731 695
rect 739 669 765 695
rect 869 669 895 695
rect 903 669 929 695
rect 937 669 963 695
rect 1065 669 1091 695
rect 1099 669 1125 695
rect 1133 669 1159 695
rect 1263 669 1289 695
rect 1297 669 1323 695
rect 1331 669 1357 695
rect 78 569 104 595
rect 112 569 138 595
rect 146 569 172 595
rect 277 569 303 595
rect 311 569 337 595
rect 345 569 371 595
rect 472 569 498 595
rect 506 569 532 595
rect 540 569 566 595
rect 671 569 697 595
rect 705 569 731 595
rect 739 569 765 595
rect 869 569 895 595
rect 903 569 929 595
rect 937 569 963 595
rect 1065 569 1091 595
rect 1099 569 1125 595
rect 1133 569 1159 595
rect 1263 569 1289 595
rect 1297 569 1323 595
rect 1331 569 1357 595
rect 77 6 103 32
rect 112 6 138 32
rect 147 6 173 32
rect 274 6 300 32
rect 309 6 335 32
rect 344 6 370 32
rect 471 6 497 32
rect 506 6 532 32
rect 541 6 567 32
rect 668 6 694 32
rect 703 6 729 32
rect 738 6 764 32
rect 865 6 891 32
rect 900 6 926 32
rect 935 6 961 32
rect 1062 6 1088 32
rect 1097 6 1123 32
rect 1132 6 1158 32
rect 1259 6 1285 32
rect 1294 6 1320 32
rect 1329 6 1355 32
rect -175 -135 -149 -109
rect -135 -135 -109 -109
rect -95 -135 -69 -109
rect -55 -135 -29 -109
rect -15 -135 11 -109
rect 25 -135 51 -109
rect 65 -135 91 -109
rect -175 -175 -149 -149
rect -135 -175 -109 -149
rect -95 -175 -69 -149
rect -55 -175 -29 -149
rect -15 -175 11 -149
rect 25 -175 51 -149
rect 65 -175 91 -149
rect -175 -215 -149 -189
rect -135 -215 -109 -189
rect -95 -215 -69 -189
rect -55 -215 -29 -189
rect -15 -215 11 -189
rect 25 -215 51 -189
rect 65 -215 91 -189
rect -175 -255 -149 -229
rect -135 -255 -109 -229
rect -95 -255 -69 -229
rect -55 -255 -29 -229
rect -15 -255 11 -229
rect 25 -255 51 -229
rect 65 -255 91 -229
rect -175 -295 -149 -269
rect -135 -295 -109 -269
rect -95 -295 -69 -269
rect -55 -295 -29 -269
rect -15 -295 11 -269
rect 25 -295 51 -269
rect 65 -295 91 -269
rect -175 -335 -149 -309
rect -135 -335 -109 -309
rect -95 -335 -69 -309
rect -55 -335 -29 -309
rect -15 -335 11 -309
rect 25 -335 51 -309
rect 65 -335 91 -309
rect 583 -135 609 -109
rect 623 -135 649 -109
rect 663 -135 689 -109
rect 703 -135 729 -109
rect 743 -135 769 -109
rect 783 -135 809 -109
rect 823 -135 849 -109
rect 583 -175 609 -149
rect 623 -175 649 -149
rect 663 -175 689 -149
rect 703 -175 729 -149
rect 743 -175 769 -149
rect 783 -175 809 -149
rect 823 -175 849 -149
rect 583 -215 609 -189
rect 623 -215 649 -189
rect 663 -215 689 -189
rect 703 -215 729 -189
rect 743 -215 769 -189
rect 783 -215 809 -189
rect 823 -215 849 -189
rect 583 -255 609 -229
rect 623 -255 649 -229
rect 663 -255 689 -229
rect 703 -255 729 -229
rect 743 -255 769 -229
rect 783 -255 809 -229
rect 823 -255 849 -229
rect 583 -295 609 -269
rect 623 -295 649 -269
rect 663 -295 689 -269
rect 703 -295 729 -269
rect 743 -295 769 -269
rect 783 -295 809 -269
rect 823 -295 849 -269
rect 583 -335 609 -309
rect 623 -335 649 -309
rect 663 -335 689 -309
rect 703 -335 729 -309
rect 743 -335 769 -309
rect 783 -335 809 -309
rect 823 -335 849 -309
rect 1371 -135 1397 -109
rect 1411 -135 1437 -109
rect 1451 -135 1477 -109
rect 1491 -135 1517 -109
rect 1531 -135 1557 -109
rect 1571 -135 1597 -109
rect 1611 -135 1637 -109
rect 1371 -175 1397 -149
rect 1411 -175 1437 -149
rect 1451 -175 1477 -149
rect 1491 -175 1517 -149
rect 1531 -175 1557 -149
rect 1571 -175 1597 -149
rect 1611 -175 1637 -149
rect 1371 -215 1397 -189
rect 1411 -215 1437 -189
rect 1451 -215 1477 -189
rect 1491 -215 1517 -189
rect 1531 -215 1557 -189
rect 1571 -215 1597 -189
rect 1611 -215 1637 -189
rect 1371 -255 1397 -229
rect 1411 -255 1437 -229
rect 1451 -255 1477 -229
rect 1491 -255 1517 -229
rect 1531 -255 1557 -229
rect 1571 -255 1597 -229
rect 1611 -255 1637 -229
rect 1371 -295 1397 -269
rect 1411 -295 1437 -269
rect 1451 -295 1477 -269
rect 1491 -295 1517 -269
rect 1531 -295 1557 -269
rect 1571 -295 1597 -269
rect 1611 -295 1637 -269
rect 1371 -335 1397 -309
rect 1411 -335 1437 -309
rect 1451 -335 1477 -309
rect 1491 -335 1517 -309
rect 1531 -335 1557 -309
rect 1571 -335 1597 -309
rect 1611 -335 1637 -309
<< metal2 >>
rect 271 1324 373 1327
rect 271 1296 276 1324
rect 304 1296 340 1324
rect 368 1296 373 1324
rect 74 1260 176 1263
rect 74 1259 79 1260
rect 107 1259 143 1260
rect 171 1259 176 1260
rect 74 1233 77 1259
rect 107 1233 112 1259
rect 138 1233 143 1259
rect 173 1233 176 1259
rect 74 1232 79 1233
rect 107 1232 143 1233
rect 171 1232 176 1233
rect 74 1229 176 1232
rect 271 1259 373 1296
rect 665 1324 767 1327
rect 665 1296 670 1324
rect 698 1296 734 1324
rect 762 1296 767 1324
rect 271 1233 274 1259
rect 300 1233 309 1259
rect 335 1233 344 1259
rect 370 1233 373 1259
rect 271 1229 373 1233
rect 468 1260 570 1263
rect 468 1259 473 1260
rect 501 1259 537 1260
rect 565 1259 570 1260
rect 468 1233 471 1259
rect 501 1233 506 1259
rect 532 1233 537 1259
rect 567 1233 570 1259
rect 468 1232 473 1233
rect 501 1232 537 1233
rect 565 1232 570 1233
rect 468 1229 570 1232
rect 665 1259 767 1296
rect 1059 1324 1161 1327
rect 1059 1296 1064 1324
rect 1092 1296 1128 1324
rect 1156 1296 1161 1324
rect 665 1233 668 1259
rect 694 1233 703 1259
rect 729 1233 738 1259
rect 764 1233 767 1259
rect 665 1229 767 1233
rect 862 1260 964 1263
rect 862 1259 867 1260
rect 895 1259 931 1260
rect 959 1259 964 1260
rect 862 1233 865 1259
rect 895 1233 900 1259
rect 926 1233 931 1259
rect 961 1233 964 1259
rect 862 1232 867 1233
rect 895 1232 931 1233
rect 959 1232 964 1233
rect 862 1229 964 1232
rect 1059 1259 1161 1296
rect 1059 1233 1062 1259
rect 1088 1233 1097 1259
rect 1123 1233 1132 1259
rect 1158 1233 1161 1259
rect 1059 1229 1161 1233
rect 1256 1260 1358 1263
rect 1256 1259 1261 1260
rect 1289 1259 1325 1260
rect 1353 1259 1358 1260
rect 1256 1233 1259 1259
rect 1289 1233 1294 1259
rect 1320 1233 1325 1259
rect 1355 1233 1358 1259
rect 1256 1232 1261 1233
rect 1289 1232 1325 1233
rect 1353 1232 1358 1233
rect 1256 1229 1358 1232
rect 70 939 184 950
rect 70 911 73 939
rect 101 911 113 939
rect 141 911 153 939
rect 181 911 184 939
rect 70 899 184 911
rect 70 871 73 899
rect 101 871 113 899
rect 141 871 153 899
rect 181 871 184 899
rect 70 860 184 871
rect 464 939 578 950
rect 464 911 467 939
rect 495 911 507 939
rect 535 911 547 939
rect 575 911 578 939
rect 464 899 578 911
rect 464 871 467 899
rect 495 871 507 899
rect 535 871 547 899
rect 575 871 578 899
rect 464 860 578 871
rect 858 939 972 950
rect 858 911 861 939
rect 889 911 901 939
rect 929 911 941 939
rect 969 911 972 939
rect 858 899 972 911
rect 858 871 861 899
rect 889 871 901 899
rect 929 871 941 899
rect 969 871 972 899
rect 858 860 972 871
rect 1252 939 1366 950
rect 1252 911 1255 939
rect 1283 911 1295 939
rect 1323 911 1335 939
rect 1363 911 1366 939
rect 1252 899 1366 911
rect 1252 871 1255 899
rect 1283 871 1295 899
rect 1323 871 1335 899
rect 1363 871 1366 899
rect 1252 860 1366 871
rect 267 807 381 818
rect 267 779 270 807
rect 298 779 310 807
rect 338 779 350 807
rect 378 779 381 807
rect 267 767 381 779
rect 267 739 270 767
rect 298 739 310 767
rect 338 739 350 767
rect 378 739 381 767
rect 267 728 381 739
rect 661 807 775 818
rect 661 779 664 807
rect 692 779 704 807
rect 732 779 744 807
rect 772 779 775 807
rect 661 767 775 779
rect 661 739 664 767
rect 692 739 704 767
rect 732 739 744 767
rect 772 739 775 767
rect 661 728 775 739
rect 1055 807 1169 818
rect 1055 779 1058 807
rect 1086 779 1098 807
rect 1126 779 1138 807
rect 1166 779 1169 807
rect 1055 767 1169 779
rect 1055 739 1058 767
rect 1086 739 1098 767
rect 1126 739 1138 767
rect 1166 739 1169 767
rect 1055 728 1169 739
rect 273 698 375 699
rect 471 698 573 699
rect 667 698 769 699
rect 865 698 967 699
rect 1061 698 1163 699
rect 1259 698 1361 699
rect 76 695 178 698
rect 76 694 93 695
rect 121 694 133 695
rect 161 694 178 695
rect 76 668 80 694
rect 174 668 178 694
rect 76 667 93 668
rect 121 667 133 668
rect 161 667 178 668
rect 76 664 178 667
rect 210 695 375 698
rect 210 669 277 695
rect 371 669 375 695
rect 210 667 289 669
rect 317 667 329 669
rect 357 667 375 669
rect 210 664 375 667
rect 407 695 573 698
rect 407 669 475 695
rect 569 669 573 695
rect 407 667 487 669
rect 515 667 527 669
rect 555 667 573 669
rect 407 664 573 667
rect 604 695 769 698
rect 604 669 671 695
rect 765 669 769 695
rect 604 667 683 669
rect 711 667 723 669
rect 751 667 769 669
rect 604 664 769 667
rect 801 695 967 698
rect 801 669 869 695
rect 963 669 967 695
rect 801 667 881 669
rect 909 667 921 669
rect 949 667 967 669
rect 801 664 967 667
rect 998 695 1163 698
rect 998 669 1065 695
rect 1159 669 1163 695
rect 998 667 1077 669
rect 1105 667 1117 669
rect 1145 667 1163 669
rect 998 664 1163 667
rect 1195 695 1361 698
rect 1195 669 1263 695
rect 1357 669 1361 695
rect 1195 667 1275 669
rect 1303 667 1315 669
rect 1343 667 1361 669
rect 1195 664 1361 667
rect 210 599 241 664
rect 407 599 438 664
rect 604 599 635 664
rect 801 599 832 664
rect 998 599 1029 664
rect 1195 599 1226 664
rect 74 596 241 599
rect 74 595 93 596
rect 121 595 133 596
rect 161 595 241 596
rect 74 569 78 595
rect 172 569 241 595
rect 74 568 93 569
rect 121 568 133 569
rect 161 568 241 569
rect 74 565 241 568
rect 273 596 438 599
rect 273 595 289 596
rect 317 595 329 596
rect 357 595 438 596
rect 273 569 277 595
rect 371 569 438 595
rect 273 568 289 569
rect 317 568 329 569
rect 357 568 438 569
rect 273 565 438 568
rect 468 596 635 599
rect 468 595 487 596
rect 515 595 527 596
rect 555 595 635 596
rect 468 569 472 595
rect 566 569 635 595
rect 468 568 487 569
rect 515 568 527 569
rect 555 568 635 569
rect 468 565 635 568
rect 667 596 832 599
rect 667 595 683 596
rect 711 595 723 596
rect 751 595 832 596
rect 667 569 671 595
rect 765 569 832 595
rect 667 568 683 569
rect 711 568 723 569
rect 751 568 832 569
rect 667 565 832 568
rect 862 596 1029 599
rect 862 595 881 596
rect 909 595 921 596
rect 949 595 1029 596
rect 862 569 869 595
rect 963 569 1029 595
rect 862 568 881 569
rect 909 568 921 569
rect 949 568 1029 569
rect 862 565 1029 568
rect 1061 596 1226 599
rect 1061 595 1077 596
rect 1105 595 1117 596
rect 1145 595 1226 596
rect 1061 569 1065 595
rect 1159 569 1226 595
rect 1061 568 1077 569
rect 1105 568 1117 569
rect 1145 568 1226 569
rect 1061 565 1226 568
rect 1256 596 1361 599
rect 1256 595 1275 596
rect 1303 595 1315 596
rect 1343 595 1361 596
rect 1256 569 1263 595
rect 1357 569 1361 595
rect 1256 568 1275 569
rect 1303 568 1315 569
rect 1343 568 1361 569
rect 1256 565 1361 568
rect 74 564 176 565
rect 273 564 375 565
rect 468 564 570 565
rect 667 564 769 565
rect 865 564 967 565
rect 1061 564 1163 565
rect 1259 564 1361 565
rect 267 523 381 534
rect 267 495 270 523
rect 298 495 310 523
rect 338 495 350 523
rect 378 495 381 523
rect 267 483 381 495
rect 267 455 270 483
rect 298 455 310 483
rect 338 455 350 483
rect 378 455 381 483
rect 267 444 381 455
rect 661 523 775 534
rect 661 495 664 523
rect 692 495 704 523
rect 732 495 744 523
rect 772 495 775 523
rect 661 483 775 495
rect 661 455 664 483
rect 692 455 704 483
rect 732 455 744 483
rect 772 455 775 483
rect 661 444 775 455
rect 1055 523 1169 534
rect 1055 495 1058 523
rect 1086 495 1098 523
rect 1126 495 1138 523
rect 1166 495 1169 523
rect 1055 483 1169 495
rect 1055 455 1058 483
rect 1086 455 1098 483
rect 1126 455 1138 483
rect 1166 455 1169 483
rect 1055 444 1169 455
rect 70 390 184 401
rect 70 362 73 390
rect 101 362 113 390
rect 141 362 153 390
rect 181 362 184 390
rect 70 350 184 362
rect 70 322 73 350
rect 101 322 113 350
rect 141 322 153 350
rect 181 322 184 350
rect 70 311 184 322
rect 464 390 578 401
rect 464 362 467 390
rect 495 362 507 390
rect 535 362 547 390
rect 575 362 578 390
rect 464 350 578 362
rect 464 322 467 350
rect 495 322 507 350
rect 535 322 547 350
rect 575 322 578 350
rect 464 311 578 322
rect 858 390 972 401
rect 858 362 861 390
rect 889 362 901 390
rect 929 362 941 390
rect 969 362 972 390
rect 858 350 972 362
rect 858 322 861 350
rect 889 322 901 350
rect 929 322 941 350
rect 969 322 972 350
rect 858 311 972 322
rect 1252 390 1366 401
rect 1252 362 1255 390
rect 1283 362 1295 390
rect 1323 362 1335 390
rect 1363 362 1366 390
rect 1252 350 1366 362
rect 1252 322 1255 350
rect 1283 322 1295 350
rect 1323 322 1335 350
rect 1363 322 1366 350
rect 1252 311 1366 322
rect 74 33 176 36
rect 74 32 79 33
rect 107 32 143 33
rect 171 32 176 33
rect 74 6 77 32
rect 107 6 112 32
rect 138 6 143 32
rect 173 6 176 32
rect 74 5 79 6
rect 107 5 143 6
rect 171 5 176 6
rect 74 2 176 5
rect 271 32 373 36
rect 271 6 274 32
rect 300 6 309 32
rect 335 6 344 32
rect 370 6 373 32
rect 271 -31 373 6
rect 468 33 570 36
rect 468 32 473 33
rect 501 32 537 33
rect 565 32 570 33
rect 468 6 471 32
rect 501 6 506 32
rect 532 6 537 32
rect 567 6 570 32
rect 468 5 473 6
rect 501 5 537 6
rect 565 5 570 6
rect 468 2 570 5
rect 665 32 767 36
rect 665 6 668 32
rect 694 6 703 32
rect 729 6 738 32
rect 764 6 767 32
rect 271 -59 276 -31
rect 304 -59 340 -31
rect 368 -59 373 -31
rect 271 -62 373 -59
rect 665 -31 767 6
rect 862 33 964 36
rect 862 32 867 33
rect 895 32 931 33
rect 959 32 964 33
rect 862 6 865 32
rect 895 6 900 32
rect 926 6 931 32
rect 961 6 964 32
rect 862 5 867 6
rect 895 5 931 6
rect 959 5 964 6
rect 862 2 964 5
rect 1059 32 1161 36
rect 1059 6 1062 32
rect 1088 6 1097 32
rect 1123 6 1132 32
rect 1158 6 1161 32
rect 665 -59 670 -31
rect 698 -59 734 -31
rect 762 -59 767 -31
rect 665 -62 767 -59
rect 1059 -31 1161 6
rect 1256 33 1358 36
rect 1256 32 1261 33
rect 1289 32 1325 33
rect 1353 32 1358 33
rect 1256 6 1259 32
rect 1289 6 1294 32
rect 1320 6 1325 32
rect 1355 6 1358 32
rect 1256 5 1261 6
rect 1289 5 1325 6
rect 1353 5 1358 6
rect 1256 2 1358 5
rect 1059 -59 1064 -31
rect 1092 -59 1128 -31
rect 1156 -59 1161 -31
rect 1059 -62 1161 -59
rect -193 -108 109 -107
rect -193 -136 -176 -108
rect -148 -136 -136 -108
rect -108 -136 -96 -108
rect -68 -136 -56 -108
rect -28 -136 -16 -108
rect 12 -136 24 -108
rect 52 -136 64 -108
rect 92 -136 109 -108
rect -193 -148 109 -136
rect -193 -176 -176 -148
rect -148 -176 -136 -148
rect -108 -176 -96 -148
rect -68 -176 -56 -148
rect -28 -176 -16 -148
rect 12 -176 24 -148
rect 52 -176 64 -148
rect 92 -176 109 -148
rect -193 -188 109 -176
rect -193 -216 -176 -188
rect -148 -216 -136 -188
rect -108 -216 -96 -188
rect -68 -216 -56 -188
rect -28 -216 -16 -188
rect 12 -216 24 -188
rect 52 -216 64 -188
rect 92 -216 109 -188
rect -193 -228 109 -216
rect -193 -256 -176 -228
rect -148 -256 -136 -228
rect -108 -256 -96 -228
rect -68 -256 -56 -228
rect -28 -256 -16 -228
rect 12 -256 24 -228
rect 52 -256 64 -228
rect 92 -256 109 -228
rect -193 -268 109 -256
rect -193 -296 -176 -268
rect -148 -296 -136 -268
rect -108 -296 -96 -268
rect -68 -296 -56 -268
rect -28 -296 -16 -268
rect 12 -296 24 -268
rect 52 -296 64 -268
rect 92 -296 109 -268
rect -193 -308 109 -296
rect -193 -336 -176 -308
rect -148 -336 -136 -308
rect -108 -336 -96 -308
rect -68 -336 -56 -308
rect -28 -336 -16 -308
rect 12 -336 24 -308
rect 52 -336 64 -308
rect 92 -336 109 -308
rect -193 -343 109 -336
rect 565 -108 867 -107
rect 565 -136 582 -108
rect 610 -136 622 -108
rect 650 -136 662 -108
rect 690 -136 702 -108
rect 730 -136 742 -108
rect 770 -136 782 -108
rect 810 -136 822 -108
rect 850 -136 867 -108
rect 565 -148 867 -136
rect 565 -176 582 -148
rect 610 -176 622 -148
rect 650 -176 662 -148
rect 690 -176 702 -148
rect 730 -176 742 -148
rect 770 -176 782 -148
rect 810 -176 822 -148
rect 850 -176 867 -148
rect 565 -188 867 -176
rect 565 -216 582 -188
rect 610 -216 622 -188
rect 650 -216 662 -188
rect 690 -216 702 -188
rect 730 -216 742 -188
rect 770 -216 782 -188
rect 810 -216 822 -188
rect 850 -216 867 -188
rect 565 -228 867 -216
rect 565 -256 582 -228
rect 610 -256 622 -228
rect 650 -256 662 -228
rect 690 -256 702 -228
rect 730 -256 742 -228
rect 770 -256 782 -228
rect 810 -256 822 -228
rect 850 -256 867 -228
rect 565 -268 867 -256
rect 565 -296 582 -268
rect 610 -296 622 -268
rect 650 -296 662 -268
rect 690 -296 702 -268
rect 730 -296 742 -268
rect 770 -296 782 -268
rect 810 -296 822 -268
rect 850 -296 867 -268
rect 565 -308 867 -296
rect 565 -336 582 -308
rect 610 -336 622 -308
rect 650 -336 662 -308
rect 690 -336 702 -308
rect 730 -336 742 -308
rect 770 -336 782 -308
rect 810 -336 822 -308
rect 850 -336 867 -308
rect 565 -343 867 -336
rect 1353 -108 1655 -107
rect 1353 -136 1370 -108
rect 1398 -136 1410 -108
rect 1438 -136 1450 -108
rect 1478 -136 1490 -108
rect 1518 -136 1530 -108
rect 1558 -136 1570 -108
rect 1598 -136 1610 -108
rect 1638 -136 1655 -108
rect 1353 -148 1655 -136
rect 1353 -176 1370 -148
rect 1398 -176 1410 -148
rect 1438 -176 1450 -148
rect 1478 -176 1490 -148
rect 1518 -176 1530 -148
rect 1558 -176 1570 -148
rect 1598 -176 1610 -148
rect 1638 -176 1655 -148
rect 1353 -188 1655 -176
rect 1353 -216 1370 -188
rect 1398 -216 1410 -188
rect 1438 -216 1450 -188
rect 1478 -216 1490 -188
rect 1518 -216 1530 -188
rect 1558 -216 1570 -188
rect 1598 -216 1610 -188
rect 1638 -216 1655 -188
rect 1353 -228 1655 -216
rect 1353 -256 1370 -228
rect 1398 -256 1410 -228
rect 1438 -256 1450 -228
rect 1478 -256 1490 -228
rect 1518 -256 1530 -228
rect 1558 -256 1570 -228
rect 1598 -256 1610 -228
rect 1638 -256 1655 -228
rect 1353 -268 1655 -256
rect 1353 -296 1370 -268
rect 1398 -296 1410 -268
rect 1438 -296 1450 -268
rect 1478 -296 1490 -268
rect 1518 -296 1530 -268
rect 1558 -296 1570 -268
rect 1598 -296 1610 -268
rect 1638 -296 1655 -268
rect 1353 -308 1655 -296
rect 1353 -336 1370 -308
rect 1398 -336 1410 -308
rect 1438 -336 1450 -308
rect 1478 -336 1490 -308
rect 1518 -336 1530 -308
rect 1558 -336 1570 -308
rect 1598 -336 1610 -308
rect 1638 -336 1655 -308
rect 1353 -343 1655 -336
<< via2 >>
rect 276 1296 304 1324
rect 340 1296 368 1324
rect 79 1259 107 1260
rect 143 1259 171 1260
rect 79 1233 103 1259
rect 103 1233 107 1259
rect 143 1233 147 1259
rect 147 1233 171 1259
rect 79 1232 107 1233
rect 143 1232 171 1233
rect 670 1296 698 1324
rect 734 1296 762 1324
rect 473 1259 501 1260
rect 537 1259 565 1260
rect 473 1233 497 1259
rect 497 1233 501 1259
rect 537 1233 541 1259
rect 541 1233 565 1259
rect 473 1232 501 1233
rect 537 1232 565 1233
rect 1064 1296 1092 1324
rect 1128 1296 1156 1324
rect 867 1259 895 1260
rect 931 1259 959 1260
rect 867 1233 891 1259
rect 891 1233 895 1259
rect 931 1233 935 1259
rect 935 1233 959 1259
rect 867 1232 895 1233
rect 931 1232 959 1233
rect 1261 1259 1289 1260
rect 1325 1259 1353 1260
rect 1261 1233 1285 1259
rect 1285 1233 1289 1259
rect 1325 1233 1329 1259
rect 1329 1233 1353 1259
rect 1261 1232 1289 1233
rect 1325 1232 1353 1233
rect 73 1155 101 1183
rect 113 1155 141 1183
rect 153 1155 181 1183
rect 270 1155 298 1183
rect 310 1155 338 1183
rect 350 1155 378 1183
rect 467 1155 495 1183
rect 507 1155 535 1183
rect 547 1155 575 1183
rect 664 1155 692 1183
rect 704 1155 732 1183
rect 744 1155 772 1183
rect 861 1155 889 1183
rect 901 1155 929 1183
rect 941 1155 969 1183
rect 1058 1155 1086 1183
rect 1098 1155 1126 1183
rect 1138 1155 1166 1183
rect 1255 1155 1283 1183
rect 1295 1155 1323 1183
rect 1335 1155 1363 1183
rect 73 1115 101 1143
rect 113 1115 141 1143
rect 153 1115 181 1143
rect 270 1115 298 1143
rect 310 1115 338 1143
rect 350 1115 378 1143
rect 467 1115 495 1143
rect 507 1115 535 1143
rect 547 1115 575 1143
rect 664 1115 692 1143
rect 704 1115 732 1143
rect 744 1115 772 1143
rect 861 1115 889 1143
rect 901 1115 929 1143
rect 941 1115 969 1143
rect 1058 1115 1086 1143
rect 1098 1115 1126 1143
rect 1138 1115 1166 1143
rect 1255 1115 1283 1143
rect 1295 1115 1323 1143
rect 1335 1115 1363 1143
rect 73 1075 101 1103
rect 113 1075 141 1103
rect 153 1075 181 1103
rect 270 1075 298 1103
rect 310 1075 338 1103
rect 350 1075 378 1103
rect 467 1075 495 1103
rect 507 1075 535 1103
rect 547 1075 575 1103
rect 664 1075 692 1103
rect 704 1075 732 1103
rect 744 1075 772 1103
rect 861 1075 889 1103
rect 901 1075 929 1103
rect 941 1075 969 1103
rect 1058 1075 1086 1103
rect 1098 1075 1126 1103
rect 1138 1075 1166 1103
rect 1255 1075 1283 1103
rect 1295 1075 1323 1103
rect 1335 1075 1363 1103
rect 73 1035 101 1063
rect 113 1035 141 1063
rect 153 1035 181 1063
rect 270 1035 298 1063
rect 310 1035 338 1063
rect 350 1035 378 1063
rect 467 1035 495 1063
rect 507 1035 535 1063
rect 547 1035 575 1063
rect 664 1035 692 1063
rect 704 1035 732 1063
rect 744 1035 772 1063
rect 861 1035 889 1063
rect 901 1035 929 1063
rect 941 1035 969 1063
rect 1058 1035 1086 1063
rect 1098 1035 1126 1063
rect 1138 1035 1166 1063
rect 1255 1035 1283 1063
rect 1295 1035 1323 1063
rect 1335 1035 1363 1063
rect 73 995 101 1023
rect 113 995 141 1023
rect 153 995 181 1023
rect 270 995 298 1023
rect 310 995 338 1023
rect 350 995 378 1023
rect 467 995 495 1023
rect 507 995 535 1023
rect 547 995 575 1023
rect 664 995 692 1023
rect 704 995 732 1023
rect 744 995 772 1023
rect 861 995 889 1023
rect 901 995 929 1023
rect 941 995 969 1023
rect 1058 995 1086 1023
rect 1098 995 1126 1023
rect 1138 995 1166 1023
rect 1255 995 1283 1023
rect 1295 995 1323 1023
rect 1335 995 1363 1023
rect 73 911 101 939
rect 113 911 141 939
rect 153 911 181 939
rect 73 871 101 899
rect 113 871 141 899
rect 153 871 181 899
rect 467 911 495 939
rect 507 911 535 939
rect 547 911 575 939
rect 467 871 495 899
rect 507 871 535 899
rect 547 871 575 899
rect 861 911 889 939
rect 901 911 929 939
rect 941 911 969 939
rect 861 871 889 899
rect 901 871 929 899
rect 941 871 969 899
rect 1255 911 1283 939
rect 1295 911 1323 939
rect 1335 911 1363 939
rect 1255 871 1283 899
rect 1295 871 1323 899
rect 1335 871 1363 899
rect 270 779 298 807
rect 310 779 338 807
rect 350 779 378 807
rect 270 739 298 767
rect 310 739 338 767
rect 350 739 378 767
rect 664 779 692 807
rect 704 779 732 807
rect 744 779 772 807
rect 664 739 692 767
rect 704 739 732 767
rect 744 739 772 767
rect 1058 779 1086 807
rect 1098 779 1126 807
rect 1138 779 1166 807
rect 1058 739 1086 767
rect 1098 739 1126 767
rect 1138 739 1166 767
rect 93 694 121 695
rect 133 694 161 695
rect 93 668 106 694
rect 106 668 114 694
rect 114 668 121 694
rect 133 668 140 694
rect 140 668 148 694
rect 148 668 161 694
rect 93 667 121 668
rect 133 667 161 668
rect 289 669 303 695
rect 303 669 311 695
rect 311 669 317 695
rect 329 669 337 695
rect 337 669 345 695
rect 345 669 357 695
rect 289 667 317 669
rect 329 667 357 669
rect 487 669 501 695
rect 501 669 509 695
rect 509 669 515 695
rect 527 669 535 695
rect 535 669 543 695
rect 543 669 555 695
rect 487 667 515 669
rect 527 667 555 669
rect 683 669 697 695
rect 697 669 705 695
rect 705 669 711 695
rect 723 669 731 695
rect 731 669 739 695
rect 739 669 751 695
rect 683 667 711 669
rect 723 667 751 669
rect 881 669 895 695
rect 895 669 903 695
rect 903 669 909 695
rect 921 669 929 695
rect 929 669 937 695
rect 937 669 949 695
rect 881 667 909 669
rect 921 667 949 669
rect 1077 669 1091 695
rect 1091 669 1099 695
rect 1099 669 1105 695
rect 1117 669 1125 695
rect 1125 669 1133 695
rect 1133 669 1145 695
rect 1077 667 1105 669
rect 1117 667 1145 669
rect 1275 669 1289 695
rect 1289 669 1297 695
rect 1297 669 1303 695
rect 1315 669 1323 695
rect 1323 669 1331 695
rect 1331 669 1343 695
rect 1275 667 1303 669
rect 1315 667 1343 669
rect 93 595 121 596
rect 133 595 161 596
rect 93 569 104 595
rect 104 569 112 595
rect 112 569 121 595
rect 133 569 138 595
rect 138 569 146 595
rect 146 569 161 595
rect 93 568 121 569
rect 133 568 161 569
rect 289 595 317 596
rect 329 595 357 596
rect 289 569 303 595
rect 303 569 311 595
rect 311 569 317 595
rect 329 569 337 595
rect 337 569 345 595
rect 345 569 357 595
rect 289 568 317 569
rect 329 568 357 569
rect 487 595 515 596
rect 527 595 555 596
rect 487 569 498 595
rect 498 569 506 595
rect 506 569 515 595
rect 527 569 532 595
rect 532 569 540 595
rect 540 569 555 595
rect 487 568 515 569
rect 527 568 555 569
rect 683 595 711 596
rect 723 595 751 596
rect 683 569 697 595
rect 697 569 705 595
rect 705 569 711 595
rect 723 569 731 595
rect 731 569 739 595
rect 739 569 751 595
rect 683 568 711 569
rect 723 568 751 569
rect 881 595 909 596
rect 921 595 949 596
rect 881 569 895 595
rect 895 569 903 595
rect 903 569 909 595
rect 921 569 929 595
rect 929 569 937 595
rect 937 569 949 595
rect 881 568 909 569
rect 921 568 949 569
rect 1077 595 1105 596
rect 1117 595 1145 596
rect 1077 569 1091 595
rect 1091 569 1099 595
rect 1099 569 1105 595
rect 1117 569 1125 595
rect 1125 569 1133 595
rect 1133 569 1145 595
rect 1077 568 1105 569
rect 1117 568 1145 569
rect 1275 595 1303 596
rect 1315 595 1343 596
rect 1275 569 1289 595
rect 1289 569 1297 595
rect 1297 569 1303 595
rect 1315 569 1323 595
rect 1323 569 1331 595
rect 1331 569 1343 595
rect 1275 568 1303 569
rect 1315 568 1343 569
rect 270 495 298 523
rect 310 495 338 523
rect 350 495 378 523
rect 270 455 298 483
rect 310 455 338 483
rect 350 455 378 483
rect 664 495 692 523
rect 704 495 732 523
rect 744 495 772 523
rect 664 455 692 483
rect 704 455 732 483
rect 744 455 772 483
rect 1058 495 1086 523
rect 1098 495 1126 523
rect 1138 495 1166 523
rect 1058 455 1086 483
rect 1098 455 1126 483
rect 1138 455 1166 483
rect 73 362 101 390
rect 113 362 141 390
rect 153 362 181 390
rect 73 322 101 350
rect 113 322 141 350
rect 153 322 181 350
rect 467 362 495 390
rect 507 362 535 390
rect 547 362 575 390
rect 467 322 495 350
rect 507 322 535 350
rect 547 322 575 350
rect 861 362 889 390
rect 901 362 929 390
rect 941 362 969 390
rect 861 322 889 350
rect 901 322 929 350
rect 941 322 969 350
rect 1255 362 1283 390
rect 1295 362 1323 390
rect 1335 362 1363 390
rect 1255 322 1283 350
rect 1295 322 1323 350
rect 1335 322 1363 350
rect 73 233 101 261
rect 113 233 141 261
rect 153 233 181 261
rect 270 233 298 261
rect 310 233 338 261
rect 350 233 378 261
rect 467 233 495 261
rect 507 233 535 261
rect 547 233 575 261
rect 664 233 692 261
rect 704 233 732 261
rect 744 233 772 261
rect 861 233 889 261
rect 901 233 929 261
rect 941 233 969 261
rect 1058 233 1086 261
rect 1098 233 1126 261
rect 1138 233 1166 261
rect 1255 233 1283 261
rect 1295 233 1323 261
rect 1335 233 1363 261
rect 73 193 101 221
rect 113 193 141 221
rect 153 193 181 221
rect 270 193 298 221
rect 310 193 338 221
rect 350 193 378 221
rect 467 193 495 221
rect 507 193 535 221
rect 547 193 575 221
rect 664 193 692 221
rect 704 193 732 221
rect 744 193 772 221
rect 861 193 889 221
rect 901 193 929 221
rect 941 193 969 221
rect 1058 193 1086 221
rect 1098 193 1126 221
rect 1138 193 1166 221
rect 1255 193 1283 221
rect 1295 193 1323 221
rect 1335 193 1363 221
rect 73 153 101 181
rect 113 153 141 181
rect 153 153 181 181
rect 270 153 298 181
rect 310 153 338 181
rect 350 153 378 181
rect 467 153 495 181
rect 507 153 535 181
rect 547 153 575 181
rect 664 153 692 181
rect 704 153 732 181
rect 744 153 772 181
rect 861 153 889 181
rect 901 153 929 181
rect 941 153 969 181
rect 1058 153 1086 181
rect 1098 153 1126 181
rect 1138 153 1166 181
rect 1255 153 1283 181
rect 1295 153 1323 181
rect 1335 153 1363 181
rect 73 113 101 141
rect 113 113 141 141
rect 153 113 181 141
rect 270 113 298 141
rect 310 113 338 141
rect 350 113 378 141
rect 467 113 495 141
rect 507 113 535 141
rect 547 113 575 141
rect 664 113 692 141
rect 704 113 732 141
rect 744 113 772 141
rect 861 113 889 141
rect 901 113 929 141
rect 941 113 969 141
rect 1058 113 1086 141
rect 1098 113 1126 141
rect 1138 113 1166 141
rect 1255 113 1283 141
rect 1295 113 1323 141
rect 1335 113 1363 141
rect 73 73 101 101
rect 113 73 141 101
rect 153 73 181 101
rect 270 73 298 101
rect 310 73 338 101
rect 350 73 378 101
rect 467 73 495 101
rect 507 73 535 101
rect 547 73 575 101
rect 664 73 692 101
rect 704 73 732 101
rect 744 73 772 101
rect 861 73 889 101
rect 901 73 929 101
rect 941 73 969 101
rect 1058 73 1086 101
rect 1098 73 1126 101
rect 1138 73 1166 101
rect 1255 73 1283 101
rect 1295 73 1323 101
rect 1335 73 1363 101
rect 79 32 107 33
rect 143 32 171 33
rect 79 6 103 32
rect 103 6 107 32
rect 143 6 147 32
rect 147 6 171 32
rect 79 5 107 6
rect 143 5 171 6
rect 473 32 501 33
rect 537 32 565 33
rect 473 6 497 32
rect 497 6 501 32
rect 537 6 541 32
rect 541 6 565 32
rect 473 5 501 6
rect 537 5 565 6
rect 276 -59 304 -31
rect 340 -59 368 -31
rect 867 32 895 33
rect 931 32 959 33
rect 867 6 891 32
rect 891 6 895 32
rect 931 6 935 32
rect 935 6 959 32
rect 867 5 895 6
rect 931 5 959 6
rect 670 -59 698 -31
rect 734 -59 762 -31
rect 1261 32 1289 33
rect 1325 32 1353 33
rect 1261 6 1285 32
rect 1285 6 1289 32
rect 1325 6 1329 32
rect 1329 6 1353 32
rect 1261 5 1289 6
rect 1325 5 1353 6
rect 1064 -59 1092 -31
rect 1128 -59 1156 -31
rect -176 -109 -148 -108
rect -176 -135 -175 -109
rect -175 -135 -149 -109
rect -149 -135 -148 -109
rect -176 -136 -148 -135
rect -136 -109 -108 -108
rect -136 -135 -135 -109
rect -135 -135 -109 -109
rect -109 -135 -108 -109
rect -136 -136 -108 -135
rect -96 -109 -68 -108
rect -96 -135 -95 -109
rect -95 -135 -69 -109
rect -69 -135 -68 -109
rect -96 -136 -68 -135
rect -56 -109 -28 -108
rect -56 -135 -55 -109
rect -55 -135 -29 -109
rect -29 -135 -28 -109
rect -56 -136 -28 -135
rect -16 -109 12 -108
rect -16 -135 -15 -109
rect -15 -135 11 -109
rect 11 -135 12 -109
rect -16 -136 12 -135
rect 24 -109 52 -108
rect 24 -135 25 -109
rect 25 -135 51 -109
rect 51 -135 52 -109
rect 24 -136 52 -135
rect 64 -109 92 -108
rect 64 -135 65 -109
rect 65 -135 91 -109
rect 91 -135 92 -109
rect 64 -136 92 -135
rect -176 -149 -148 -148
rect -176 -175 -175 -149
rect -175 -175 -149 -149
rect -149 -175 -148 -149
rect -176 -176 -148 -175
rect -136 -149 -108 -148
rect -136 -175 -135 -149
rect -135 -175 -109 -149
rect -109 -175 -108 -149
rect -136 -176 -108 -175
rect -96 -149 -68 -148
rect -96 -175 -95 -149
rect -95 -175 -69 -149
rect -69 -175 -68 -149
rect -96 -176 -68 -175
rect -56 -149 -28 -148
rect -56 -175 -55 -149
rect -55 -175 -29 -149
rect -29 -175 -28 -149
rect -56 -176 -28 -175
rect -16 -149 12 -148
rect -16 -175 -15 -149
rect -15 -175 11 -149
rect 11 -175 12 -149
rect -16 -176 12 -175
rect 24 -149 52 -148
rect 24 -175 25 -149
rect 25 -175 51 -149
rect 51 -175 52 -149
rect 24 -176 52 -175
rect 64 -149 92 -148
rect 64 -175 65 -149
rect 65 -175 91 -149
rect 91 -175 92 -149
rect 64 -176 92 -175
rect -176 -189 -148 -188
rect -176 -215 -175 -189
rect -175 -215 -149 -189
rect -149 -215 -148 -189
rect -176 -216 -148 -215
rect -136 -189 -108 -188
rect -136 -215 -135 -189
rect -135 -215 -109 -189
rect -109 -215 -108 -189
rect -136 -216 -108 -215
rect -96 -189 -68 -188
rect -96 -215 -95 -189
rect -95 -215 -69 -189
rect -69 -215 -68 -189
rect -96 -216 -68 -215
rect -56 -189 -28 -188
rect -56 -215 -55 -189
rect -55 -215 -29 -189
rect -29 -215 -28 -189
rect -56 -216 -28 -215
rect -16 -189 12 -188
rect -16 -215 -15 -189
rect -15 -215 11 -189
rect 11 -215 12 -189
rect -16 -216 12 -215
rect 24 -189 52 -188
rect 24 -215 25 -189
rect 25 -215 51 -189
rect 51 -215 52 -189
rect 24 -216 52 -215
rect 64 -189 92 -188
rect 64 -215 65 -189
rect 65 -215 91 -189
rect 91 -215 92 -189
rect 64 -216 92 -215
rect -176 -229 -148 -228
rect -176 -255 -175 -229
rect -175 -255 -149 -229
rect -149 -255 -148 -229
rect -176 -256 -148 -255
rect -136 -229 -108 -228
rect -136 -255 -135 -229
rect -135 -255 -109 -229
rect -109 -255 -108 -229
rect -136 -256 -108 -255
rect -96 -229 -68 -228
rect -96 -255 -95 -229
rect -95 -255 -69 -229
rect -69 -255 -68 -229
rect -96 -256 -68 -255
rect -56 -229 -28 -228
rect -56 -255 -55 -229
rect -55 -255 -29 -229
rect -29 -255 -28 -229
rect -56 -256 -28 -255
rect -16 -229 12 -228
rect -16 -255 -15 -229
rect -15 -255 11 -229
rect 11 -255 12 -229
rect -16 -256 12 -255
rect 24 -229 52 -228
rect 24 -255 25 -229
rect 25 -255 51 -229
rect 51 -255 52 -229
rect 24 -256 52 -255
rect 64 -229 92 -228
rect 64 -255 65 -229
rect 65 -255 91 -229
rect 91 -255 92 -229
rect 64 -256 92 -255
rect -176 -269 -148 -268
rect -176 -295 -175 -269
rect -175 -295 -149 -269
rect -149 -295 -148 -269
rect -176 -296 -148 -295
rect -136 -269 -108 -268
rect -136 -295 -135 -269
rect -135 -295 -109 -269
rect -109 -295 -108 -269
rect -136 -296 -108 -295
rect -96 -269 -68 -268
rect -96 -295 -95 -269
rect -95 -295 -69 -269
rect -69 -295 -68 -269
rect -96 -296 -68 -295
rect -56 -269 -28 -268
rect -56 -295 -55 -269
rect -55 -295 -29 -269
rect -29 -295 -28 -269
rect -56 -296 -28 -295
rect -16 -269 12 -268
rect -16 -295 -15 -269
rect -15 -295 11 -269
rect 11 -295 12 -269
rect -16 -296 12 -295
rect 24 -269 52 -268
rect 24 -295 25 -269
rect 25 -295 51 -269
rect 51 -295 52 -269
rect 24 -296 52 -295
rect 64 -269 92 -268
rect 64 -295 65 -269
rect 65 -295 91 -269
rect 91 -295 92 -269
rect 64 -296 92 -295
rect -176 -309 -148 -308
rect -176 -335 -175 -309
rect -175 -335 -149 -309
rect -149 -335 -148 -309
rect -176 -336 -148 -335
rect -136 -309 -108 -308
rect -136 -335 -135 -309
rect -135 -335 -109 -309
rect -109 -335 -108 -309
rect -136 -336 -108 -335
rect -96 -309 -68 -308
rect -96 -335 -95 -309
rect -95 -335 -69 -309
rect -69 -335 -68 -309
rect -96 -336 -68 -335
rect -56 -309 -28 -308
rect -56 -335 -55 -309
rect -55 -335 -29 -309
rect -29 -335 -28 -309
rect -56 -336 -28 -335
rect -16 -309 12 -308
rect -16 -335 -15 -309
rect -15 -335 11 -309
rect 11 -335 12 -309
rect -16 -336 12 -335
rect 24 -309 52 -308
rect 24 -335 25 -309
rect 25 -335 51 -309
rect 51 -335 52 -309
rect 24 -336 52 -335
rect 64 -309 92 -308
rect 64 -335 65 -309
rect 65 -335 91 -309
rect 91 -335 92 -309
rect 64 -336 92 -335
rect 582 -109 610 -108
rect 582 -135 583 -109
rect 583 -135 609 -109
rect 609 -135 610 -109
rect 582 -136 610 -135
rect 622 -109 650 -108
rect 622 -135 623 -109
rect 623 -135 649 -109
rect 649 -135 650 -109
rect 622 -136 650 -135
rect 662 -109 690 -108
rect 662 -135 663 -109
rect 663 -135 689 -109
rect 689 -135 690 -109
rect 662 -136 690 -135
rect 702 -109 730 -108
rect 702 -135 703 -109
rect 703 -135 729 -109
rect 729 -135 730 -109
rect 702 -136 730 -135
rect 742 -109 770 -108
rect 742 -135 743 -109
rect 743 -135 769 -109
rect 769 -135 770 -109
rect 742 -136 770 -135
rect 782 -109 810 -108
rect 782 -135 783 -109
rect 783 -135 809 -109
rect 809 -135 810 -109
rect 782 -136 810 -135
rect 822 -109 850 -108
rect 822 -135 823 -109
rect 823 -135 849 -109
rect 849 -135 850 -109
rect 822 -136 850 -135
rect 582 -149 610 -148
rect 582 -175 583 -149
rect 583 -175 609 -149
rect 609 -175 610 -149
rect 582 -176 610 -175
rect 622 -149 650 -148
rect 622 -175 623 -149
rect 623 -175 649 -149
rect 649 -175 650 -149
rect 622 -176 650 -175
rect 662 -149 690 -148
rect 662 -175 663 -149
rect 663 -175 689 -149
rect 689 -175 690 -149
rect 662 -176 690 -175
rect 702 -149 730 -148
rect 702 -175 703 -149
rect 703 -175 729 -149
rect 729 -175 730 -149
rect 702 -176 730 -175
rect 742 -149 770 -148
rect 742 -175 743 -149
rect 743 -175 769 -149
rect 769 -175 770 -149
rect 742 -176 770 -175
rect 782 -149 810 -148
rect 782 -175 783 -149
rect 783 -175 809 -149
rect 809 -175 810 -149
rect 782 -176 810 -175
rect 822 -149 850 -148
rect 822 -175 823 -149
rect 823 -175 849 -149
rect 849 -175 850 -149
rect 822 -176 850 -175
rect 582 -189 610 -188
rect 582 -215 583 -189
rect 583 -215 609 -189
rect 609 -215 610 -189
rect 582 -216 610 -215
rect 622 -189 650 -188
rect 622 -215 623 -189
rect 623 -215 649 -189
rect 649 -215 650 -189
rect 622 -216 650 -215
rect 662 -189 690 -188
rect 662 -215 663 -189
rect 663 -215 689 -189
rect 689 -215 690 -189
rect 662 -216 690 -215
rect 702 -189 730 -188
rect 702 -215 703 -189
rect 703 -215 729 -189
rect 729 -215 730 -189
rect 702 -216 730 -215
rect 742 -189 770 -188
rect 742 -215 743 -189
rect 743 -215 769 -189
rect 769 -215 770 -189
rect 742 -216 770 -215
rect 782 -189 810 -188
rect 782 -215 783 -189
rect 783 -215 809 -189
rect 809 -215 810 -189
rect 782 -216 810 -215
rect 822 -189 850 -188
rect 822 -215 823 -189
rect 823 -215 849 -189
rect 849 -215 850 -189
rect 822 -216 850 -215
rect 582 -229 610 -228
rect 582 -255 583 -229
rect 583 -255 609 -229
rect 609 -255 610 -229
rect 582 -256 610 -255
rect 622 -229 650 -228
rect 622 -255 623 -229
rect 623 -255 649 -229
rect 649 -255 650 -229
rect 622 -256 650 -255
rect 662 -229 690 -228
rect 662 -255 663 -229
rect 663 -255 689 -229
rect 689 -255 690 -229
rect 662 -256 690 -255
rect 702 -229 730 -228
rect 702 -255 703 -229
rect 703 -255 729 -229
rect 729 -255 730 -229
rect 702 -256 730 -255
rect 742 -229 770 -228
rect 742 -255 743 -229
rect 743 -255 769 -229
rect 769 -255 770 -229
rect 742 -256 770 -255
rect 782 -229 810 -228
rect 782 -255 783 -229
rect 783 -255 809 -229
rect 809 -255 810 -229
rect 782 -256 810 -255
rect 822 -229 850 -228
rect 822 -255 823 -229
rect 823 -255 849 -229
rect 849 -255 850 -229
rect 822 -256 850 -255
rect 582 -269 610 -268
rect 582 -295 583 -269
rect 583 -295 609 -269
rect 609 -295 610 -269
rect 582 -296 610 -295
rect 622 -269 650 -268
rect 622 -295 623 -269
rect 623 -295 649 -269
rect 649 -295 650 -269
rect 622 -296 650 -295
rect 662 -269 690 -268
rect 662 -295 663 -269
rect 663 -295 689 -269
rect 689 -295 690 -269
rect 662 -296 690 -295
rect 702 -269 730 -268
rect 702 -295 703 -269
rect 703 -295 729 -269
rect 729 -295 730 -269
rect 702 -296 730 -295
rect 742 -269 770 -268
rect 742 -295 743 -269
rect 743 -295 769 -269
rect 769 -295 770 -269
rect 742 -296 770 -295
rect 782 -269 810 -268
rect 782 -295 783 -269
rect 783 -295 809 -269
rect 809 -295 810 -269
rect 782 -296 810 -295
rect 822 -269 850 -268
rect 822 -295 823 -269
rect 823 -295 849 -269
rect 849 -295 850 -269
rect 822 -296 850 -295
rect 582 -309 610 -308
rect 582 -335 583 -309
rect 583 -335 609 -309
rect 609 -335 610 -309
rect 582 -336 610 -335
rect 622 -309 650 -308
rect 622 -335 623 -309
rect 623 -335 649 -309
rect 649 -335 650 -309
rect 622 -336 650 -335
rect 662 -309 690 -308
rect 662 -335 663 -309
rect 663 -335 689 -309
rect 689 -335 690 -309
rect 662 -336 690 -335
rect 702 -309 730 -308
rect 702 -335 703 -309
rect 703 -335 729 -309
rect 729 -335 730 -309
rect 702 -336 730 -335
rect 742 -309 770 -308
rect 742 -335 743 -309
rect 743 -335 769 -309
rect 769 -335 770 -309
rect 742 -336 770 -335
rect 782 -309 810 -308
rect 782 -335 783 -309
rect 783 -335 809 -309
rect 809 -335 810 -309
rect 782 -336 810 -335
rect 822 -309 850 -308
rect 822 -335 823 -309
rect 823 -335 849 -309
rect 849 -335 850 -309
rect 822 -336 850 -335
rect 1370 -109 1398 -108
rect 1370 -135 1371 -109
rect 1371 -135 1397 -109
rect 1397 -135 1398 -109
rect 1370 -136 1398 -135
rect 1410 -109 1438 -108
rect 1410 -135 1411 -109
rect 1411 -135 1437 -109
rect 1437 -135 1438 -109
rect 1410 -136 1438 -135
rect 1450 -109 1478 -108
rect 1450 -135 1451 -109
rect 1451 -135 1477 -109
rect 1477 -135 1478 -109
rect 1450 -136 1478 -135
rect 1490 -109 1518 -108
rect 1490 -135 1491 -109
rect 1491 -135 1517 -109
rect 1517 -135 1518 -109
rect 1490 -136 1518 -135
rect 1530 -109 1558 -108
rect 1530 -135 1531 -109
rect 1531 -135 1557 -109
rect 1557 -135 1558 -109
rect 1530 -136 1558 -135
rect 1570 -109 1598 -108
rect 1570 -135 1571 -109
rect 1571 -135 1597 -109
rect 1597 -135 1598 -109
rect 1570 -136 1598 -135
rect 1610 -109 1638 -108
rect 1610 -135 1611 -109
rect 1611 -135 1637 -109
rect 1637 -135 1638 -109
rect 1610 -136 1638 -135
rect 1370 -149 1398 -148
rect 1370 -175 1371 -149
rect 1371 -175 1397 -149
rect 1397 -175 1398 -149
rect 1370 -176 1398 -175
rect 1410 -149 1438 -148
rect 1410 -175 1411 -149
rect 1411 -175 1437 -149
rect 1437 -175 1438 -149
rect 1410 -176 1438 -175
rect 1450 -149 1478 -148
rect 1450 -175 1451 -149
rect 1451 -175 1477 -149
rect 1477 -175 1478 -149
rect 1450 -176 1478 -175
rect 1490 -149 1518 -148
rect 1490 -175 1491 -149
rect 1491 -175 1517 -149
rect 1517 -175 1518 -149
rect 1490 -176 1518 -175
rect 1530 -149 1558 -148
rect 1530 -175 1531 -149
rect 1531 -175 1557 -149
rect 1557 -175 1558 -149
rect 1530 -176 1558 -175
rect 1570 -149 1598 -148
rect 1570 -175 1571 -149
rect 1571 -175 1597 -149
rect 1597 -175 1598 -149
rect 1570 -176 1598 -175
rect 1610 -149 1638 -148
rect 1610 -175 1611 -149
rect 1611 -175 1637 -149
rect 1637 -175 1638 -149
rect 1610 -176 1638 -175
rect 1370 -189 1398 -188
rect 1370 -215 1371 -189
rect 1371 -215 1397 -189
rect 1397 -215 1398 -189
rect 1370 -216 1398 -215
rect 1410 -189 1438 -188
rect 1410 -215 1411 -189
rect 1411 -215 1437 -189
rect 1437 -215 1438 -189
rect 1410 -216 1438 -215
rect 1450 -189 1478 -188
rect 1450 -215 1451 -189
rect 1451 -215 1477 -189
rect 1477 -215 1478 -189
rect 1450 -216 1478 -215
rect 1490 -189 1518 -188
rect 1490 -215 1491 -189
rect 1491 -215 1517 -189
rect 1517 -215 1518 -189
rect 1490 -216 1518 -215
rect 1530 -189 1558 -188
rect 1530 -215 1531 -189
rect 1531 -215 1557 -189
rect 1557 -215 1558 -189
rect 1530 -216 1558 -215
rect 1570 -189 1598 -188
rect 1570 -215 1571 -189
rect 1571 -215 1597 -189
rect 1597 -215 1598 -189
rect 1570 -216 1598 -215
rect 1610 -189 1638 -188
rect 1610 -215 1611 -189
rect 1611 -215 1637 -189
rect 1637 -215 1638 -189
rect 1610 -216 1638 -215
rect 1370 -229 1398 -228
rect 1370 -255 1371 -229
rect 1371 -255 1397 -229
rect 1397 -255 1398 -229
rect 1370 -256 1398 -255
rect 1410 -229 1438 -228
rect 1410 -255 1411 -229
rect 1411 -255 1437 -229
rect 1437 -255 1438 -229
rect 1410 -256 1438 -255
rect 1450 -229 1478 -228
rect 1450 -255 1451 -229
rect 1451 -255 1477 -229
rect 1477 -255 1478 -229
rect 1450 -256 1478 -255
rect 1490 -229 1518 -228
rect 1490 -255 1491 -229
rect 1491 -255 1517 -229
rect 1517 -255 1518 -229
rect 1490 -256 1518 -255
rect 1530 -229 1558 -228
rect 1530 -255 1531 -229
rect 1531 -255 1557 -229
rect 1557 -255 1558 -229
rect 1530 -256 1558 -255
rect 1570 -229 1598 -228
rect 1570 -255 1571 -229
rect 1571 -255 1597 -229
rect 1597 -255 1598 -229
rect 1570 -256 1598 -255
rect 1610 -229 1638 -228
rect 1610 -255 1611 -229
rect 1611 -255 1637 -229
rect 1637 -255 1638 -229
rect 1610 -256 1638 -255
rect 1370 -269 1398 -268
rect 1370 -295 1371 -269
rect 1371 -295 1397 -269
rect 1397 -295 1398 -269
rect 1370 -296 1398 -295
rect 1410 -269 1438 -268
rect 1410 -295 1411 -269
rect 1411 -295 1437 -269
rect 1437 -295 1438 -269
rect 1410 -296 1438 -295
rect 1450 -269 1478 -268
rect 1450 -295 1451 -269
rect 1451 -295 1477 -269
rect 1477 -295 1478 -269
rect 1450 -296 1478 -295
rect 1490 -269 1518 -268
rect 1490 -295 1491 -269
rect 1491 -295 1517 -269
rect 1517 -295 1518 -269
rect 1490 -296 1518 -295
rect 1530 -269 1558 -268
rect 1530 -295 1531 -269
rect 1531 -295 1557 -269
rect 1557 -295 1558 -269
rect 1530 -296 1558 -295
rect 1570 -269 1598 -268
rect 1570 -295 1571 -269
rect 1571 -295 1597 -269
rect 1597 -295 1598 -269
rect 1570 -296 1598 -295
rect 1610 -269 1638 -268
rect 1610 -295 1611 -269
rect 1611 -295 1637 -269
rect 1637 -295 1638 -269
rect 1610 -296 1638 -295
rect 1370 -309 1398 -308
rect 1370 -335 1371 -309
rect 1371 -335 1397 -309
rect 1397 -335 1398 -309
rect 1370 -336 1398 -335
rect 1410 -309 1438 -308
rect 1410 -335 1411 -309
rect 1411 -335 1437 -309
rect 1437 -335 1438 -309
rect 1410 -336 1438 -335
rect 1450 -309 1478 -308
rect 1450 -335 1451 -309
rect 1451 -335 1477 -309
rect 1477 -335 1478 -309
rect 1450 -336 1478 -335
rect 1490 -309 1518 -308
rect 1490 -335 1491 -309
rect 1491 -335 1517 -309
rect 1517 -335 1518 -309
rect 1490 -336 1518 -335
rect 1530 -309 1558 -308
rect 1530 -335 1531 -309
rect 1531 -335 1557 -309
rect 1557 -335 1558 -309
rect 1530 -336 1558 -335
rect 1570 -309 1598 -308
rect 1570 -335 1571 -309
rect 1571 -335 1597 -309
rect 1597 -335 1598 -309
rect 1570 -336 1598 -335
rect 1610 -309 1638 -308
rect 1610 -335 1611 -309
rect 1611 -335 1637 -309
rect 1637 -335 1638 -309
rect 1610 -336 1638 -335
<< metal3 >>
rect 1630 1374 1720 1383
rect 1630 1342 1638 1374
rect 1670 1342 1678 1374
rect 1710 1342 1720 1374
rect 1630 1334 1720 1342
rect 1630 1327 1638 1334
rect 271 1324 1638 1327
rect 271 1296 276 1324
rect 304 1296 340 1324
rect 368 1296 670 1324
rect 698 1296 734 1324
rect 762 1296 1064 1324
rect 1092 1296 1128 1324
rect 1156 1302 1638 1324
rect 1670 1302 1678 1334
rect 1710 1302 1720 1334
rect 1156 1296 1720 1302
rect 271 1293 1720 1296
rect 74 1260 1846 1263
rect 74 1232 79 1260
rect 107 1232 143 1260
rect 171 1232 473 1260
rect 501 1232 537 1260
rect 565 1232 867 1260
rect 895 1232 931 1260
rect 959 1232 1261 1260
rect 1289 1232 1325 1260
rect 1353 1254 1846 1260
rect 1353 1232 1758 1254
rect 74 1229 1758 1232
rect 1750 1222 1758 1229
rect 1790 1222 1798 1254
rect 1830 1229 1846 1254
rect 1830 1222 1840 1229
rect 1750 1214 1840 1222
rect 70 1186 183 1188
rect 267 1186 380 1188
rect 464 1186 577 1188
rect 661 1186 774 1188
rect 858 1186 971 1188
rect 1055 1186 1168 1188
rect 1252 1186 1365 1188
rect 70 1185 184 1186
rect 70 1153 71 1185
rect 103 1153 111 1185
rect 143 1153 151 1185
rect 183 1153 184 1185
rect 70 1145 184 1153
rect 70 1113 71 1145
rect 103 1113 111 1145
rect 143 1113 151 1145
rect 183 1113 184 1145
rect 70 1105 184 1113
rect 70 1073 71 1105
rect 103 1073 111 1105
rect 143 1073 151 1105
rect 183 1073 184 1105
rect 70 1065 184 1073
rect 70 1033 71 1065
rect 103 1033 111 1065
rect 143 1033 151 1065
rect 183 1033 184 1065
rect 70 1025 184 1033
rect 70 993 71 1025
rect 103 993 111 1025
rect 143 993 151 1025
rect 183 993 184 1025
rect 70 992 184 993
rect 267 1185 381 1186
rect 267 1153 268 1185
rect 300 1153 308 1185
rect 340 1153 348 1185
rect 380 1153 381 1185
rect 267 1145 381 1153
rect 267 1113 268 1145
rect 300 1113 308 1145
rect 340 1113 348 1145
rect 380 1113 381 1145
rect 267 1105 381 1113
rect 267 1073 268 1105
rect 300 1073 308 1105
rect 340 1073 348 1105
rect 380 1073 381 1105
rect 267 1065 381 1073
rect 267 1033 268 1065
rect 300 1033 308 1065
rect 340 1033 348 1065
rect 380 1033 381 1065
rect 267 1025 381 1033
rect 267 993 268 1025
rect 300 993 308 1025
rect 340 993 348 1025
rect 380 993 381 1025
rect 267 992 381 993
rect 70 990 183 992
rect 268 990 381 992
rect 464 1185 578 1186
rect 464 1153 465 1185
rect 497 1153 505 1185
rect 537 1153 545 1185
rect 577 1153 578 1185
rect 464 1145 578 1153
rect 464 1113 465 1145
rect 497 1113 505 1145
rect 537 1113 545 1145
rect 577 1113 578 1145
rect 464 1105 578 1113
rect 464 1073 465 1105
rect 497 1073 505 1105
rect 537 1073 545 1105
rect 577 1073 578 1105
rect 464 1065 578 1073
rect 464 1033 465 1065
rect 497 1033 505 1065
rect 537 1033 545 1065
rect 577 1033 578 1065
rect 464 1025 578 1033
rect 464 993 465 1025
rect 497 993 505 1025
rect 537 993 545 1025
rect 577 993 578 1025
rect 464 992 578 993
rect 661 1185 775 1186
rect 661 1153 662 1185
rect 694 1153 702 1185
rect 734 1153 742 1185
rect 774 1153 775 1185
rect 661 1145 775 1153
rect 661 1113 662 1145
rect 694 1113 702 1145
rect 734 1113 742 1145
rect 774 1113 775 1145
rect 661 1105 775 1113
rect 661 1073 662 1105
rect 694 1073 702 1105
rect 734 1073 742 1105
rect 774 1073 775 1105
rect 661 1065 775 1073
rect 661 1033 662 1065
rect 694 1033 702 1065
rect 734 1033 742 1065
rect 774 1033 775 1065
rect 661 1025 775 1033
rect 661 993 662 1025
rect 694 993 702 1025
rect 734 993 742 1025
rect 774 993 775 1025
rect 661 992 775 993
rect 858 1185 972 1186
rect 858 1153 859 1185
rect 891 1153 899 1185
rect 931 1153 939 1185
rect 971 1153 972 1185
rect 858 1145 972 1153
rect 858 1113 859 1145
rect 891 1113 899 1145
rect 931 1113 939 1145
rect 971 1113 972 1145
rect 858 1105 972 1113
rect 858 1073 859 1105
rect 891 1073 899 1105
rect 931 1073 939 1105
rect 971 1073 972 1105
rect 858 1065 972 1073
rect 858 1033 859 1065
rect 891 1033 899 1065
rect 931 1033 939 1065
rect 971 1033 972 1065
rect 858 1025 972 1033
rect 858 993 859 1025
rect 891 993 899 1025
rect 931 993 939 1025
rect 971 993 972 1025
rect 858 992 972 993
rect 1055 1185 1169 1186
rect 1055 1153 1056 1185
rect 1088 1153 1096 1185
rect 1128 1153 1136 1185
rect 1168 1153 1169 1185
rect 1055 1145 1169 1153
rect 1055 1113 1056 1145
rect 1088 1113 1096 1145
rect 1128 1113 1136 1145
rect 1168 1113 1169 1145
rect 1055 1105 1169 1113
rect 1055 1073 1056 1105
rect 1088 1073 1096 1105
rect 1128 1073 1136 1105
rect 1168 1073 1169 1105
rect 1055 1065 1169 1073
rect 1055 1033 1056 1065
rect 1088 1033 1096 1065
rect 1128 1033 1136 1065
rect 1168 1033 1169 1065
rect 1055 1025 1169 1033
rect 1055 993 1056 1025
rect 1088 993 1096 1025
rect 1128 993 1136 1025
rect 1168 993 1169 1025
rect 1055 992 1169 993
rect 1252 1185 1366 1186
rect 1252 1153 1253 1185
rect 1285 1153 1293 1185
rect 1325 1153 1333 1185
rect 1365 1153 1366 1185
rect 1750 1182 1758 1214
rect 1790 1182 1798 1214
rect 1830 1182 1840 1214
rect 1750 1173 1840 1182
rect 1252 1145 1366 1153
rect 1252 1113 1253 1145
rect 1285 1113 1293 1145
rect 1325 1113 1333 1145
rect 1365 1113 1366 1145
rect 1252 1105 1366 1113
rect 1252 1073 1253 1105
rect 1285 1073 1293 1105
rect 1325 1073 1333 1105
rect 1365 1073 1366 1105
rect 1252 1065 1366 1073
rect 1252 1033 1253 1065
rect 1285 1033 1293 1065
rect 1325 1033 1333 1065
rect 1365 1033 1366 1065
rect 1252 1025 1366 1033
rect 1252 993 1253 1025
rect 1285 993 1293 1025
rect 1325 993 1333 1025
rect 1365 993 1366 1025
rect 1252 992 1366 993
rect 464 990 577 992
rect 661 990 774 992
rect 858 990 971 992
rect 1055 990 1168 992
rect 1252 990 1365 992
rect 70 941 1840 950
rect 70 939 1638 941
rect 70 911 73 939
rect 101 911 113 939
rect 141 911 153 939
rect 181 911 467 939
rect 495 911 507 939
rect 535 911 547 939
rect 575 911 861 939
rect 889 911 901 939
rect 929 911 941 939
rect 969 911 1255 939
rect 1283 911 1295 939
rect 1323 911 1335 939
rect 1363 911 1638 939
rect 70 909 1638 911
rect 1670 909 1678 941
rect 1710 909 1840 941
rect 70 901 1840 909
rect 70 899 1638 901
rect 70 871 73 899
rect 101 871 113 899
rect 141 871 153 899
rect 181 871 467 899
rect 495 871 507 899
rect 535 871 547 899
rect 575 871 861 899
rect 889 871 901 899
rect 929 871 941 899
rect 969 871 1255 899
rect 1283 871 1295 899
rect 1323 871 1335 899
rect 1363 871 1638 899
rect 70 869 1638 871
rect 1670 869 1678 901
rect 1710 869 1840 901
rect 70 860 1840 869
rect 70 809 1840 818
rect 70 807 1758 809
rect 70 779 270 807
rect 298 779 310 807
rect 338 779 350 807
rect 378 779 664 807
rect 692 779 704 807
rect 732 779 744 807
rect 772 779 1058 807
rect 1086 779 1098 807
rect 1126 779 1138 807
rect 1166 779 1758 807
rect 70 777 1758 779
rect 1790 777 1798 809
rect 1830 777 1840 809
rect 70 769 1840 777
rect 70 767 1758 769
rect 70 739 270 767
rect 298 739 310 767
rect 338 739 350 767
rect 378 739 664 767
rect 692 739 704 767
rect 732 739 744 767
rect 772 739 1058 767
rect 1086 739 1098 767
rect 1126 739 1138 767
rect 1166 739 1758 767
rect 70 737 1758 739
rect 1790 737 1798 769
rect 1830 737 1840 769
rect 70 729 1840 737
rect 70 728 1758 729
rect 1750 698 1758 728
rect 43 695 241 698
rect 43 667 93 695
rect 121 667 133 695
rect 161 667 241 695
rect 43 664 241 667
rect 273 695 438 698
rect 273 667 289 695
rect 317 667 329 695
rect 357 667 438 695
rect 273 664 438 667
rect 469 695 635 698
rect 469 667 487 695
rect 515 667 527 695
rect 555 667 635 695
rect 469 664 635 667
rect 667 695 832 698
rect 667 667 683 695
rect 711 667 723 695
rect 751 667 832 695
rect 667 664 832 667
rect 863 695 1029 698
rect 863 667 881 695
rect 909 667 921 695
rect 949 667 1029 695
rect 863 664 1029 667
rect 1061 695 1226 698
rect 1061 667 1077 695
rect 1105 667 1117 695
rect 1145 667 1226 695
rect 1061 664 1226 667
rect 1257 697 1758 698
rect 1790 697 1798 729
rect 1830 697 1840 729
rect 1257 695 1840 697
rect 1257 667 1275 695
rect 1303 667 1315 695
rect 1343 667 1840 695
rect 1257 664 1840 667
rect 210 599 241 664
rect 407 599 438 664
rect 604 599 635 664
rect 801 599 832 664
rect 998 599 1029 664
rect 1195 599 1226 664
rect 43 596 177 599
rect 43 568 93 596
rect 121 568 133 596
rect 161 568 177 596
rect 43 565 177 568
rect 210 596 376 599
rect 210 568 289 596
rect 317 568 329 596
rect 357 568 376 596
rect 210 565 376 568
rect 407 596 571 599
rect 407 568 487 596
rect 515 568 527 596
rect 555 568 571 596
rect 407 565 571 568
rect 604 596 770 599
rect 604 568 683 596
rect 711 568 723 596
rect 751 568 770 596
rect 604 565 770 568
rect 801 596 965 599
rect 801 568 881 596
rect 909 568 921 596
rect 949 568 965 596
rect 801 565 965 568
rect 998 596 1164 599
rect 998 568 1077 596
rect 1105 568 1117 596
rect 1145 568 1164 596
rect 998 565 1164 568
rect 1195 596 1720 599
rect 1195 568 1275 596
rect 1303 568 1315 596
rect 1343 568 1720 596
rect 1195 565 1720 568
rect 43 564 77 565
rect 1630 534 1638 565
rect 70 533 1638 534
rect 1670 533 1678 565
rect 1710 533 1720 565
rect 70 525 1720 533
rect 70 523 1638 525
rect 70 495 270 523
rect 298 495 310 523
rect 338 495 350 523
rect 378 495 664 523
rect 692 495 704 523
rect 732 495 744 523
rect 772 495 1058 523
rect 1086 495 1098 523
rect 1126 495 1138 523
rect 1166 495 1638 523
rect 70 493 1638 495
rect 1670 493 1678 525
rect 1710 493 1720 525
rect 70 485 1720 493
rect 70 483 1638 485
rect 70 455 270 483
rect 298 455 310 483
rect 338 455 350 483
rect 378 455 664 483
rect 692 455 704 483
rect 732 455 744 483
rect 772 455 1058 483
rect 1086 455 1098 483
rect 1126 455 1138 483
rect 1166 455 1638 483
rect 70 453 1638 455
rect 1670 453 1678 485
rect 1710 453 1720 485
rect 70 444 1720 453
rect 70 392 1840 401
rect 70 390 1758 392
rect 70 362 73 390
rect 101 362 113 390
rect 141 362 153 390
rect 181 362 467 390
rect 495 362 507 390
rect 535 362 547 390
rect 575 362 861 390
rect 889 362 901 390
rect 929 362 941 390
rect 969 362 1255 390
rect 1283 362 1295 390
rect 1323 362 1335 390
rect 1363 362 1758 390
rect 70 360 1758 362
rect 1790 360 1798 392
rect 1830 360 1840 392
rect 70 352 1840 360
rect 70 350 1758 352
rect 70 322 73 350
rect 101 322 113 350
rect 141 322 153 350
rect 181 322 467 350
rect 495 322 507 350
rect 535 322 547 350
rect 575 322 861 350
rect 889 322 901 350
rect 929 322 941 350
rect 969 322 1255 350
rect 1283 322 1295 350
rect 1323 322 1335 350
rect 1363 322 1758 350
rect 70 320 1758 322
rect 1790 320 1798 352
rect 1830 320 1840 352
rect 70 311 1840 320
rect 70 264 183 266
rect 267 264 380 266
rect 464 264 577 266
rect 661 264 774 266
rect 858 264 971 266
rect 1055 264 1168 266
rect 1252 264 1365 266
rect 70 263 184 264
rect 70 231 71 263
rect 103 231 111 263
rect 143 231 151 263
rect 183 231 184 263
rect 70 223 184 231
rect 70 191 71 223
rect 103 191 111 223
rect 143 191 151 223
rect 183 191 184 223
rect 70 183 184 191
rect 70 151 71 183
rect 103 151 111 183
rect 143 151 151 183
rect 183 151 184 183
rect 70 143 184 151
rect 70 111 71 143
rect 103 111 111 143
rect 143 111 151 143
rect 183 111 184 143
rect 70 103 184 111
rect 70 71 71 103
rect 103 71 111 103
rect 143 71 151 103
rect 183 71 184 103
rect 70 70 184 71
rect 267 263 381 264
rect 267 231 268 263
rect 300 231 308 263
rect 340 231 348 263
rect 380 231 381 263
rect 267 223 381 231
rect 267 191 268 223
rect 300 191 308 223
rect 340 191 348 223
rect 380 191 381 223
rect 267 183 381 191
rect 267 151 268 183
rect 300 151 308 183
rect 340 151 348 183
rect 380 151 381 183
rect 267 143 381 151
rect 267 111 268 143
rect 300 111 308 143
rect 340 111 348 143
rect 380 111 381 143
rect 267 103 381 111
rect 267 71 268 103
rect 300 71 308 103
rect 340 71 348 103
rect 380 71 381 103
rect 267 70 381 71
rect 464 263 578 264
rect 464 231 465 263
rect 497 231 505 263
rect 537 231 545 263
rect 577 231 578 263
rect 464 223 578 231
rect 464 191 465 223
rect 497 191 505 223
rect 537 191 545 223
rect 577 191 578 223
rect 464 183 578 191
rect 464 151 465 183
rect 497 151 505 183
rect 537 151 545 183
rect 577 151 578 183
rect 464 143 578 151
rect 464 111 465 143
rect 497 111 505 143
rect 537 111 545 143
rect 577 111 578 143
rect 464 103 578 111
rect 464 71 465 103
rect 497 71 505 103
rect 537 71 545 103
rect 577 71 578 103
rect 464 70 578 71
rect 661 263 775 264
rect 661 231 662 263
rect 694 231 702 263
rect 734 231 742 263
rect 774 231 775 263
rect 661 223 775 231
rect 661 191 662 223
rect 694 191 702 223
rect 734 191 742 223
rect 774 191 775 223
rect 661 183 775 191
rect 661 151 662 183
rect 694 151 702 183
rect 734 151 742 183
rect 774 151 775 183
rect 661 143 775 151
rect 661 111 662 143
rect 694 111 702 143
rect 734 111 742 143
rect 774 111 775 143
rect 661 103 775 111
rect 661 71 662 103
rect 694 71 702 103
rect 734 71 742 103
rect 774 71 775 103
rect 661 70 775 71
rect 858 263 972 264
rect 858 231 859 263
rect 891 231 899 263
rect 931 231 939 263
rect 971 231 972 263
rect 858 223 972 231
rect 858 191 859 223
rect 891 191 899 223
rect 931 191 939 223
rect 971 191 972 223
rect 858 183 972 191
rect 858 151 859 183
rect 891 151 899 183
rect 931 151 939 183
rect 971 151 972 183
rect 858 143 972 151
rect 858 111 859 143
rect 891 111 899 143
rect 931 111 939 143
rect 971 111 972 143
rect 858 103 972 111
rect 858 71 859 103
rect 891 71 899 103
rect 931 71 939 103
rect 971 71 972 103
rect 858 70 972 71
rect 1055 263 1169 264
rect 1055 231 1056 263
rect 1088 231 1096 263
rect 1128 231 1136 263
rect 1168 231 1169 263
rect 1055 223 1169 231
rect 1055 191 1056 223
rect 1088 191 1096 223
rect 1128 191 1136 223
rect 1168 191 1169 223
rect 1055 183 1169 191
rect 1055 151 1056 183
rect 1088 151 1096 183
rect 1128 151 1136 183
rect 1168 151 1169 183
rect 1055 143 1169 151
rect 1055 111 1056 143
rect 1088 111 1096 143
rect 1128 111 1136 143
rect 1168 111 1169 143
rect 1055 103 1169 111
rect 1055 71 1056 103
rect 1088 71 1096 103
rect 1128 71 1136 103
rect 1168 71 1169 103
rect 1055 70 1169 71
rect 1252 263 1366 264
rect 1252 231 1253 263
rect 1285 231 1293 263
rect 1325 231 1333 263
rect 1365 231 1366 263
rect 1252 223 1366 231
rect 1252 191 1253 223
rect 1285 191 1293 223
rect 1325 191 1333 223
rect 1365 191 1366 223
rect 1252 183 1366 191
rect 1252 151 1253 183
rect 1285 151 1293 183
rect 1325 151 1333 183
rect 1365 151 1366 183
rect 1252 143 1366 151
rect 1252 111 1253 143
rect 1285 111 1293 143
rect 1325 111 1333 143
rect 1365 111 1366 143
rect 1252 103 1366 111
rect 1252 71 1253 103
rect 1285 71 1293 103
rect 1325 71 1333 103
rect 1365 71 1366 103
rect 1252 70 1366 71
rect 1630 83 1720 92
rect 70 68 183 70
rect 267 68 380 70
rect 464 68 577 70
rect 661 68 774 70
rect 858 68 971 70
rect 1055 68 1168 70
rect 1252 68 1365 70
rect 1630 51 1638 83
rect 1670 51 1678 83
rect 1710 51 1720 83
rect 1630 43 1720 51
rect 1630 36 1638 43
rect 74 33 1638 36
rect 74 5 79 33
rect 107 5 143 33
rect 171 5 473 33
rect 501 5 537 33
rect 565 5 867 33
rect 895 5 931 33
rect 959 5 1261 33
rect 1289 5 1325 33
rect 1353 11 1638 33
rect 1670 11 1678 43
rect 1710 11 1720 43
rect 1353 5 1720 11
rect 74 2 1720 5
rect 1750 19 1840 36
rect 1750 -13 1758 19
rect 1790 -13 1798 19
rect 1830 -13 1840 19
rect 1750 -21 1840 -13
rect 1750 -28 1758 -21
rect 271 -31 1758 -28
rect 271 -59 276 -31
rect 304 -59 340 -31
rect 368 -59 670 -31
rect 698 -59 734 -31
rect 762 -59 1064 -31
rect 1092 -59 1128 -31
rect 1156 -53 1758 -31
rect 1790 -53 1798 -21
rect 1830 -53 1840 -21
rect 1156 -59 1840 -53
rect 271 -62 1840 -59
rect -193 -106 109 -103
rect -193 -138 -178 -106
rect -146 -138 -138 -106
rect -106 -138 -98 -106
rect -66 -138 -58 -106
rect -26 -138 -18 -106
rect 14 -138 22 -106
rect 54 -138 62 -106
rect 94 -138 109 -106
rect -193 -146 109 -138
rect -193 -178 -178 -146
rect -146 -178 -138 -146
rect -106 -178 -98 -146
rect -66 -178 -58 -146
rect -26 -178 -18 -146
rect 14 -178 22 -146
rect 54 -178 62 -146
rect 94 -178 109 -146
rect -193 -186 109 -178
rect -193 -218 -178 -186
rect -146 -218 -138 -186
rect -106 -218 -98 -186
rect -66 -218 -58 -186
rect -26 -218 -18 -186
rect 14 -218 22 -186
rect 54 -218 62 -186
rect 94 -218 109 -186
rect -193 -226 109 -218
rect -193 -258 -178 -226
rect -146 -258 -138 -226
rect -106 -258 -98 -226
rect -66 -258 -58 -226
rect -26 -258 -18 -226
rect 14 -258 22 -226
rect 54 -258 62 -226
rect 94 -258 109 -226
rect -193 -266 109 -258
rect -193 -298 -178 -266
rect -146 -298 -138 -266
rect -106 -298 -98 -266
rect -66 -298 -58 -266
rect -26 -298 -18 -266
rect 14 -298 22 -266
rect 54 -298 62 -266
rect 94 -298 109 -266
rect -193 -306 109 -298
rect -193 -338 -178 -306
rect -146 -338 -138 -306
rect -106 -338 -98 -306
rect -66 -338 -58 -306
rect -26 -338 -18 -306
rect 14 -338 22 -306
rect 54 -338 62 -306
rect 94 -338 109 -306
rect -193 -343 109 -338
rect 565 -106 867 -103
rect 565 -138 580 -106
rect 612 -138 620 -106
rect 652 -138 660 -106
rect 692 -138 700 -106
rect 732 -138 740 -106
rect 772 -138 780 -106
rect 812 -138 820 -106
rect 852 -138 867 -106
rect 565 -146 867 -138
rect 565 -178 580 -146
rect 612 -178 620 -146
rect 652 -178 660 -146
rect 692 -178 700 -146
rect 732 -178 740 -146
rect 772 -178 780 -146
rect 812 -178 820 -146
rect 852 -178 867 -146
rect 565 -186 867 -178
rect 565 -218 580 -186
rect 612 -218 620 -186
rect 652 -218 660 -186
rect 692 -218 700 -186
rect 732 -218 740 -186
rect 772 -218 780 -186
rect 812 -218 820 -186
rect 852 -218 867 -186
rect 565 -226 867 -218
rect 565 -258 580 -226
rect 612 -258 620 -226
rect 652 -258 660 -226
rect 692 -258 700 -226
rect 732 -258 740 -226
rect 772 -258 780 -226
rect 812 -258 820 -226
rect 852 -258 867 -226
rect 565 -266 867 -258
rect 565 -298 580 -266
rect 612 -298 620 -266
rect 652 -298 660 -266
rect 692 -298 700 -266
rect 732 -298 740 -266
rect 772 -298 780 -266
rect 812 -298 820 -266
rect 852 -298 867 -266
rect 565 -306 867 -298
rect 565 -338 580 -306
rect 612 -338 620 -306
rect 652 -338 660 -306
rect 692 -338 700 -306
rect 732 -338 740 -306
rect 772 -338 780 -306
rect 812 -338 820 -306
rect 852 -338 867 -306
rect 565 -343 867 -338
rect 1353 -106 1655 -103
rect 1353 -138 1368 -106
rect 1400 -138 1408 -106
rect 1440 -138 1448 -106
rect 1480 -138 1488 -106
rect 1520 -138 1528 -106
rect 1560 -138 1568 -106
rect 1600 -138 1608 -106
rect 1640 -138 1655 -106
rect 1353 -146 1655 -138
rect 1353 -178 1368 -146
rect 1400 -178 1408 -146
rect 1440 -178 1448 -146
rect 1480 -178 1488 -146
rect 1520 -178 1528 -146
rect 1560 -178 1568 -146
rect 1600 -178 1608 -146
rect 1640 -178 1655 -146
rect 1353 -186 1655 -178
rect 1353 -218 1368 -186
rect 1400 -218 1408 -186
rect 1440 -218 1448 -186
rect 1480 -218 1488 -186
rect 1520 -218 1528 -186
rect 1560 -218 1568 -186
rect 1600 -218 1608 -186
rect 1640 -218 1655 -186
rect 1353 -226 1655 -218
rect 1353 -258 1368 -226
rect 1400 -258 1408 -226
rect 1440 -258 1448 -226
rect 1480 -258 1488 -226
rect 1520 -258 1528 -226
rect 1560 -258 1568 -226
rect 1600 -258 1608 -226
rect 1640 -258 1655 -226
rect 1353 -266 1655 -258
rect 1353 -298 1368 -266
rect 1400 -298 1408 -266
rect 1440 -298 1448 -266
rect 1480 -298 1488 -266
rect 1520 -298 1528 -266
rect 1560 -298 1568 -266
rect 1600 -298 1608 -266
rect 1640 -298 1655 -266
rect 1353 -306 1655 -298
rect 1353 -338 1368 -306
rect 1400 -338 1408 -306
rect 1440 -338 1448 -306
rect 1480 -338 1488 -306
rect 1520 -338 1528 -306
rect 1560 -338 1568 -306
rect 1600 -338 1608 -306
rect 1640 -338 1655 -306
rect 1353 -343 1655 -338
<< via3 >>
rect 1638 1342 1670 1374
rect 1678 1342 1710 1374
rect 1638 1302 1670 1334
rect 1678 1302 1710 1334
rect 1758 1222 1790 1254
rect 1798 1222 1830 1254
rect 71 1183 103 1185
rect 71 1155 73 1183
rect 73 1155 101 1183
rect 101 1155 103 1183
rect 71 1153 103 1155
rect 111 1183 143 1185
rect 111 1155 113 1183
rect 113 1155 141 1183
rect 141 1155 143 1183
rect 111 1153 143 1155
rect 151 1183 183 1185
rect 151 1155 153 1183
rect 153 1155 181 1183
rect 181 1155 183 1183
rect 151 1153 183 1155
rect 71 1143 103 1145
rect 71 1115 73 1143
rect 73 1115 101 1143
rect 101 1115 103 1143
rect 71 1113 103 1115
rect 111 1143 143 1145
rect 111 1115 113 1143
rect 113 1115 141 1143
rect 141 1115 143 1143
rect 111 1113 143 1115
rect 151 1143 183 1145
rect 151 1115 153 1143
rect 153 1115 181 1143
rect 181 1115 183 1143
rect 151 1113 183 1115
rect 71 1103 103 1105
rect 71 1075 73 1103
rect 73 1075 101 1103
rect 101 1075 103 1103
rect 71 1073 103 1075
rect 111 1103 143 1105
rect 111 1075 113 1103
rect 113 1075 141 1103
rect 141 1075 143 1103
rect 111 1073 143 1075
rect 151 1103 183 1105
rect 151 1075 153 1103
rect 153 1075 181 1103
rect 181 1075 183 1103
rect 151 1073 183 1075
rect 71 1063 103 1065
rect 71 1035 73 1063
rect 73 1035 101 1063
rect 101 1035 103 1063
rect 71 1033 103 1035
rect 111 1063 143 1065
rect 111 1035 113 1063
rect 113 1035 141 1063
rect 141 1035 143 1063
rect 111 1033 143 1035
rect 151 1063 183 1065
rect 151 1035 153 1063
rect 153 1035 181 1063
rect 181 1035 183 1063
rect 151 1033 183 1035
rect 71 1023 103 1025
rect 71 995 73 1023
rect 73 995 101 1023
rect 101 995 103 1023
rect 71 993 103 995
rect 111 1023 143 1025
rect 111 995 113 1023
rect 113 995 141 1023
rect 141 995 143 1023
rect 111 993 143 995
rect 151 1023 183 1025
rect 151 995 153 1023
rect 153 995 181 1023
rect 181 995 183 1023
rect 151 993 183 995
rect 268 1183 300 1185
rect 268 1155 270 1183
rect 270 1155 298 1183
rect 298 1155 300 1183
rect 268 1153 300 1155
rect 308 1183 340 1185
rect 308 1155 310 1183
rect 310 1155 338 1183
rect 338 1155 340 1183
rect 308 1153 340 1155
rect 348 1183 380 1185
rect 348 1155 350 1183
rect 350 1155 378 1183
rect 378 1155 380 1183
rect 348 1153 380 1155
rect 268 1143 300 1145
rect 268 1115 270 1143
rect 270 1115 298 1143
rect 298 1115 300 1143
rect 268 1113 300 1115
rect 308 1143 340 1145
rect 308 1115 310 1143
rect 310 1115 338 1143
rect 338 1115 340 1143
rect 308 1113 340 1115
rect 348 1143 380 1145
rect 348 1115 350 1143
rect 350 1115 378 1143
rect 378 1115 380 1143
rect 348 1113 380 1115
rect 268 1103 300 1105
rect 268 1075 270 1103
rect 270 1075 298 1103
rect 298 1075 300 1103
rect 268 1073 300 1075
rect 308 1103 340 1105
rect 308 1075 310 1103
rect 310 1075 338 1103
rect 338 1075 340 1103
rect 308 1073 340 1075
rect 348 1103 380 1105
rect 348 1075 350 1103
rect 350 1075 378 1103
rect 378 1075 380 1103
rect 348 1073 380 1075
rect 268 1063 300 1065
rect 268 1035 270 1063
rect 270 1035 298 1063
rect 298 1035 300 1063
rect 268 1033 300 1035
rect 308 1063 340 1065
rect 308 1035 310 1063
rect 310 1035 338 1063
rect 338 1035 340 1063
rect 308 1033 340 1035
rect 348 1063 380 1065
rect 348 1035 350 1063
rect 350 1035 378 1063
rect 378 1035 380 1063
rect 348 1033 380 1035
rect 268 1023 300 1025
rect 268 995 270 1023
rect 270 995 298 1023
rect 298 995 300 1023
rect 268 993 300 995
rect 308 1023 340 1025
rect 308 995 310 1023
rect 310 995 338 1023
rect 338 995 340 1023
rect 308 993 340 995
rect 348 1023 380 1025
rect 348 995 350 1023
rect 350 995 378 1023
rect 378 995 380 1023
rect 348 993 380 995
rect 465 1183 497 1185
rect 465 1155 467 1183
rect 467 1155 495 1183
rect 495 1155 497 1183
rect 465 1153 497 1155
rect 505 1183 537 1185
rect 505 1155 507 1183
rect 507 1155 535 1183
rect 535 1155 537 1183
rect 505 1153 537 1155
rect 545 1183 577 1185
rect 545 1155 547 1183
rect 547 1155 575 1183
rect 575 1155 577 1183
rect 545 1153 577 1155
rect 465 1143 497 1145
rect 465 1115 467 1143
rect 467 1115 495 1143
rect 495 1115 497 1143
rect 465 1113 497 1115
rect 505 1143 537 1145
rect 505 1115 507 1143
rect 507 1115 535 1143
rect 535 1115 537 1143
rect 505 1113 537 1115
rect 545 1143 577 1145
rect 545 1115 547 1143
rect 547 1115 575 1143
rect 575 1115 577 1143
rect 545 1113 577 1115
rect 465 1103 497 1105
rect 465 1075 467 1103
rect 467 1075 495 1103
rect 495 1075 497 1103
rect 465 1073 497 1075
rect 505 1103 537 1105
rect 505 1075 507 1103
rect 507 1075 535 1103
rect 535 1075 537 1103
rect 505 1073 537 1075
rect 545 1103 577 1105
rect 545 1075 547 1103
rect 547 1075 575 1103
rect 575 1075 577 1103
rect 545 1073 577 1075
rect 465 1063 497 1065
rect 465 1035 467 1063
rect 467 1035 495 1063
rect 495 1035 497 1063
rect 465 1033 497 1035
rect 505 1063 537 1065
rect 505 1035 507 1063
rect 507 1035 535 1063
rect 535 1035 537 1063
rect 505 1033 537 1035
rect 545 1063 577 1065
rect 545 1035 547 1063
rect 547 1035 575 1063
rect 575 1035 577 1063
rect 545 1033 577 1035
rect 465 1023 497 1025
rect 465 995 467 1023
rect 467 995 495 1023
rect 495 995 497 1023
rect 465 993 497 995
rect 505 1023 537 1025
rect 505 995 507 1023
rect 507 995 535 1023
rect 535 995 537 1023
rect 505 993 537 995
rect 545 1023 577 1025
rect 545 995 547 1023
rect 547 995 575 1023
rect 575 995 577 1023
rect 545 993 577 995
rect 662 1183 694 1185
rect 662 1155 664 1183
rect 664 1155 692 1183
rect 692 1155 694 1183
rect 662 1153 694 1155
rect 702 1183 734 1185
rect 702 1155 704 1183
rect 704 1155 732 1183
rect 732 1155 734 1183
rect 702 1153 734 1155
rect 742 1183 774 1185
rect 742 1155 744 1183
rect 744 1155 772 1183
rect 772 1155 774 1183
rect 742 1153 774 1155
rect 662 1143 694 1145
rect 662 1115 664 1143
rect 664 1115 692 1143
rect 692 1115 694 1143
rect 662 1113 694 1115
rect 702 1143 734 1145
rect 702 1115 704 1143
rect 704 1115 732 1143
rect 732 1115 734 1143
rect 702 1113 734 1115
rect 742 1143 774 1145
rect 742 1115 744 1143
rect 744 1115 772 1143
rect 772 1115 774 1143
rect 742 1113 774 1115
rect 662 1103 694 1105
rect 662 1075 664 1103
rect 664 1075 692 1103
rect 692 1075 694 1103
rect 662 1073 694 1075
rect 702 1103 734 1105
rect 702 1075 704 1103
rect 704 1075 732 1103
rect 732 1075 734 1103
rect 702 1073 734 1075
rect 742 1103 774 1105
rect 742 1075 744 1103
rect 744 1075 772 1103
rect 772 1075 774 1103
rect 742 1073 774 1075
rect 662 1063 694 1065
rect 662 1035 664 1063
rect 664 1035 692 1063
rect 692 1035 694 1063
rect 662 1033 694 1035
rect 702 1063 734 1065
rect 702 1035 704 1063
rect 704 1035 732 1063
rect 732 1035 734 1063
rect 702 1033 734 1035
rect 742 1063 774 1065
rect 742 1035 744 1063
rect 744 1035 772 1063
rect 772 1035 774 1063
rect 742 1033 774 1035
rect 662 1023 694 1025
rect 662 995 664 1023
rect 664 995 692 1023
rect 692 995 694 1023
rect 662 993 694 995
rect 702 1023 734 1025
rect 702 995 704 1023
rect 704 995 732 1023
rect 732 995 734 1023
rect 702 993 734 995
rect 742 1023 774 1025
rect 742 995 744 1023
rect 744 995 772 1023
rect 772 995 774 1023
rect 742 993 774 995
rect 859 1183 891 1185
rect 859 1155 861 1183
rect 861 1155 889 1183
rect 889 1155 891 1183
rect 859 1153 891 1155
rect 899 1183 931 1185
rect 899 1155 901 1183
rect 901 1155 929 1183
rect 929 1155 931 1183
rect 899 1153 931 1155
rect 939 1183 971 1185
rect 939 1155 941 1183
rect 941 1155 969 1183
rect 969 1155 971 1183
rect 939 1153 971 1155
rect 859 1143 891 1145
rect 859 1115 861 1143
rect 861 1115 889 1143
rect 889 1115 891 1143
rect 859 1113 891 1115
rect 899 1143 931 1145
rect 899 1115 901 1143
rect 901 1115 929 1143
rect 929 1115 931 1143
rect 899 1113 931 1115
rect 939 1143 971 1145
rect 939 1115 941 1143
rect 941 1115 969 1143
rect 969 1115 971 1143
rect 939 1113 971 1115
rect 859 1103 891 1105
rect 859 1075 861 1103
rect 861 1075 889 1103
rect 889 1075 891 1103
rect 859 1073 891 1075
rect 899 1103 931 1105
rect 899 1075 901 1103
rect 901 1075 929 1103
rect 929 1075 931 1103
rect 899 1073 931 1075
rect 939 1103 971 1105
rect 939 1075 941 1103
rect 941 1075 969 1103
rect 969 1075 971 1103
rect 939 1073 971 1075
rect 859 1063 891 1065
rect 859 1035 861 1063
rect 861 1035 889 1063
rect 889 1035 891 1063
rect 859 1033 891 1035
rect 899 1063 931 1065
rect 899 1035 901 1063
rect 901 1035 929 1063
rect 929 1035 931 1063
rect 899 1033 931 1035
rect 939 1063 971 1065
rect 939 1035 941 1063
rect 941 1035 969 1063
rect 969 1035 971 1063
rect 939 1033 971 1035
rect 859 1023 891 1025
rect 859 995 861 1023
rect 861 995 889 1023
rect 889 995 891 1023
rect 859 993 891 995
rect 899 1023 931 1025
rect 899 995 901 1023
rect 901 995 929 1023
rect 929 995 931 1023
rect 899 993 931 995
rect 939 1023 971 1025
rect 939 995 941 1023
rect 941 995 969 1023
rect 969 995 971 1023
rect 939 993 971 995
rect 1056 1183 1088 1185
rect 1056 1155 1058 1183
rect 1058 1155 1086 1183
rect 1086 1155 1088 1183
rect 1056 1153 1088 1155
rect 1096 1183 1128 1185
rect 1096 1155 1098 1183
rect 1098 1155 1126 1183
rect 1126 1155 1128 1183
rect 1096 1153 1128 1155
rect 1136 1183 1168 1185
rect 1136 1155 1138 1183
rect 1138 1155 1166 1183
rect 1166 1155 1168 1183
rect 1136 1153 1168 1155
rect 1056 1143 1088 1145
rect 1056 1115 1058 1143
rect 1058 1115 1086 1143
rect 1086 1115 1088 1143
rect 1056 1113 1088 1115
rect 1096 1143 1128 1145
rect 1096 1115 1098 1143
rect 1098 1115 1126 1143
rect 1126 1115 1128 1143
rect 1096 1113 1128 1115
rect 1136 1143 1168 1145
rect 1136 1115 1138 1143
rect 1138 1115 1166 1143
rect 1166 1115 1168 1143
rect 1136 1113 1168 1115
rect 1056 1103 1088 1105
rect 1056 1075 1058 1103
rect 1058 1075 1086 1103
rect 1086 1075 1088 1103
rect 1056 1073 1088 1075
rect 1096 1103 1128 1105
rect 1096 1075 1098 1103
rect 1098 1075 1126 1103
rect 1126 1075 1128 1103
rect 1096 1073 1128 1075
rect 1136 1103 1168 1105
rect 1136 1075 1138 1103
rect 1138 1075 1166 1103
rect 1166 1075 1168 1103
rect 1136 1073 1168 1075
rect 1056 1063 1088 1065
rect 1056 1035 1058 1063
rect 1058 1035 1086 1063
rect 1086 1035 1088 1063
rect 1056 1033 1088 1035
rect 1096 1063 1128 1065
rect 1096 1035 1098 1063
rect 1098 1035 1126 1063
rect 1126 1035 1128 1063
rect 1096 1033 1128 1035
rect 1136 1063 1168 1065
rect 1136 1035 1138 1063
rect 1138 1035 1166 1063
rect 1166 1035 1168 1063
rect 1136 1033 1168 1035
rect 1056 1023 1088 1025
rect 1056 995 1058 1023
rect 1058 995 1086 1023
rect 1086 995 1088 1023
rect 1056 993 1088 995
rect 1096 1023 1128 1025
rect 1096 995 1098 1023
rect 1098 995 1126 1023
rect 1126 995 1128 1023
rect 1096 993 1128 995
rect 1136 1023 1168 1025
rect 1136 995 1138 1023
rect 1138 995 1166 1023
rect 1166 995 1168 1023
rect 1136 993 1168 995
rect 1253 1183 1285 1185
rect 1253 1155 1255 1183
rect 1255 1155 1283 1183
rect 1283 1155 1285 1183
rect 1253 1153 1285 1155
rect 1293 1183 1325 1185
rect 1293 1155 1295 1183
rect 1295 1155 1323 1183
rect 1323 1155 1325 1183
rect 1293 1153 1325 1155
rect 1333 1183 1365 1185
rect 1333 1155 1335 1183
rect 1335 1155 1363 1183
rect 1363 1155 1365 1183
rect 1333 1153 1365 1155
rect 1758 1182 1790 1214
rect 1798 1182 1830 1214
rect 1253 1143 1285 1145
rect 1253 1115 1255 1143
rect 1255 1115 1283 1143
rect 1283 1115 1285 1143
rect 1253 1113 1285 1115
rect 1293 1143 1325 1145
rect 1293 1115 1295 1143
rect 1295 1115 1323 1143
rect 1323 1115 1325 1143
rect 1293 1113 1325 1115
rect 1333 1143 1365 1145
rect 1333 1115 1335 1143
rect 1335 1115 1363 1143
rect 1363 1115 1365 1143
rect 1333 1113 1365 1115
rect 1253 1103 1285 1105
rect 1253 1075 1255 1103
rect 1255 1075 1283 1103
rect 1283 1075 1285 1103
rect 1253 1073 1285 1075
rect 1293 1103 1325 1105
rect 1293 1075 1295 1103
rect 1295 1075 1323 1103
rect 1323 1075 1325 1103
rect 1293 1073 1325 1075
rect 1333 1103 1365 1105
rect 1333 1075 1335 1103
rect 1335 1075 1363 1103
rect 1363 1075 1365 1103
rect 1333 1073 1365 1075
rect 1253 1063 1285 1065
rect 1253 1035 1255 1063
rect 1255 1035 1283 1063
rect 1283 1035 1285 1063
rect 1253 1033 1285 1035
rect 1293 1063 1325 1065
rect 1293 1035 1295 1063
rect 1295 1035 1323 1063
rect 1323 1035 1325 1063
rect 1293 1033 1325 1035
rect 1333 1063 1365 1065
rect 1333 1035 1335 1063
rect 1335 1035 1363 1063
rect 1363 1035 1365 1063
rect 1333 1033 1365 1035
rect 1253 1023 1285 1025
rect 1253 995 1255 1023
rect 1255 995 1283 1023
rect 1283 995 1285 1023
rect 1253 993 1285 995
rect 1293 1023 1325 1025
rect 1293 995 1295 1023
rect 1295 995 1323 1023
rect 1323 995 1325 1023
rect 1293 993 1325 995
rect 1333 1023 1365 1025
rect 1333 995 1335 1023
rect 1335 995 1363 1023
rect 1363 995 1365 1023
rect 1333 993 1365 995
rect 1638 909 1670 941
rect 1678 909 1710 941
rect 1638 869 1670 901
rect 1678 869 1710 901
rect 1758 777 1790 809
rect 1798 777 1830 809
rect 1758 737 1790 769
rect 1798 737 1830 769
rect 1758 697 1790 729
rect 1798 697 1830 729
rect 1638 533 1670 565
rect 1678 533 1710 565
rect 1638 493 1670 525
rect 1678 493 1710 525
rect 1638 453 1670 485
rect 1678 453 1710 485
rect 1758 360 1790 392
rect 1798 360 1830 392
rect 1758 320 1790 352
rect 1798 320 1830 352
rect 71 261 103 263
rect 71 233 73 261
rect 73 233 101 261
rect 101 233 103 261
rect 71 231 103 233
rect 111 261 143 263
rect 111 233 113 261
rect 113 233 141 261
rect 141 233 143 261
rect 111 231 143 233
rect 151 261 183 263
rect 151 233 153 261
rect 153 233 181 261
rect 181 233 183 261
rect 151 231 183 233
rect 71 221 103 223
rect 71 193 73 221
rect 73 193 101 221
rect 101 193 103 221
rect 71 191 103 193
rect 111 221 143 223
rect 111 193 113 221
rect 113 193 141 221
rect 141 193 143 221
rect 111 191 143 193
rect 151 221 183 223
rect 151 193 153 221
rect 153 193 181 221
rect 181 193 183 221
rect 151 191 183 193
rect 71 181 103 183
rect 71 153 73 181
rect 73 153 101 181
rect 101 153 103 181
rect 71 151 103 153
rect 111 181 143 183
rect 111 153 113 181
rect 113 153 141 181
rect 141 153 143 181
rect 111 151 143 153
rect 151 181 183 183
rect 151 153 153 181
rect 153 153 181 181
rect 181 153 183 181
rect 151 151 183 153
rect 71 141 103 143
rect 71 113 73 141
rect 73 113 101 141
rect 101 113 103 141
rect 71 111 103 113
rect 111 141 143 143
rect 111 113 113 141
rect 113 113 141 141
rect 141 113 143 141
rect 111 111 143 113
rect 151 141 183 143
rect 151 113 153 141
rect 153 113 181 141
rect 181 113 183 141
rect 151 111 183 113
rect 71 101 103 103
rect 71 73 73 101
rect 73 73 101 101
rect 101 73 103 101
rect 71 71 103 73
rect 111 101 143 103
rect 111 73 113 101
rect 113 73 141 101
rect 141 73 143 101
rect 111 71 143 73
rect 151 101 183 103
rect 151 73 153 101
rect 153 73 181 101
rect 181 73 183 101
rect 151 71 183 73
rect 268 261 300 263
rect 268 233 270 261
rect 270 233 298 261
rect 298 233 300 261
rect 268 231 300 233
rect 308 261 340 263
rect 308 233 310 261
rect 310 233 338 261
rect 338 233 340 261
rect 308 231 340 233
rect 348 261 380 263
rect 348 233 350 261
rect 350 233 378 261
rect 378 233 380 261
rect 348 231 380 233
rect 268 221 300 223
rect 268 193 270 221
rect 270 193 298 221
rect 298 193 300 221
rect 268 191 300 193
rect 308 221 340 223
rect 308 193 310 221
rect 310 193 338 221
rect 338 193 340 221
rect 308 191 340 193
rect 348 221 380 223
rect 348 193 350 221
rect 350 193 378 221
rect 378 193 380 221
rect 348 191 380 193
rect 268 181 300 183
rect 268 153 270 181
rect 270 153 298 181
rect 298 153 300 181
rect 268 151 300 153
rect 308 181 340 183
rect 308 153 310 181
rect 310 153 338 181
rect 338 153 340 181
rect 308 151 340 153
rect 348 181 380 183
rect 348 153 350 181
rect 350 153 378 181
rect 378 153 380 181
rect 348 151 380 153
rect 268 141 300 143
rect 268 113 270 141
rect 270 113 298 141
rect 298 113 300 141
rect 268 111 300 113
rect 308 141 340 143
rect 308 113 310 141
rect 310 113 338 141
rect 338 113 340 141
rect 308 111 340 113
rect 348 141 380 143
rect 348 113 350 141
rect 350 113 378 141
rect 378 113 380 141
rect 348 111 380 113
rect 268 101 300 103
rect 268 73 270 101
rect 270 73 298 101
rect 298 73 300 101
rect 268 71 300 73
rect 308 101 340 103
rect 308 73 310 101
rect 310 73 338 101
rect 338 73 340 101
rect 308 71 340 73
rect 348 101 380 103
rect 348 73 350 101
rect 350 73 378 101
rect 378 73 380 101
rect 348 71 380 73
rect 465 261 497 263
rect 465 233 467 261
rect 467 233 495 261
rect 495 233 497 261
rect 465 231 497 233
rect 505 261 537 263
rect 505 233 507 261
rect 507 233 535 261
rect 535 233 537 261
rect 505 231 537 233
rect 545 261 577 263
rect 545 233 547 261
rect 547 233 575 261
rect 575 233 577 261
rect 545 231 577 233
rect 465 221 497 223
rect 465 193 467 221
rect 467 193 495 221
rect 495 193 497 221
rect 465 191 497 193
rect 505 221 537 223
rect 505 193 507 221
rect 507 193 535 221
rect 535 193 537 221
rect 505 191 537 193
rect 545 221 577 223
rect 545 193 547 221
rect 547 193 575 221
rect 575 193 577 221
rect 545 191 577 193
rect 465 181 497 183
rect 465 153 467 181
rect 467 153 495 181
rect 495 153 497 181
rect 465 151 497 153
rect 505 181 537 183
rect 505 153 507 181
rect 507 153 535 181
rect 535 153 537 181
rect 505 151 537 153
rect 545 181 577 183
rect 545 153 547 181
rect 547 153 575 181
rect 575 153 577 181
rect 545 151 577 153
rect 465 141 497 143
rect 465 113 467 141
rect 467 113 495 141
rect 495 113 497 141
rect 465 111 497 113
rect 505 141 537 143
rect 505 113 507 141
rect 507 113 535 141
rect 535 113 537 141
rect 505 111 537 113
rect 545 141 577 143
rect 545 113 547 141
rect 547 113 575 141
rect 575 113 577 141
rect 545 111 577 113
rect 465 101 497 103
rect 465 73 467 101
rect 467 73 495 101
rect 495 73 497 101
rect 465 71 497 73
rect 505 101 537 103
rect 505 73 507 101
rect 507 73 535 101
rect 535 73 537 101
rect 505 71 537 73
rect 545 101 577 103
rect 545 73 547 101
rect 547 73 575 101
rect 575 73 577 101
rect 545 71 577 73
rect 662 261 694 263
rect 662 233 664 261
rect 664 233 692 261
rect 692 233 694 261
rect 662 231 694 233
rect 702 261 734 263
rect 702 233 704 261
rect 704 233 732 261
rect 732 233 734 261
rect 702 231 734 233
rect 742 261 774 263
rect 742 233 744 261
rect 744 233 772 261
rect 772 233 774 261
rect 742 231 774 233
rect 662 221 694 223
rect 662 193 664 221
rect 664 193 692 221
rect 692 193 694 221
rect 662 191 694 193
rect 702 221 734 223
rect 702 193 704 221
rect 704 193 732 221
rect 732 193 734 221
rect 702 191 734 193
rect 742 221 774 223
rect 742 193 744 221
rect 744 193 772 221
rect 772 193 774 221
rect 742 191 774 193
rect 662 181 694 183
rect 662 153 664 181
rect 664 153 692 181
rect 692 153 694 181
rect 662 151 694 153
rect 702 181 734 183
rect 702 153 704 181
rect 704 153 732 181
rect 732 153 734 181
rect 702 151 734 153
rect 742 181 774 183
rect 742 153 744 181
rect 744 153 772 181
rect 772 153 774 181
rect 742 151 774 153
rect 662 141 694 143
rect 662 113 664 141
rect 664 113 692 141
rect 692 113 694 141
rect 662 111 694 113
rect 702 141 734 143
rect 702 113 704 141
rect 704 113 732 141
rect 732 113 734 141
rect 702 111 734 113
rect 742 141 774 143
rect 742 113 744 141
rect 744 113 772 141
rect 772 113 774 141
rect 742 111 774 113
rect 662 101 694 103
rect 662 73 664 101
rect 664 73 692 101
rect 692 73 694 101
rect 662 71 694 73
rect 702 101 734 103
rect 702 73 704 101
rect 704 73 732 101
rect 732 73 734 101
rect 702 71 734 73
rect 742 101 774 103
rect 742 73 744 101
rect 744 73 772 101
rect 772 73 774 101
rect 742 71 774 73
rect 859 261 891 263
rect 859 233 861 261
rect 861 233 889 261
rect 889 233 891 261
rect 859 231 891 233
rect 899 261 931 263
rect 899 233 901 261
rect 901 233 929 261
rect 929 233 931 261
rect 899 231 931 233
rect 939 261 971 263
rect 939 233 941 261
rect 941 233 969 261
rect 969 233 971 261
rect 939 231 971 233
rect 859 221 891 223
rect 859 193 861 221
rect 861 193 889 221
rect 889 193 891 221
rect 859 191 891 193
rect 899 221 931 223
rect 899 193 901 221
rect 901 193 929 221
rect 929 193 931 221
rect 899 191 931 193
rect 939 221 971 223
rect 939 193 941 221
rect 941 193 969 221
rect 969 193 971 221
rect 939 191 971 193
rect 859 181 891 183
rect 859 153 861 181
rect 861 153 889 181
rect 889 153 891 181
rect 859 151 891 153
rect 899 181 931 183
rect 899 153 901 181
rect 901 153 929 181
rect 929 153 931 181
rect 899 151 931 153
rect 939 181 971 183
rect 939 153 941 181
rect 941 153 969 181
rect 969 153 971 181
rect 939 151 971 153
rect 859 141 891 143
rect 859 113 861 141
rect 861 113 889 141
rect 889 113 891 141
rect 859 111 891 113
rect 899 141 931 143
rect 899 113 901 141
rect 901 113 929 141
rect 929 113 931 141
rect 899 111 931 113
rect 939 141 971 143
rect 939 113 941 141
rect 941 113 969 141
rect 969 113 971 141
rect 939 111 971 113
rect 859 101 891 103
rect 859 73 861 101
rect 861 73 889 101
rect 889 73 891 101
rect 859 71 891 73
rect 899 101 931 103
rect 899 73 901 101
rect 901 73 929 101
rect 929 73 931 101
rect 899 71 931 73
rect 939 101 971 103
rect 939 73 941 101
rect 941 73 969 101
rect 969 73 971 101
rect 939 71 971 73
rect 1056 261 1088 263
rect 1056 233 1058 261
rect 1058 233 1086 261
rect 1086 233 1088 261
rect 1056 231 1088 233
rect 1096 261 1128 263
rect 1096 233 1098 261
rect 1098 233 1126 261
rect 1126 233 1128 261
rect 1096 231 1128 233
rect 1136 261 1168 263
rect 1136 233 1138 261
rect 1138 233 1166 261
rect 1166 233 1168 261
rect 1136 231 1168 233
rect 1056 221 1088 223
rect 1056 193 1058 221
rect 1058 193 1086 221
rect 1086 193 1088 221
rect 1056 191 1088 193
rect 1096 221 1128 223
rect 1096 193 1098 221
rect 1098 193 1126 221
rect 1126 193 1128 221
rect 1096 191 1128 193
rect 1136 221 1168 223
rect 1136 193 1138 221
rect 1138 193 1166 221
rect 1166 193 1168 221
rect 1136 191 1168 193
rect 1056 181 1088 183
rect 1056 153 1058 181
rect 1058 153 1086 181
rect 1086 153 1088 181
rect 1056 151 1088 153
rect 1096 181 1128 183
rect 1096 153 1098 181
rect 1098 153 1126 181
rect 1126 153 1128 181
rect 1096 151 1128 153
rect 1136 181 1168 183
rect 1136 153 1138 181
rect 1138 153 1166 181
rect 1166 153 1168 181
rect 1136 151 1168 153
rect 1056 141 1088 143
rect 1056 113 1058 141
rect 1058 113 1086 141
rect 1086 113 1088 141
rect 1056 111 1088 113
rect 1096 141 1128 143
rect 1096 113 1098 141
rect 1098 113 1126 141
rect 1126 113 1128 141
rect 1096 111 1128 113
rect 1136 141 1168 143
rect 1136 113 1138 141
rect 1138 113 1166 141
rect 1166 113 1168 141
rect 1136 111 1168 113
rect 1056 101 1088 103
rect 1056 73 1058 101
rect 1058 73 1086 101
rect 1086 73 1088 101
rect 1056 71 1088 73
rect 1096 101 1128 103
rect 1096 73 1098 101
rect 1098 73 1126 101
rect 1126 73 1128 101
rect 1096 71 1128 73
rect 1136 101 1168 103
rect 1136 73 1138 101
rect 1138 73 1166 101
rect 1166 73 1168 101
rect 1136 71 1168 73
rect 1253 261 1285 263
rect 1253 233 1255 261
rect 1255 233 1283 261
rect 1283 233 1285 261
rect 1253 231 1285 233
rect 1293 261 1325 263
rect 1293 233 1295 261
rect 1295 233 1323 261
rect 1323 233 1325 261
rect 1293 231 1325 233
rect 1333 261 1365 263
rect 1333 233 1335 261
rect 1335 233 1363 261
rect 1363 233 1365 261
rect 1333 231 1365 233
rect 1253 221 1285 223
rect 1253 193 1255 221
rect 1255 193 1283 221
rect 1283 193 1285 221
rect 1253 191 1285 193
rect 1293 221 1325 223
rect 1293 193 1295 221
rect 1295 193 1323 221
rect 1323 193 1325 221
rect 1293 191 1325 193
rect 1333 221 1365 223
rect 1333 193 1335 221
rect 1335 193 1363 221
rect 1363 193 1365 221
rect 1333 191 1365 193
rect 1253 181 1285 183
rect 1253 153 1255 181
rect 1255 153 1283 181
rect 1283 153 1285 181
rect 1253 151 1285 153
rect 1293 181 1325 183
rect 1293 153 1295 181
rect 1295 153 1323 181
rect 1323 153 1325 181
rect 1293 151 1325 153
rect 1333 181 1365 183
rect 1333 153 1335 181
rect 1335 153 1363 181
rect 1363 153 1365 181
rect 1333 151 1365 153
rect 1253 141 1285 143
rect 1253 113 1255 141
rect 1255 113 1283 141
rect 1283 113 1285 141
rect 1253 111 1285 113
rect 1293 141 1325 143
rect 1293 113 1295 141
rect 1295 113 1323 141
rect 1323 113 1325 141
rect 1293 111 1325 113
rect 1333 141 1365 143
rect 1333 113 1335 141
rect 1335 113 1363 141
rect 1363 113 1365 141
rect 1333 111 1365 113
rect 1253 101 1285 103
rect 1253 73 1255 101
rect 1255 73 1283 101
rect 1283 73 1285 101
rect 1253 71 1285 73
rect 1293 101 1325 103
rect 1293 73 1295 101
rect 1295 73 1323 101
rect 1323 73 1325 101
rect 1293 71 1325 73
rect 1333 101 1365 103
rect 1333 73 1335 101
rect 1335 73 1363 101
rect 1363 73 1365 101
rect 1333 71 1365 73
rect 1638 51 1670 83
rect 1678 51 1710 83
rect 1638 11 1670 43
rect 1678 11 1710 43
rect 1758 -13 1790 19
rect 1798 -13 1830 19
rect 1758 -53 1790 -21
rect 1798 -53 1830 -21
rect -178 -108 -146 -106
rect -178 -136 -176 -108
rect -176 -136 -148 -108
rect -148 -136 -146 -108
rect -178 -138 -146 -136
rect -138 -108 -106 -106
rect -138 -136 -136 -108
rect -136 -136 -108 -108
rect -108 -136 -106 -108
rect -138 -138 -106 -136
rect -98 -108 -66 -106
rect -98 -136 -96 -108
rect -96 -136 -68 -108
rect -68 -136 -66 -108
rect -98 -138 -66 -136
rect -58 -108 -26 -106
rect -58 -136 -56 -108
rect -56 -136 -28 -108
rect -28 -136 -26 -108
rect -58 -138 -26 -136
rect -18 -108 14 -106
rect -18 -136 -16 -108
rect -16 -136 12 -108
rect 12 -136 14 -108
rect -18 -138 14 -136
rect 22 -108 54 -106
rect 22 -136 24 -108
rect 24 -136 52 -108
rect 52 -136 54 -108
rect 22 -138 54 -136
rect 62 -108 94 -106
rect 62 -136 64 -108
rect 64 -136 92 -108
rect 92 -136 94 -108
rect 62 -138 94 -136
rect -178 -148 -146 -146
rect -178 -176 -176 -148
rect -176 -176 -148 -148
rect -148 -176 -146 -148
rect -178 -178 -146 -176
rect -138 -148 -106 -146
rect -138 -176 -136 -148
rect -136 -176 -108 -148
rect -108 -176 -106 -148
rect -138 -178 -106 -176
rect -98 -148 -66 -146
rect -98 -176 -96 -148
rect -96 -176 -68 -148
rect -68 -176 -66 -148
rect -98 -178 -66 -176
rect -58 -148 -26 -146
rect -58 -176 -56 -148
rect -56 -176 -28 -148
rect -28 -176 -26 -148
rect -58 -178 -26 -176
rect -18 -148 14 -146
rect -18 -176 -16 -148
rect -16 -176 12 -148
rect 12 -176 14 -148
rect -18 -178 14 -176
rect 22 -148 54 -146
rect 22 -176 24 -148
rect 24 -176 52 -148
rect 52 -176 54 -148
rect 22 -178 54 -176
rect 62 -148 94 -146
rect 62 -176 64 -148
rect 64 -176 92 -148
rect 92 -176 94 -148
rect 62 -178 94 -176
rect -178 -188 -146 -186
rect -178 -216 -176 -188
rect -176 -216 -148 -188
rect -148 -216 -146 -188
rect -178 -218 -146 -216
rect -138 -188 -106 -186
rect -138 -216 -136 -188
rect -136 -216 -108 -188
rect -108 -216 -106 -188
rect -138 -218 -106 -216
rect -98 -188 -66 -186
rect -98 -216 -96 -188
rect -96 -216 -68 -188
rect -68 -216 -66 -188
rect -98 -218 -66 -216
rect -58 -188 -26 -186
rect -58 -216 -56 -188
rect -56 -216 -28 -188
rect -28 -216 -26 -188
rect -58 -218 -26 -216
rect -18 -188 14 -186
rect -18 -216 -16 -188
rect -16 -216 12 -188
rect 12 -216 14 -188
rect -18 -218 14 -216
rect 22 -188 54 -186
rect 22 -216 24 -188
rect 24 -216 52 -188
rect 52 -216 54 -188
rect 22 -218 54 -216
rect 62 -188 94 -186
rect 62 -216 64 -188
rect 64 -216 92 -188
rect 92 -216 94 -188
rect 62 -218 94 -216
rect -178 -228 -146 -226
rect -178 -256 -176 -228
rect -176 -256 -148 -228
rect -148 -256 -146 -228
rect -178 -258 -146 -256
rect -138 -228 -106 -226
rect -138 -256 -136 -228
rect -136 -256 -108 -228
rect -108 -256 -106 -228
rect -138 -258 -106 -256
rect -98 -228 -66 -226
rect -98 -256 -96 -228
rect -96 -256 -68 -228
rect -68 -256 -66 -228
rect -98 -258 -66 -256
rect -58 -228 -26 -226
rect -58 -256 -56 -228
rect -56 -256 -28 -228
rect -28 -256 -26 -228
rect -58 -258 -26 -256
rect -18 -228 14 -226
rect -18 -256 -16 -228
rect -16 -256 12 -228
rect 12 -256 14 -228
rect -18 -258 14 -256
rect 22 -228 54 -226
rect 22 -256 24 -228
rect 24 -256 52 -228
rect 52 -256 54 -228
rect 22 -258 54 -256
rect 62 -228 94 -226
rect 62 -256 64 -228
rect 64 -256 92 -228
rect 92 -256 94 -228
rect 62 -258 94 -256
rect -178 -268 -146 -266
rect -178 -296 -176 -268
rect -176 -296 -148 -268
rect -148 -296 -146 -268
rect -178 -298 -146 -296
rect -138 -268 -106 -266
rect -138 -296 -136 -268
rect -136 -296 -108 -268
rect -108 -296 -106 -268
rect -138 -298 -106 -296
rect -98 -268 -66 -266
rect -98 -296 -96 -268
rect -96 -296 -68 -268
rect -68 -296 -66 -268
rect -98 -298 -66 -296
rect -58 -268 -26 -266
rect -58 -296 -56 -268
rect -56 -296 -28 -268
rect -28 -296 -26 -268
rect -58 -298 -26 -296
rect -18 -268 14 -266
rect -18 -296 -16 -268
rect -16 -296 12 -268
rect 12 -296 14 -268
rect -18 -298 14 -296
rect 22 -268 54 -266
rect 22 -296 24 -268
rect 24 -296 52 -268
rect 52 -296 54 -268
rect 22 -298 54 -296
rect 62 -268 94 -266
rect 62 -296 64 -268
rect 64 -296 92 -268
rect 92 -296 94 -268
rect 62 -298 94 -296
rect -178 -308 -146 -306
rect -178 -336 -176 -308
rect -176 -336 -148 -308
rect -148 -336 -146 -308
rect -178 -338 -146 -336
rect -138 -308 -106 -306
rect -138 -336 -136 -308
rect -136 -336 -108 -308
rect -108 -336 -106 -308
rect -138 -338 -106 -336
rect -98 -308 -66 -306
rect -98 -336 -96 -308
rect -96 -336 -68 -308
rect -68 -336 -66 -308
rect -98 -338 -66 -336
rect -58 -308 -26 -306
rect -58 -336 -56 -308
rect -56 -336 -28 -308
rect -28 -336 -26 -308
rect -58 -338 -26 -336
rect -18 -308 14 -306
rect -18 -336 -16 -308
rect -16 -336 12 -308
rect 12 -336 14 -308
rect -18 -338 14 -336
rect 22 -308 54 -306
rect 22 -336 24 -308
rect 24 -336 52 -308
rect 52 -336 54 -308
rect 22 -338 54 -336
rect 62 -308 94 -306
rect 62 -336 64 -308
rect 64 -336 92 -308
rect 92 -336 94 -308
rect 62 -338 94 -336
rect 580 -108 612 -106
rect 580 -136 582 -108
rect 582 -136 610 -108
rect 610 -136 612 -108
rect 580 -138 612 -136
rect 620 -108 652 -106
rect 620 -136 622 -108
rect 622 -136 650 -108
rect 650 -136 652 -108
rect 620 -138 652 -136
rect 660 -108 692 -106
rect 660 -136 662 -108
rect 662 -136 690 -108
rect 690 -136 692 -108
rect 660 -138 692 -136
rect 700 -108 732 -106
rect 700 -136 702 -108
rect 702 -136 730 -108
rect 730 -136 732 -108
rect 700 -138 732 -136
rect 740 -108 772 -106
rect 740 -136 742 -108
rect 742 -136 770 -108
rect 770 -136 772 -108
rect 740 -138 772 -136
rect 780 -108 812 -106
rect 780 -136 782 -108
rect 782 -136 810 -108
rect 810 -136 812 -108
rect 780 -138 812 -136
rect 820 -108 852 -106
rect 820 -136 822 -108
rect 822 -136 850 -108
rect 850 -136 852 -108
rect 820 -138 852 -136
rect 580 -148 612 -146
rect 580 -176 582 -148
rect 582 -176 610 -148
rect 610 -176 612 -148
rect 580 -178 612 -176
rect 620 -148 652 -146
rect 620 -176 622 -148
rect 622 -176 650 -148
rect 650 -176 652 -148
rect 620 -178 652 -176
rect 660 -148 692 -146
rect 660 -176 662 -148
rect 662 -176 690 -148
rect 690 -176 692 -148
rect 660 -178 692 -176
rect 700 -148 732 -146
rect 700 -176 702 -148
rect 702 -176 730 -148
rect 730 -176 732 -148
rect 700 -178 732 -176
rect 740 -148 772 -146
rect 740 -176 742 -148
rect 742 -176 770 -148
rect 770 -176 772 -148
rect 740 -178 772 -176
rect 780 -148 812 -146
rect 780 -176 782 -148
rect 782 -176 810 -148
rect 810 -176 812 -148
rect 780 -178 812 -176
rect 820 -148 852 -146
rect 820 -176 822 -148
rect 822 -176 850 -148
rect 850 -176 852 -148
rect 820 -178 852 -176
rect 580 -188 612 -186
rect 580 -216 582 -188
rect 582 -216 610 -188
rect 610 -216 612 -188
rect 580 -218 612 -216
rect 620 -188 652 -186
rect 620 -216 622 -188
rect 622 -216 650 -188
rect 650 -216 652 -188
rect 620 -218 652 -216
rect 660 -188 692 -186
rect 660 -216 662 -188
rect 662 -216 690 -188
rect 690 -216 692 -188
rect 660 -218 692 -216
rect 700 -188 732 -186
rect 700 -216 702 -188
rect 702 -216 730 -188
rect 730 -216 732 -188
rect 700 -218 732 -216
rect 740 -188 772 -186
rect 740 -216 742 -188
rect 742 -216 770 -188
rect 770 -216 772 -188
rect 740 -218 772 -216
rect 780 -188 812 -186
rect 780 -216 782 -188
rect 782 -216 810 -188
rect 810 -216 812 -188
rect 780 -218 812 -216
rect 820 -188 852 -186
rect 820 -216 822 -188
rect 822 -216 850 -188
rect 850 -216 852 -188
rect 820 -218 852 -216
rect 580 -228 612 -226
rect 580 -256 582 -228
rect 582 -256 610 -228
rect 610 -256 612 -228
rect 580 -258 612 -256
rect 620 -228 652 -226
rect 620 -256 622 -228
rect 622 -256 650 -228
rect 650 -256 652 -228
rect 620 -258 652 -256
rect 660 -228 692 -226
rect 660 -256 662 -228
rect 662 -256 690 -228
rect 690 -256 692 -228
rect 660 -258 692 -256
rect 700 -228 732 -226
rect 700 -256 702 -228
rect 702 -256 730 -228
rect 730 -256 732 -228
rect 700 -258 732 -256
rect 740 -228 772 -226
rect 740 -256 742 -228
rect 742 -256 770 -228
rect 770 -256 772 -228
rect 740 -258 772 -256
rect 780 -228 812 -226
rect 780 -256 782 -228
rect 782 -256 810 -228
rect 810 -256 812 -228
rect 780 -258 812 -256
rect 820 -228 852 -226
rect 820 -256 822 -228
rect 822 -256 850 -228
rect 850 -256 852 -228
rect 820 -258 852 -256
rect 580 -268 612 -266
rect 580 -296 582 -268
rect 582 -296 610 -268
rect 610 -296 612 -268
rect 580 -298 612 -296
rect 620 -268 652 -266
rect 620 -296 622 -268
rect 622 -296 650 -268
rect 650 -296 652 -268
rect 620 -298 652 -296
rect 660 -268 692 -266
rect 660 -296 662 -268
rect 662 -296 690 -268
rect 690 -296 692 -268
rect 660 -298 692 -296
rect 700 -268 732 -266
rect 700 -296 702 -268
rect 702 -296 730 -268
rect 730 -296 732 -268
rect 700 -298 732 -296
rect 740 -268 772 -266
rect 740 -296 742 -268
rect 742 -296 770 -268
rect 770 -296 772 -268
rect 740 -298 772 -296
rect 780 -268 812 -266
rect 780 -296 782 -268
rect 782 -296 810 -268
rect 810 -296 812 -268
rect 780 -298 812 -296
rect 820 -268 852 -266
rect 820 -296 822 -268
rect 822 -296 850 -268
rect 850 -296 852 -268
rect 820 -298 852 -296
rect 580 -308 612 -306
rect 580 -336 582 -308
rect 582 -336 610 -308
rect 610 -336 612 -308
rect 580 -338 612 -336
rect 620 -308 652 -306
rect 620 -336 622 -308
rect 622 -336 650 -308
rect 650 -336 652 -308
rect 620 -338 652 -336
rect 660 -308 692 -306
rect 660 -336 662 -308
rect 662 -336 690 -308
rect 690 -336 692 -308
rect 660 -338 692 -336
rect 700 -308 732 -306
rect 700 -336 702 -308
rect 702 -336 730 -308
rect 730 -336 732 -308
rect 700 -338 732 -336
rect 740 -308 772 -306
rect 740 -336 742 -308
rect 742 -336 770 -308
rect 770 -336 772 -308
rect 740 -338 772 -336
rect 780 -308 812 -306
rect 780 -336 782 -308
rect 782 -336 810 -308
rect 810 -336 812 -308
rect 780 -338 812 -336
rect 820 -308 852 -306
rect 820 -336 822 -308
rect 822 -336 850 -308
rect 850 -336 852 -308
rect 820 -338 852 -336
rect 1368 -108 1400 -106
rect 1368 -136 1370 -108
rect 1370 -136 1398 -108
rect 1398 -136 1400 -108
rect 1368 -138 1400 -136
rect 1408 -108 1440 -106
rect 1408 -136 1410 -108
rect 1410 -136 1438 -108
rect 1438 -136 1440 -108
rect 1408 -138 1440 -136
rect 1448 -108 1480 -106
rect 1448 -136 1450 -108
rect 1450 -136 1478 -108
rect 1478 -136 1480 -108
rect 1448 -138 1480 -136
rect 1488 -108 1520 -106
rect 1488 -136 1490 -108
rect 1490 -136 1518 -108
rect 1518 -136 1520 -108
rect 1488 -138 1520 -136
rect 1528 -108 1560 -106
rect 1528 -136 1530 -108
rect 1530 -136 1558 -108
rect 1558 -136 1560 -108
rect 1528 -138 1560 -136
rect 1568 -108 1600 -106
rect 1568 -136 1570 -108
rect 1570 -136 1598 -108
rect 1598 -136 1600 -108
rect 1568 -138 1600 -136
rect 1608 -108 1640 -106
rect 1608 -136 1610 -108
rect 1610 -136 1638 -108
rect 1638 -136 1640 -108
rect 1608 -138 1640 -136
rect 1368 -148 1400 -146
rect 1368 -176 1370 -148
rect 1370 -176 1398 -148
rect 1398 -176 1400 -148
rect 1368 -178 1400 -176
rect 1408 -148 1440 -146
rect 1408 -176 1410 -148
rect 1410 -176 1438 -148
rect 1438 -176 1440 -148
rect 1408 -178 1440 -176
rect 1448 -148 1480 -146
rect 1448 -176 1450 -148
rect 1450 -176 1478 -148
rect 1478 -176 1480 -148
rect 1448 -178 1480 -176
rect 1488 -148 1520 -146
rect 1488 -176 1490 -148
rect 1490 -176 1518 -148
rect 1518 -176 1520 -148
rect 1488 -178 1520 -176
rect 1528 -148 1560 -146
rect 1528 -176 1530 -148
rect 1530 -176 1558 -148
rect 1558 -176 1560 -148
rect 1528 -178 1560 -176
rect 1568 -148 1600 -146
rect 1568 -176 1570 -148
rect 1570 -176 1598 -148
rect 1598 -176 1600 -148
rect 1568 -178 1600 -176
rect 1608 -148 1640 -146
rect 1608 -176 1610 -148
rect 1610 -176 1638 -148
rect 1638 -176 1640 -148
rect 1608 -178 1640 -176
rect 1368 -188 1400 -186
rect 1368 -216 1370 -188
rect 1370 -216 1398 -188
rect 1398 -216 1400 -188
rect 1368 -218 1400 -216
rect 1408 -188 1440 -186
rect 1408 -216 1410 -188
rect 1410 -216 1438 -188
rect 1438 -216 1440 -188
rect 1408 -218 1440 -216
rect 1448 -188 1480 -186
rect 1448 -216 1450 -188
rect 1450 -216 1478 -188
rect 1478 -216 1480 -188
rect 1448 -218 1480 -216
rect 1488 -188 1520 -186
rect 1488 -216 1490 -188
rect 1490 -216 1518 -188
rect 1518 -216 1520 -188
rect 1488 -218 1520 -216
rect 1528 -188 1560 -186
rect 1528 -216 1530 -188
rect 1530 -216 1558 -188
rect 1558 -216 1560 -188
rect 1528 -218 1560 -216
rect 1568 -188 1600 -186
rect 1568 -216 1570 -188
rect 1570 -216 1598 -188
rect 1598 -216 1600 -188
rect 1568 -218 1600 -216
rect 1608 -188 1640 -186
rect 1608 -216 1610 -188
rect 1610 -216 1638 -188
rect 1638 -216 1640 -188
rect 1608 -218 1640 -216
rect 1368 -228 1400 -226
rect 1368 -256 1370 -228
rect 1370 -256 1398 -228
rect 1398 -256 1400 -228
rect 1368 -258 1400 -256
rect 1408 -228 1440 -226
rect 1408 -256 1410 -228
rect 1410 -256 1438 -228
rect 1438 -256 1440 -228
rect 1408 -258 1440 -256
rect 1448 -228 1480 -226
rect 1448 -256 1450 -228
rect 1450 -256 1478 -228
rect 1478 -256 1480 -228
rect 1448 -258 1480 -256
rect 1488 -228 1520 -226
rect 1488 -256 1490 -228
rect 1490 -256 1518 -228
rect 1518 -256 1520 -228
rect 1488 -258 1520 -256
rect 1528 -228 1560 -226
rect 1528 -256 1530 -228
rect 1530 -256 1558 -228
rect 1558 -256 1560 -228
rect 1528 -258 1560 -256
rect 1568 -228 1600 -226
rect 1568 -256 1570 -228
rect 1570 -256 1598 -228
rect 1598 -256 1600 -228
rect 1568 -258 1600 -256
rect 1608 -228 1640 -226
rect 1608 -256 1610 -228
rect 1610 -256 1638 -228
rect 1638 -256 1640 -228
rect 1608 -258 1640 -256
rect 1368 -268 1400 -266
rect 1368 -296 1370 -268
rect 1370 -296 1398 -268
rect 1398 -296 1400 -268
rect 1368 -298 1400 -296
rect 1408 -268 1440 -266
rect 1408 -296 1410 -268
rect 1410 -296 1438 -268
rect 1438 -296 1440 -268
rect 1408 -298 1440 -296
rect 1448 -268 1480 -266
rect 1448 -296 1450 -268
rect 1450 -296 1478 -268
rect 1478 -296 1480 -268
rect 1448 -298 1480 -296
rect 1488 -268 1520 -266
rect 1488 -296 1490 -268
rect 1490 -296 1518 -268
rect 1518 -296 1520 -268
rect 1488 -298 1520 -296
rect 1528 -268 1560 -266
rect 1528 -296 1530 -268
rect 1530 -296 1558 -268
rect 1558 -296 1560 -268
rect 1528 -298 1560 -296
rect 1568 -268 1600 -266
rect 1568 -296 1570 -268
rect 1570 -296 1598 -268
rect 1598 -296 1600 -268
rect 1568 -298 1600 -296
rect 1608 -268 1640 -266
rect 1608 -296 1610 -268
rect 1610 -296 1638 -268
rect 1638 -296 1640 -268
rect 1608 -298 1640 -296
rect 1368 -308 1400 -306
rect 1368 -336 1370 -308
rect 1370 -336 1398 -308
rect 1398 -336 1400 -308
rect 1368 -338 1400 -336
rect 1408 -308 1440 -306
rect 1408 -336 1410 -308
rect 1410 -336 1438 -308
rect 1438 -336 1440 -308
rect 1408 -338 1440 -336
rect 1448 -308 1480 -306
rect 1448 -336 1450 -308
rect 1450 -336 1478 -308
rect 1478 -336 1480 -308
rect 1448 -338 1480 -336
rect 1488 -308 1520 -306
rect 1488 -336 1490 -308
rect 1490 -336 1518 -308
rect 1518 -336 1520 -308
rect 1488 -338 1520 -336
rect 1528 -308 1560 -306
rect 1528 -336 1530 -308
rect 1530 -336 1558 -308
rect 1558 -336 1560 -308
rect 1528 -338 1560 -336
rect 1568 -308 1600 -306
rect 1568 -336 1570 -308
rect 1570 -336 1598 -308
rect 1598 -336 1600 -308
rect 1568 -338 1600 -336
rect 1608 -308 1640 -306
rect 1608 -336 1610 -308
rect 1610 -336 1638 -308
rect 1638 -336 1640 -308
rect 1608 -338 1640 -336
<< metal4 >>
rect 1630 1374 1720 1383
rect 1630 1342 1638 1374
rect 1670 1342 1678 1374
rect 1710 1342 1720 1374
rect 1630 1334 1720 1342
rect 1630 1302 1638 1334
rect 1670 1302 1678 1334
rect 1710 1302 1720 1334
rect -193 1199 200 1211
rect -193 1081 -133 1199
rect -15 1185 200 1199
rect -15 1153 71 1185
rect 103 1153 111 1185
rect 143 1153 151 1185
rect 183 1153 200 1185
rect -15 1148 200 1153
rect -15 1081 68 1148
rect -193 1039 68 1081
rect -193 921 -133 1039
rect -15 1030 68 1039
rect 186 1030 200 1148
rect -15 1025 200 1030
rect -15 993 71 1025
rect 103 993 111 1025
rect 143 993 151 1025
rect 183 993 200 1025
rect -15 975 200 993
rect 253 1185 397 1211
rect 253 1153 268 1185
rect 300 1153 308 1185
rect 340 1153 348 1185
rect 380 1153 397 1185
rect 253 1148 397 1153
rect 253 1030 265 1148
rect 383 1030 397 1148
rect 253 1025 397 1030
rect 253 993 268 1025
rect 300 993 308 1025
rect 340 993 348 1025
rect 380 993 397 1025
rect 253 975 397 993
rect 450 1185 594 1211
rect 450 1153 465 1185
rect 497 1153 505 1185
rect 537 1153 545 1185
rect 577 1153 594 1185
rect 450 1148 594 1153
rect 450 1030 462 1148
rect 580 1030 594 1148
rect 450 1025 594 1030
rect 450 993 465 1025
rect 497 993 505 1025
rect 537 993 545 1025
rect 577 993 594 1025
rect 450 975 594 993
rect 647 1185 791 1211
rect 647 1153 662 1185
rect 694 1153 702 1185
rect 734 1153 742 1185
rect 774 1153 791 1185
rect 647 1148 791 1153
rect 647 1030 659 1148
rect 777 1030 791 1148
rect 647 1025 791 1030
rect 647 993 662 1025
rect 694 993 702 1025
rect 734 993 742 1025
rect 774 993 791 1025
rect 647 975 791 993
rect 844 1185 988 1211
rect 844 1153 859 1185
rect 891 1153 899 1185
rect 931 1153 939 1185
rect 971 1153 988 1185
rect 844 1148 988 1153
rect 844 1030 856 1148
rect 974 1030 988 1148
rect 844 1025 988 1030
rect 844 993 859 1025
rect 891 993 899 1025
rect 931 993 939 1025
rect 971 993 988 1025
rect 844 975 988 993
rect 1041 1185 1185 1211
rect 1041 1153 1056 1185
rect 1088 1153 1096 1185
rect 1128 1153 1136 1185
rect 1168 1153 1185 1185
rect 1041 1148 1185 1153
rect 1041 1030 1053 1148
rect 1171 1030 1185 1148
rect 1041 1025 1185 1030
rect 1041 993 1056 1025
rect 1088 993 1096 1025
rect 1128 993 1136 1025
rect 1168 993 1185 1025
rect 1041 975 1185 993
rect 1238 1185 1382 1211
rect 1238 1153 1253 1185
rect 1285 1153 1293 1185
rect 1325 1153 1333 1185
rect 1365 1153 1382 1185
rect 1238 1148 1382 1153
rect 1238 1030 1250 1148
rect 1368 1030 1382 1148
rect 1238 1025 1382 1030
rect 1238 993 1253 1025
rect 1285 993 1293 1025
rect 1325 993 1333 1025
rect 1365 993 1382 1025
rect 1238 975 1382 993
rect -15 921 43 975
rect -193 344 43 921
rect -193 226 -133 344
rect -15 289 43 344
rect 1630 941 1720 1302
rect 1630 909 1638 941
rect 1670 909 1678 941
rect 1710 909 1720 941
rect 1630 901 1720 909
rect 1630 869 1638 901
rect 1670 869 1678 901
rect 1710 869 1720 901
rect 1630 565 1720 869
rect 1630 533 1638 565
rect 1670 533 1678 565
rect 1710 533 1720 565
rect 1630 525 1720 533
rect 1630 493 1638 525
rect 1670 493 1678 525
rect 1710 493 1720 525
rect 1630 485 1720 493
rect 1630 453 1638 485
rect 1670 453 1678 485
rect 1710 453 1720 485
rect -15 263 200 289
rect -15 231 71 263
rect 103 231 111 263
rect 143 231 151 263
rect 183 231 200 263
rect -15 226 200 231
rect -193 184 68 226
rect -193 66 -133 184
rect -15 108 68 184
rect 186 108 200 226
rect -15 103 200 108
rect -15 71 71 103
rect 103 71 111 103
rect 143 71 151 103
rect 183 71 200 103
rect -15 66 200 71
rect -193 53 200 66
rect 253 263 397 289
rect 253 231 268 263
rect 300 231 308 263
rect 340 231 348 263
rect 380 231 397 263
rect 253 226 397 231
rect 253 108 265 226
rect 383 108 397 226
rect 253 103 397 108
rect 253 71 268 103
rect 300 71 308 103
rect 340 71 348 103
rect 380 71 397 103
rect 253 53 397 71
rect 450 263 594 289
rect 450 231 465 263
rect 497 231 505 263
rect 537 231 545 263
rect 577 231 594 263
rect 450 226 594 231
rect 450 108 462 226
rect 580 108 594 226
rect 450 103 594 108
rect 450 71 465 103
rect 497 71 505 103
rect 537 71 545 103
rect 577 71 594 103
rect 450 53 594 71
rect 647 263 791 289
rect 647 231 662 263
rect 694 231 702 263
rect 734 231 742 263
rect 774 231 791 263
rect 647 226 791 231
rect 647 108 659 226
rect 777 108 791 226
rect 647 103 791 108
rect 647 71 662 103
rect 694 71 702 103
rect 734 71 742 103
rect 774 71 791 103
rect 647 53 791 71
rect 844 263 988 289
rect 844 231 859 263
rect 891 231 899 263
rect 931 231 939 263
rect 971 231 988 263
rect 844 226 988 231
rect 844 108 856 226
rect 974 108 988 226
rect 844 103 988 108
rect 844 71 859 103
rect 891 71 899 103
rect 931 71 939 103
rect 971 71 988 103
rect 844 53 988 71
rect 1041 263 1185 289
rect 1041 231 1056 263
rect 1088 231 1096 263
rect 1128 231 1136 263
rect 1168 231 1185 263
rect 1041 226 1185 231
rect 1041 108 1053 226
rect 1171 108 1185 226
rect 1041 103 1185 108
rect 1041 71 1056 103
rect 1088 71 1096 103
rect 1128 71 1136 103
rect 1168 71 1185 103
rect 1041 53 1185 71
rect 1238 263 1382 289
rect 1238 231 1253 263
rect 1285 231 1293 263
rect 1325 231 1333 263
rect 1365 231 1382 263
rect 1238 226 1382 231
rect 1238 108 1250 226
rect 1368 108 1382 226
rect 1238 103 1382 108
rect 1238 71 1253 103
rect 1285 71 1293 103
rect 1325 71 1333 103
rect 1365 71 1382 103
rect 1238 53 1382 71
rect 1630 83 1720 453
rect -193 24 43 53
rect -193 -94 -133 24
rect -15 -94 43 24
rect 1630 51 1638 83
rect 1670 51 1678 83
rect 1710 51 1720 83
rect 1630 43 1720 51
rect 1630 11 1638 43
rect 1670 11 1678 43
rect 1710 11 1720 43
rect 1630 2 1720 11
rect 1750 1254 1840 1263
rect 1750 1222 1758 1254
rect 1790 1222 1798 1254
rect 1830 1222 1840 1254
rect 1750 1214 1840 1222
rect 1750 1182 1758 1214
rect 1790 1182 1798 1214
rect 1830 1182 1840 1214
rect 1750 809 1840 1182
rect 1750 777 1758 809
rect 1790 777 1798 809
rect 1830 777 1840 809
rect 1750 769 1840 777
rect 1750 737 1758 769
rect 1790 737 1798 769
rect 1830 737 1840 769
rect 1750 729 1840 737
rect 1750 697 1758 729
rect 1790 697 1798 729
rect 1830 697 1840 729
rect 1750 392 1840 697
rect 1750 360 1758 392
rect 1790 360 1798 392
rect 1830 360 1840 392
rect 1750 352 1840 360
rect 1750 320 1758 352
rect 1790 320 1798 352
rect 1830 320 1840 352
rect 1750 19 1840 320
rect 1750 -13 1758 19
rect 1790 -13 1798 19
rect 1830 -13 1840 19
rect 1750 -21 1840 -13
rect 1750 -53 1758 -21
rect 1790 -53 1798 -21
rect 1830 -53 1840 -21
rect 1750 -62 1840 -53
rect -193 -103 43 -94
rect -193 -106 109 -103
rect -193 -138 -178 -106
rect -146 -138 -138 -106
rect -106 -136 -98 -106
rect -66 -136 -58 -106
rect -26 -136 -18 -106
rect 14 -138 22 -106
rect 54 -138 62 -106
rect 94 -138 109 -106
rect -193 -146 -133 -138
rect -15 -146 109 -138
rect -193 -178 -178 -146
rect -146 -178 -138 -146
rect 14 -178 22 -146
rect 54 -178 62 -146
rect 94 -178 109 -146
rect -193 -186 -133 -178
rect -15 -186 109 -178
rect -193 -218 -178 -186
rect -146 -218 -138 -186
rect 14 -218 22 -186
rect 54 -218 62 -186
rect 94 -218 109 -186
rect -193 -226 -133 -218
rect -15 -226 109 -218
rect -193 -258 -178 -226
rect -146 -258 -138 -226
rect -106 -258 -98 -254
rect -66 -258 -58 -254
rect -26 -258 -18 -254
rect 14 -258 22 -226
rect 54 -258 62 -226
rect 94 -258 109 -226
rect -193 -266 109 -258
rect -193 -298 -178 -266
rect -146 -298 -138 -266
rect -106 -298 -98 -266
rect -66 -298 -58 -266
rect -26 -298 -18 -266
rect 14 -298 22 -266
rect 54 -298 62 -266
rect 94 -298 109 -266
rect -193 -306 109 -298
rect -193 -338 -178 -306
rect -146 -338 -138 -306
rect -106 -338 -98 -306
rect -66 -338 -58 -306
rect -26 -338 -18 -306
rect 14 -338 22 -306
rect 54 -338 62 -306
rect 94 -338 109 -306
rect -193 -343 109 -338
rect 565 -106 867 -103
rect 565 -138 580 -106
rect 612 -138 620 -106
rect 652 -138 660 -106
rect 692 -138 700 -106
rect 732 -138 740 -106
rect 772 -138 780 -106
rect 812 -138 820 -106
rect 852 -138 867 -106
rect 565 -146 867 -138
rect 565 -166 580 -146
rect 612 -166 620 -146
rect 652 -166 660 -146
rect 692 -166 700 -146
rect 565 -284 577 -166
rect 695 -178 700 -166
rect 732 -166 740 -146
rect 772 -166 780 -146
rect 812 -166 820 -146
rect 852 -166 867 -146
rect 732 -178 737 -166
rect 695 -186 737 -178
rect 695 -218 700 -186
rect 732 -218 737 -186
rect 695 -226 737 -218
rect 695 -258 700 -226
rect 732 -258 737 -226
rect 695 -266 737 -258
rect 695 -284 700 -266
rect 565 -298 580 -284
rect 612 -298 620 -284
rect 652 -298 660 -284
rect 692 -298 700 -284
rect 732 -284 737 -266
rect 855 -284 867 -166
rect 732 -298 740 -284
rect 772 -298 780 -284
rect 812 -298 820 -284
rect 852 -298 867 -284
rect 565 -306 867 -298
rect 565 -338 580 -306
rect 612 -338 620 -306
rect 652 -338 660 -306
rect 692 -338 700 -306
rect 732 -338 740 -306
rect 772 -338 780 -306
rect 812 -338 820 -306
rect 852 -338 867 -306
rect 565 -343 867 -338
rect 1353 -106 1655 -103
rect 1353 -138 1368 -106
rect 1400 -138 1408 -106
rect 1440 -138 1448 -106
rect 1480 -138 1488 -106
rect 1520 -138 1528 -106
rect 1560 -138 1568 -106
rect 1600 -138 1608 -106
rect 1640 -138 1655 -106
rect 1353 -146 1655 -138
rect 1353 -166 1368 -146
rect 1400 -166 1408 -146
rect 1440 -166 1448 -146
rect 1480 -166 1488 -146
rect 1353 -284 1365 -166
rect 1483 -178 1488 -166
rect 1520 -166 1528 -146
rect 1560 -166 1568 -146
rect 1600 -166 1608 -146
rect 1640 -166 1655 -146
rect 1520 -178 1525 -166
rect 1483 -186 1525 -178
rect 1483 -218 1488 -186
rect 1520 -218 1525 -186
rect 1483 -226 1525 -218
rect 1483 -258 1488 -226
rect 1520 -258 1525 -226
rect 1483 -266 1525 -258
rect 1483 -284 1488 -266
rect 1353 -298 1368 -284
rect 1400 -298 1408 -284
rect 1440 -298 1448 -284
rect 1480 -298 1488 -284
rect 1520 -284 1525 -266
rect 1643 -284 1655 -166
rect 1520 -298 1528 -284
rect 1560 -298 1568 -284
rect 1600 -298 1608 -284
rect 1640 -298 1655 -284
rect 1353 -306 1655 -298
rect 1353 -338 1368 -306
rect 1400 -338 1408 -306
rect 1440 -338 1448 -306
rect 1480 -338 1488 -306
rect 1520 -338 1528 -306
rect 1560 -338 1568 -306
rect 1600 -338 1608 -306
rect 1640 -338 1655 -306
rect 1353 -343 1655 -338
<< via4 >>
rect -133 1081 -15 1199
rect 68 1145 186 1148
rect 68 1113 71 1145
rect 71 1113 103 1145
rect 103 1113 111 1145
rect 111 1113 143 1145
rect 143 1113 151 1145
rect 151 1113 183 1145
rect 183 1113 186 1145
rect 68 1105 186 1113
rect 68 1073 71 1105
rect 71 1073 103 1105
rect 103 1073 111 1105
rect 111 1073 143 1105
rect 143 1073 151 1105
rect 151 1073 183 1105
rect 183 1073 186 1105
rect 68 1065 186 1073
rect -133 921 -15 1039
rect 68 1033 71 1065
rect 71 1033 103 1065
rect 103 1033 111 1065
rect 111 1033 143 1065
rect 143 1033 151 1065
rect 151 1033 183 1065
rect 183 1033 186 1065
rect 68 1030 186 1033
rect 265 1145 383 1148
rect 265 1113 268 1145
rect 268 1113 300 1145
rect 300 1113 308 1145
rect 308 1113 340 1145
rect 340 1113 348 1145
rect 348 1113 380 1145
rect 380 1113 383 1145
rect 265 1105 383 1113
rect 265 1073 268 1105
rect 268 1073 300 1105
rect 300 1073 308 1105
rect 308 1073 340 1105
rect 340 1073 348 1105
rect 348 1073 380 1105
rect 380 1073 383 1105
rect 265 1065 383 1073
rect 265 1033 268 1065
rect 268 1033 300 1065
rect 300 1033 308 1065
rect 308 1033 340 1065
rect 340 1033 348 1065
rect 348 1033 380 1065
rect 380 1033 383 1065
rect 265 1030 383 1033
rect 462 1145 580 1148
rect 462 1113 465 1145
rect 465 1113 497 1145
rect 497 1113 505 1145
rect 505 1113 537 1145
rect 537 1113 545 1145
rect 545 1113 577 1145
rect 577 1113 580 1145
rect 462 1105 580 1113
rect 462 1073 465 1105
rect 465 1073 497 1105
rect 497 1073 505 1105
rect 505 1073 537 1105
rect 537 1073 545 1105
rect 545 1073 577 1105
rect 577 1073 580 1105
rect 462 1065 580 1073
rect 462 1033 465 1065
rect 465 1033 497 1065
rect 497 1033 505 1065
rect 505 1033 537 1065
rect 537 1033 545 1065
rect 545 1033 577 1065
rect 577 1033 580 1065
rect 462 1030 580 1033
rect 659 1145 777 1148
rect 659 1113 662 1145
rect 662 1113 694 1145
rect 694 1113 702 1145
rect 702 1113 734 1145
rect 734 1113 742 1145
rect 742 1113 774 1145
rect 774 1113 777 1145
rect 659 1105 777 1113
rect 659 1073 662 1105
rect 662 1073 694 1105
rect 694 1073 702 1105
rect 702 1073 734 1105
rect 734 1073 742 1105
rect 742 1073 774 1105
rect 774 1073 777 1105
rect 659 1065 777 1073
rect 659 1033 662 1065
rect 662 1033 694 1065
rect 694 1033 702 1065
rect 702 1033 734 1065
rect 734 1033 742 1065
rect 742 1033 774 1065
rect 774 1033 777 1065
rect 659 1030 777 1033
rect 856 1145 974 1148
rect 856 1113 859 1145
rect 859 1113 891 1145
rect 891 1113 899 1145
rect 899 1113 931 1145
rect 931 1113 939 1145
rect 939 1113 971 1145
rect 971 1113 974 1145
rect 856 1105 974 1113
rect 856 1073 859 1105
rect 859 1073 891 1105
rect 891 1073 899 1105
rect 899 1073 931 1105
rect 931 1073 939 1105
rect 939 1073 971 1105
rect 971 1073 974 1105
rect 856 1065 974 1073
rect 856 1033 859 1065
rect 859 1033 891 1065
rect 891 1033 899 1065
rect 899 1033 931 1065
rect 931 1033 939 1065
rect 939 1033 971 1065
rect 971 1033 974 1065
rect 856 1030 974 1033
rect 1053 1145 1171 1148
rect 1053 1113 1056 1145
rect 1056 1113 1088 1145
rect 1088 1113 1096 1145
rect 1096 1113 1128 1145
rect 1128 1113 1136 1145
rect 1136 1113 1168 1145
rect 1168 1113 1171 1145
rect 1053 1105 1171 1113
rect 1053 1073 1056 1105
rect 1056 1073 1088 1105
rect 1088 1073 1096 1105
rect 1096 1073 1128 1105
rect 1128 1073 1136 1105
rect 1136 1073 1168 1105
rect 1168 1073 1171 1105
rect 1053 1065 1171 1073
rect 1053 1033 1056 1065
rect 1056 1033 1088 1065
rect 1088 1033 1096 1065
rect 1096 1033 1128 1065
rect 1128 1033 1136 1065
rect 1136 1033 1168 1065
rect 1168 1033 1171 1065
rect 1053 1030 1171 1033
rect 1250 1145 1368 1148
rect 1250 1113 1253 1145
rect 1253 1113 1285 1145
rect 1285 1113 1293 1145
rect 1293 1113 1325 1145
rect 1325 1113 1333 1145
rect 1333 1113 1365 1145
rect 1365 1113 1368 1145
rect 1250 1105 1368 1113
rect 1250 1073 1253 1105
rect 1253 1073 1285 1105
rect 1285 1073 1293 1105
rect 1293 1073 1325 1105
rect 1325 1073 1333 1105
rect 1333 1073 1365 1105
rect 1365 1073 1368 1105
rect 1250 1065 1368 1073
rect 1250 1033 1253 1065
rect 1253 1033 1285 1065
rect 1285 1033 1293 1065
rect 1293 1033 1325 1065
rect 1325 1033 1333 1065
rect 1333 1033 1365 1065
rect 1365 1033 1368 1065
rect 1250 1030 1368 1033
rect -133 226 -15 344
rect 68 223 186 226
rect 68 191 71 223
rect 71 191 103 223
rect 103 191 111 223
rect 111 191 143 223
rect 143 191 151 223
rect 151 191 183 223
rect 183 191 186 223
rect -133 66 -15 184
rect 68 183 186 191
rect 68 151 71 183
rect 71 151 103 183
rect 103 151 111 183
rect 111 151 143 183
rect 143 151 151 183
rect 151 151 183 183
rect 183 151 186 183
rect 68 143 186 151
rect 68 111 71 143
rect 71 111 103 143
rect 103 111 111 143
rect 111 111 143 143
rect 143 111 151 143
rect 151 111 183 143
rect 183 111 186 143
rect 68 108 186 111
rect 265 223 383 226
rect 265 191 268 223
rect 268 191 300 223
rect 300 191 308 223
rect 308 191 340 223
rect 340 191 348 223
rect 348 191 380 223
rect 380 191 383 223
rect 265 183 383 191
rect 265 151 268 183
rect 268 151 300 183
rect 300 151 308 183
rect 308 151 340 183
rect 340 151 348 183
rect 348 151 380 183
rect 380 151 383 183
rect 265 143 383 151
rect 265 111 268 143
rect 268 111 300 143
rect 300 111 308 143
rect 308 111 340 143
rect 340 111 348 143
rect 348 111 380 143
rect 380 111 383 143
rect 265 108 383 111
rect 462 223 580 226
rect 462 191 465 223
rect 465 191 497 223
rect 497 191 505 223
rect 505 191 537 223
rect 537 191 545 223
rect 545 191 577 223
rect 577 191 580 223
rect 462 183 580 191
rect 462 151 465 183
rect 465 151 497 183
rect 497 151 505 183
rect 505 151 537 183
rect 537 151 545 183
rect 545 151 577 183
rect 577 151 580 183
rect 462 143 580 151
rect 462 111 465 143
rect 465 111 497 143
rect 497 111 505 143
rect 505 111 537 143
rect 537 111 545 143
rect 545 111 577 143
rect 577 111 580 143
rect 462 108 580 111
rect 659 223 777 226
rect 659 191 662 223
rect 662 191 694 223
rect 694 191 702 223
rect 702 191 734 223
rect 734 191 742 223
rect 742 191 774 223
rect 774 191 777 223
rect 659 183 777 191
rect 659 151 662 183
rect 662 151 694 183
rect 694 151 702 183
rect 702 151 734 183
rect 734 151 742 183
rect 742 151 774 183
rect 774 151 777 183
rect 659 143 777 151
rect 659 111 662 143
rect 662 111 694 143
rect 694 111 702 143
rect 702 111 734 143
rect 734 111 742 143
rect 742 111 774 143
rect 774 111 777 143
rect 659 108 777 111
rect 856 223 974 226
rect 856 191 859 223
rect 859 191 891 223
rect 891 191 899 223
rect 899 191 931 223
rect 931 191 939 223
rect 939 191 971 223
rect 971 191 974 223
rect 856 183 974 191
rect 856 151 859 183
rect 859 151 891 183
rect 891 151 899 183
rect 899 151 931 183
rect 931 151 939 183
rect 939 151 971 183
rect 971 151 974 183
rect 856 143 974 151
rect 856 111 859 143
rect 859 111 891 143
rect 891 111 899 143
rect 899 111 931 143
rect 931 111 939 143
rect 939 111 971 143
rect 971 111 974 143
rect 856 108 974 111
rect 1053 223 1171 226
rect 1053 191 1056 223
rect 1056 191 1088 223
rect 1088 191 1096 223
rect 1096 191 1128 223
rect 1128 191 1136 223
rect 1136 191 1168 223
rect 1168 191 1171 223
rect 1053 183 1171 191
rect 1053 151 1056 183
rect 1056 151 1088 183
rect 1088 151 1096 183
rect 1096 151 1128 183
rect 1128 151 1136 183
rect 1136 151 1168 183
rect 1168 151 1171 183
rect 1053 143 1171 151
rect 1053 111 1056 143
rect 1056 111 1088 143
rect 1088 111 1096 143
rect 1096 111 1128 143
rect 1128 111 1136 143
rect 1136 111 1168 143
rect 1168 111 1171 143
rect 1053 108 1171 111
rect 1250 223 1368 226
rect 1250 191 1253 223
rect 1253 191 1285 223
rect 1285 191 1293 223
rect 1293 191 1325 223
rect 1325 191 1333 223
rect 1333 191 1365 223
rect 1365 191 1368 223
rect 1250 183 1368 191
rect 1250 151 1253 183
rect 1253 151 1285 183
rect 1285 151 1293 183
rect 1293 151 1325 183
rect 1325 151 1333 183
rect 1333 151 1365 183
rect 1365 151 1368 183
rect 1250 143 1368 151
rect 1250 111 1253 143
rect 1253 111 1285 143
rect 1285 111 1293 143
rect 1293 111 1325 143
rect 1325 111 1333 143
rect 1333 111 1365 143
rect 1365 111 1368 143
rect 1250 108 1368 111
rect -133 -94 -15 24
rect -133 -138 -106 -136
rect -106 -138 -98 -136
rect -98 -138 -66 -136
rect -66 -138 -58 -136
rect -58 -138 -26 -136
rect -26 -138 -18 -136
rect -18 -138 -15 -136
rect -133 -146 -15 -138
rect -133 -178 -106 -146
rect -106 -178 -98 -146
rect -98 -178 -66 -146
rect -66 -178 -58 -146
rect -58 -178 -26 -146
rect -26 -178 -18 -146
rect -18 -178 -15 -146
rect -133 -186 -15 -178
rect -133 -218 -106 -186
rect -106 -218 -98 -186
rect -98 -218 -66 -186
rect -66 -218 -58 -186
rect -58 -218 -26 -186
rect -26 -218 -18 -186
rect -18 -218 -15 -186
rect -133 -226 -15 -218
rect -133 -254 -106 -226
rect -106 -254 -98 -226
rect -98 -254 -66 -226
rect -66 -254 -58 -226
rect -58 -254 -26 -226
rect -26 -254 -18 -226
rect -18 -254 -15 -226
rect 577 -178 580 -166
rect 580 -178 612 -166
rect 612 -178 620 -166
rect 620 -178 652 -166
rect 652 -178 660 -166
rect 660 -178 692 -166
rect 692 -178 695 -166
rect 737 -178 740 -166
rect 740 -178 772 -166
rect 772 -178 780 -166
rect 780 -178 812 -166
rect 812 -178 820 -166
rect 820 -178 852 -166
rect 852 -178 855 -166
rect 577 -186 695 -178
rect 737 -186 855 -178
rect 577 -218 580 -186
rect 580 -218 612 -186
rect 612 -218 620 -186
rect 620 -218 652 -186
rect 652 -218 660 -186
rect 660 -218 692 -186
rect 692 -218 695 -186
rect 737 -218 740 -186
rect 740 -218 772 -186
rect 772 -218 780 -186
rect 780 -218 812 -186
rect 812 -218 820 -186
rect 820 -218 852 -186
rect 852 -218 855 -186
rect 577 -226 695 -218
rect 737 -226 855 -218
rect 577 -258 580 -226
rect 580 -258 612 -226
rect 612 -258 620 -226
rect 620 -258 652 -226
rect 652 -258 660 -226
rect 660 -258 692 -226
rect 692 -258 695 -226
rect 737 -258 740 -226
rect 740 -258 772 -226
rect 772 -258 780 -226
rect 780 -258 812 -226
rect 812 -258 820 -226
rect 820 -258 852 -226
rect 852 -258 855 -226
rect 577 -266 695 -258
rect 737 -266 855 -258
rect 577 -284 580 -266
rect 580 -284 612 -266
rect 612 -284 620 -266
rect 620 -284 652 -266
rect 652 -284 660 -266
rect 660 -284 692 -266
rect 692 -284 695 -266
rect 737 -284 740 -266
rect 740 -284 772 -266
rect 772 -284 780 -266
rect 780 -284 812 -266
rect 812 -284 820 -266
rect 820 -284 852 -266
rect 852 -284 855 -266
rect 1365 -178 1368 -166
rect 1368 -178 1400 -166
rect 1400 -178 1408 -166
rect 1408 -178 1440 -166
rect 1440 -178 1448 -166
rect 1448 -178 1480 -166
rect 1480 -178 1483 -166
rect 1525 -178 1528 -166
rect 1528 -178 1560 -166
rect 1560 -178 1568 -166
rect 1568 -178 1600 -166
rect 1600 -178 1608 -166
rect 1608 -178 1640 -166
rect 1640 -178 1643 -166
rect 1365 -186 1483 -178
rect 1525 -186 1643 -178
rect 1365 -218 1368 -186
rect 1368 -218 1400 -186
rect 1400 -218 1408 -186
rect 1408 -218 1440 -186
rect 1440 -218 1448 -186
rect 1448 -218 1480 -186
rect 1480 -218 1483 -186
rect 1525 -218 1528 -186
rect 1528 -218 1560 -186
rect 1560 -218 1568 -186
rect 1568 -218 1600 -186
rect 1600 -218 1608 -186
rect 1608 -218 1640 -186
rect 1640 -218 1643 -186
rect 1365 -226 1483 -218
rect 1525 -226 1643 -218
rect 1365 -258 1368 -226
rect 1368 -258 1400 -226
rect 1400 -258 1408 -226
rect 1408 -258 1440 -226
rect 1440 -258 1448 -226
rect 1448 -258 1480 -226
rect 1480 -258 1483 -226
rect 1525 -258 1528 -226
rect 1528 -258 1560 -226
rect 1560 -258 1568 -226
rect 1568 -258 1600 -226
rect 1600 -258 1608 -226
rect 1608 -258 1640 -226
rect 1640 -258 1643 -226
rect 1365 -266 1483 -258
rect 1525 -266 1643 -258
rect 1365 -284 1368 -266
rect 1368 -284 1400 -266
rect 1400 -284 1408 -266
rect 1408 -284 1440 -266
rect 1440 -284 1448 -266
rect 1448 -284 1480 -266
rect 1480 -284 1483 -266
rect 1525 -284 1528 -266
rect 1528 -284 1560 -266
rect 1560 -284 1568 -266
rect 1568 -284 1600 -266
rect 1600 -284 1608 -266
rect 1608 -284 1640 -266
rect 1640 -284 1643 -266
<< metal5 >>
rect -193 1199 1393 1211
rect -193 1081 -133 1199
rect -15 1148 1393 1199
rect -15 1081 68 1148
rect -193 1039 68 1081
rect -193 921 -133 1039
rect -15 1030 68 1039
rect 186 1030 265 1148
rect 383 1030 462 1148
rect 580 1030 659 1148
rect 777 1030 856 1148
rect 974 1030 1053 1148
rect 1171 1030 1250 1148
rect 1368 1030 1393 1148
rect -15 975 1393 1030
rect -15 921 43 975
rect -193 908 43 921
rect -193 344 43 356
rect -193 226 -133 344
rect -15 289 43 344
rect -15 226 1393 289
rect -193 184 68 226
rect -193 66 -133 184
rect -15 108 68 184
rect 186 108 265 226
rect 383 108 462 226
rect 580 108 659 226
rect 777 108 856 226
rect 974 108 1053 226
rect 1171 108 1250 226
rect 1368 108 1393 226
rect -15 66 1393 108
rect -193 53 1393 66
rect -193 24 43 53
rect -193 -94 -133 24
rect -15 -94 43 24
rect -193 -107 43 -94
rect -193 -136 1840 -107
rect -193 -254 -133 -136
rect -15 -166 1840 -136
rect -15 -254 577 -166
rect -193 -284 577 -254
rect 695 -284 737 -166
rect 855 -284 1365 -166
rect 1483 -284 1525 -166
rect 1643 -284 1840 -166
rect -193 -343 1840 -284
use vco_pair_base  vco_pair_base_0
timestamp 1654635176
transform 1 0 -1 0 1 666
box -197 -707 1631 640
<< labels >>
flabel metal5 s 247 -242 253 -226 0 FreeSans 800 0 0 0 GND
port 0 nsew
flabel metal3 s 1819 896 1825 912 0 FreeSans 800 0 0 0 OUT_P
port 1 nsew
flabel metal3 s 1826 766 1832 782 0 FreeSans 800 0 0 0 OUT_N
port 3 nsew
<< end >>
