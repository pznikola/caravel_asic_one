magic
tech sky130B
magscale 1 2
timestamp 1654038913
<< metal3 >>
rect -480 402 479 430
rect -480 -402 395 402
rect 459 -402 479 402
rect -480 -430 479 -402
<< via3 >>
rect 395 -402 459 402
<< mimcap >>
rect -380 290 280 330
rect -380 -290 -340 290
rect 240 -290 280 290
rect -380 -330 280 -290
<< mimcapcontact >>
rect -340 -290 240 290
<< metal4 >>
rect 379 402 475 418
rect -341 290 241 291
rect -341 -290 -340 290
rect 240 -290 241 290
rect -341 -291 241 -290
rect 379 -402 395 402
rect 459 -402 475 402
rect 379 -418 475 -402
<< properties >>
string FIXED_BBOX -480 -430 380 430
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.3 l 3.3 val 24.287 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
