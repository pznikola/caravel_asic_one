* NGSPICE file created from vco_pmirr_pex.ext - technology: sky130B

.subckt vco_pmirr_pex VBIAS IND_CT VDD GND
X0 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t4 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t3 VDD.t66 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X1 VDD VDD.t37 VDD VDD.t1 sky130_fd_pr__pfet_01v8 ad=2.78124e+13p pd=2.1714e+08u as=0p ps=0u w=3.01e+06u l=150000u
X2 VDD.t65 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t5 IND_CT.t15 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X3 VDD.t36 VDD.t34 VDD.t35 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X4 VDD.t33 VDD.t30 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X5 IND_CT.t14 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t6 VDD.t64 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X6 VDD VDD.t25 VDD VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X7 VDD.t63 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t1 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t2 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X8 IND_CT.t13 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t7 VDD.t62 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X9 IND_CT.t12 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t8 VDD.t61 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X10 VDD VDD.t21 VDD VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X11 VBIAS.t0 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t0 GND.t0 sky130_fd_pr__res_high_po_2p85 l=3.5e+06u
X12 IND_CT.t11 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t9 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X13 VDD.t58 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t10 IND_CT.t10 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X14 VDD.t57 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t11 IND_CT.t9 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X15 IND_CT.t8 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t12 VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X16 VDD.t54 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t13 IND_CT.t7 VDD.t53 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X17 VDD.t51 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t14 IND_CT.t6 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X18 VDD.t52 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t15 IND_CT.t5 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X19 VDD.t49 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t16 IND_CT.t4 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X20 VDD.t20 VDD.t17 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X21 VDD.t47 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t17 IND_CT.t3 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X22 IND_CT.t2 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t18 VDD.t45 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X23 VDD VDD.t12 VDD VDD.t13 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X24 VDD.t11 VDD.t9 VDD.t10 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X25 IND_CT.t1 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t19 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X26 IND_CT.t0 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t20 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X27 VDD.t8 VDD.t5 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
X28 VDD VDD.t0 VDD VDD.t1 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
C0 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE IND_CT 9.77fF
C1 VDD VBIAS 0.52fF
C2 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE VBIAS 0.69fF
C3 VDD vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE 22.87fF
C4 IND_CT VBIAS 0.01fF
C5 VDD IND_CT 23.96fF
R0 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n54 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t3 535.019
R1 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n67 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t1 535.019
R2 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n943 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t15 535.019
R3 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n964 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t6 535.019
R4 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n905 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t5 535.019
R5 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n926 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t19 535.019
R6 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1000 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t12 535.019
R7 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n981 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t17 535.019
R8 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n438 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t16 535.019
R9 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n459 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t20 535.019
R10 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n385 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t13 535.019
R11 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n406 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t18 535.019
R12 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n510 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t7 535.019
R13 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n491 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t10 535.019
R14 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n346 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t11 535.019
R15 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n328 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t9 535.019
R16 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n880 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t14 535.019
R17 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n862 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t8 535.019
R18 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n68 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n67 25.02
R19 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n258 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n257 24.875
R20 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n206 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n205 24.875
R21 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n154 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n153 24.875
R22 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n675 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n674 24.875
R23 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n781 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n780 24.875
R24 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n439 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n438 24.875
R25 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n386 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n385 24.875
R26 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n492 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n491 24.875
R27 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n728 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n727 24.875
R28 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n622 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n621 24.875
R29 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n906 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n905 24.733
R30 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n944 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n943 24.733
R31 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n982 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n981 24.733
R32 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n56 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n55 20.259
R33 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n697 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n696 20.259
R34 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n750 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n747 20.259
R35 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n966 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n965 20.259
R36 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n644 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n641 20.259
R37 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n928 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n927 20.259
R38 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1004 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1001 20.259
R39 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n803 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n802 20.259
R40 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n227 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n224 20.259
R41 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n461 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n460 20.259
R42 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n175 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n172 20.259
R43 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n408 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n407 20.259
R44 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n514 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n511 20.259
R45 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n279 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n278 20.259
R46 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n116 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n115 20.259
R47 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n98 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n95 20.259
R48 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n348 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n347 20.259
R49 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n330 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n329 20.259
R50 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n584 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n583 20.259
R51 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n566 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n563 20.259
R52 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n882 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n881 20.259
R53 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n864 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n863 20.259
R54 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n686 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n685 9.3
R55 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n689 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n688 9.3
R56 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n739 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n738 9.3
R57 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n742 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n741 9.3
R58 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n633 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n632 9.3
R59 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n636 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n635 9.3
R60 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n792 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n791 9.3
R61 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n795 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n794 9.3
R62 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n217 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n216 9.3
R63 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n220 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n219 9.3
R64 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n453 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n452 9.3
R65 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n450 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n449 9.3
R66 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n165 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n164 9.3
R67 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n168 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n167 9.3
R68 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n400 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n399 9.3
R69 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n397 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n396 9.3
R70 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n503 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n502 9.3
R71 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n506 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n505 9.3
R72 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n269 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n268 9.3
R73 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n272 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n271 9.3
R74 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n11 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n10 9.3
R75 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n42 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n41 9.3
R76 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n27 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n26 9.3
R77 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n13 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n12 9.3
R78 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n31 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n30 9.3
R79 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n17 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n16 9.3
R80 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n45 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n44 9.3
R81 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n3 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t2 9.162
R82 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n3 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t4 9.162
R83 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n684 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n683 9
R84 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n691 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n690 9
R85 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n737 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n736 9
R86 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n744 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n743 9
R87 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n960 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n959 9
R88 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n952 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n951 9
R89 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n631 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n630 9
R90 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n638 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n637 9
R91 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n922 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n921 9
R92 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n914 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n908 9
R93 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n998 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n997 9
R94 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n990 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n989 9
R95 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n790 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n789 9
R96 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n797 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n796 9
R97 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n215 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n214 9
R98 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n222 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n221 9
R99 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n448 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n447 9
R100 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n455 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n454 9
R101 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n163 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n162 9
R102 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n170 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n169 9
R103 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n395 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n394 9
R104 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n402 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n401 9
R105 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n501 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n500 9
R106 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n508 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n507 9
R107 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n267 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n266 9
R108 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n274 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n273 9
R109 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n122 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n121 9
R110 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n127 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n126 9
R111 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n356 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n355 9
R112 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n359 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n358 9
R113 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n590 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n589 9
R114 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n595 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n594 9
R115 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n888 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n887 9
R116 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n893 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n892 9
R117 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n51 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n50 9
R118 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n65 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n64 9
R119 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n20 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n19 9
R120 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n34 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n33 9
R121 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n47 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n46 9
R122 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n62 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n61 8.764
R123 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n688 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n687 8.764
R124 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n741 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n740 8.764
R125 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n948 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n947 8.764
R126 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n635 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n634 8.764
R127 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n911 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n910 8.764
R128 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n986 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n985 8.764
R129 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n794 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n793 8.764
R130 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n219 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n218 8.764
R131 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n452 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n451 8.764
R132 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n167 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n166 8.764
R133 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n399 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n398 8.764
R134 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n505 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n504 8.764
R135 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n271 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n270 8.764
R136 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n124 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n123 8.764
R137 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n352 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n351 8.764
R138 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n592 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n591 8.764
R139 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n890 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n889 8.764
R140 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n6 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n5 7.816
R141 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n55 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n54 6.885
R142 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n696 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n695 6.885
R143 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n747 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n746 6.885
R144 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n965 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n964 6.885
R145 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n641 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n640 6.885
R146 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n927 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n926 6.885
R147 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1001 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1000 6.885
R148 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n802 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n801 6.885
R149 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n224 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n223 6.885
R150 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n460 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n459 6.885
R151 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n172 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n171 6.885
R152 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n407 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n406 6.885
R153 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n511 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n510 6.885
R154 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n278 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n277 6.885
R155 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n115 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n114 6.885
R156 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n95 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n94 6.885
R157 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n347 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n346 6.885
R158 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n329 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n328 6.885
R159 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n583 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n582 6.885
R160 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n563 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n562 6.885
R161 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n881 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n880 6.885
R162 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n863 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n862 6.885
R163 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n79 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t0 4.829
R164 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n63 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n62 4.65
R165 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n949 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n948 4.65
R166 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n912 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n911 4.65
R167 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n987 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n986 4.65
R168 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n125 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n124 4.65
R169 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n357 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n352 4.65
R170 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n593 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n592 4.65
R171 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n891 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n890 4.65
R172 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1035 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n70 4.498
R173 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1037 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n60 4.491
R174 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1037 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n66 4.491
R175 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n698 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n697 4.452
R176 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n751 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n750 4.452
R177 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n645 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n644 4.452
R178 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n804 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n803 4.452
R179 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n462 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n461 4.452
R180 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n409 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n408 4.452
R181 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n515 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n514 4.452
R182 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n57 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n56 4.451
R183 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n228 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n227 4.451
R184 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n176 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n175 4.451
R185 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n280 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n279 4.451
R186 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n99 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n98 4.451
R187 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n331 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n330 4.451
R188 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n567 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n566 4.451
R189 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n865 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n864 4.451
R190 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n349 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n348 4.388
R191 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n117 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n116 4.387
R192 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n585 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n584 4.387
R193 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n883 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n882 4.387
R194 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n116 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n113 3.711
R195 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n348 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n345 3.711
R196 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n584 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n581 3.711
R197 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n882 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n879 3.711
R198 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n6 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n3 3.634
R199 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n56 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n53 3.335
R200 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n697 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n694 3.335
R201 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n750 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n749 3.335
R202 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n966 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n963 3.335
R203 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n644 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n643 3.335
R204 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n928 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n925 3.335
R205 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1004 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1003 3.335
R206 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n803 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n800 3.335
R207 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n227 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n226 3.335
R208 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n461 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n458 3.335
R209 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n175 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n174 3.335
R210 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n408 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n405 3.335
R211 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n514 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n513 3.335
R212 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n279 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n276 3.335
R213 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n98 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n97 3.335
R214 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n330 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n327 3.335
R215 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n566 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n565 3.335
R216 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n864 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n861 3.335
R217 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n967 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n966 3.272
R218 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n929 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n928 3.272
R219 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1005 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1004 3.272
R220 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n259 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n258 3.078
R221 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n207 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n206 3.078
R222 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n155 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n154 3.078
R223 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n676 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n675 3.077
R224 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n782 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n781 3.077
R225 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n440 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n439 3.077
R226 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n387 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n386 3.077
R227 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n493 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n492 3.077
R228 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n729 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n728 3.077
R229 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n623 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n622 3.077
R230 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n53 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n52 3.011
R231 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n694 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n693 3.011
R232 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n749 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n748 3.011
R233 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n963 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n962 3.011
R234 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n643 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n642 3.011
R235 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n925 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n924 3.011
R236 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1003 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1002 3.011
R237 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n800 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n799 3.011
R238 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n226 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n225 3.011
R239 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n458 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n457 3.011
R240 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n174 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n173 3.011
R241 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n405 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n404 3.011
R242 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n513 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n512 3.011
R243 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n276 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n275 3.011
R244 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n97 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n96 3.011
R245 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n327 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n326 3.011
R246 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n565 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n564 3.011
R247 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n861 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n860 3.011
R248 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n8 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n7 3.008
R249 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n103 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n102 3
R250 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n131 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n130 3
R251 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n363 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n362 3
R252 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n335 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n334 3
R253 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n599 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n598 3
R254 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n571 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n570 3
R255 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n869 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n868 3
R256 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n897 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n896 3
R257 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n21 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n20 3
R258 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n35 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n34 3
R259 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n48 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n47 3
R260 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n69 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n68 2.86
R261 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n113 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n112 2.635
R262 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n345 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n344 2.635
R263 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n581 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n580 2.635
R264 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n879 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n878 2.635
R265 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n907 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n906 2.566
R266 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n983 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n982 2.565
R267 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n945 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n944 2.565
R268 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n812 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n811 1.94
R269 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n759 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n758 1.94
R270 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n706 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n705 1.94
R271 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n653 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n652 1.94
R272 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n417 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n416 1.94
R273 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n470 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n469 1.94
R274 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n523 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n522 1.94
R275 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n288 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n287 1.94
R276 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n236 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n235 1.94
R277 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n184 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n183 1.94
R278 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n558 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n322 1.352
R279 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1032 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n856 1.284
R280 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n692 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/GATE 1.031
R281 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n745 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/GATE 1.031
R282 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n639 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE 1.031
R283 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n798 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/GATE 1.031
R284 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n509 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE 1.031
R285 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n456 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/GATE 1.031
R286 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n403 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/GATE 1.031
R287 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1033 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1032 0.971
R288 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1031 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1030 0.881
R289 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n855 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n854 0.881
R290 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n557 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n556 0.881
R291 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n322 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n321 0.881
R292 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n815 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n813 0.853
R293 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n820 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n772 0.853
R294 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n824 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n760 0.853
R295 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n829 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n719 0.853
R296 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n833 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n707 0.853
R297 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n838 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n666 0.853
R298 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n842 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n654 0.853
R299 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n847 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n613 0.853
R300 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n544 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n418 0.853
R301 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n535 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n471 0.853
R302 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n526 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n524 0.853
R303 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n291 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n289 0.853
R304 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n296 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n249 0.853
R305 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n300 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n237 0.853
R306 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n305 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n197 0.853
R307 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n309 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n185 0.853
R308 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n314 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n145 0.853
R309 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n549 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n377 0.853
R310 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n540 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n430 0.853
R311 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n531 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n483 0.853
R312 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n948 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n946 0.752
R313 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n911 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n909 0.752
R314 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n986 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n984 0.752
R315 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1021 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1020 0.477
R316 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n542 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n541 0.461
R317 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n307 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n306 0.461
R318 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1034 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1033 0.282
R319 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n856 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n558 0.223
R320 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1017 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1016 0.197
R321 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n5 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n4 0.189
R322 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n822 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n821 0.181
R323 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n831 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n830 0.181
R324 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n840 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n839 0.181
R325 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n533 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n532 0.181
R326 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n298 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n297 0.181
R327 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n16 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n15 0.178
R328 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n849 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n848 0.174
R329 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n551 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n550 0.174
R330 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n316 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n315 0.174
R331 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1025 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1024 0.173
R332 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n30 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n29 0.166
R333 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n322 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n133 0.151
R334 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n557 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n365 0.151
R335 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n855 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n601 0.151
R336 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1031 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n899 0.151
R337 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n90 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n89 0.1
R338 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1014 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1013 0.083
R339 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n558 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n557 0.076
R340 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n856 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n855 0.076
R341 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1032 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1031 0.076
R342 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n7 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n6 0.071
R343 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n934 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n933 0.069
R344 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n918 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n917 0.069
R345 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n972 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n971 0.069
R346 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n956 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n955 0.069
R347 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1010 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1009 0.069
R348 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n994 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n993 0.069
R349 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1021 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n937 0.066
R350 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1017 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n975 0.066
R351 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1023 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n919 0.065
R352 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1019 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n957 0.065
R353 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1015 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n995 0.065
R354 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n80 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n79 0.055
R355 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1005 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/GATE 0.05
R356 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n967 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/GATE 0.05
R357 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n929 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE 0.05
R358 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n567 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/GATE 0.048
R359 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n57 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/GATE 0.048
R360 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n99 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/GATE 0.048
R361 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n228 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/GATE 0.048
R362 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n176 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/GATE 0.048
R363 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n280 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE 0.048
R364 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n331 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/GATE 0.048
R365 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n865 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/GATE 0.048
R366 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1008 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1007 0.043
R367 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n970 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n969 0.043
R368 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n932 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n931 0.043
R369 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n107 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n106 0.043
R370 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n339 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n338 0.043
R371 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n575 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n574 0.043
R372 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n873 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n872 0.043
R373 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n657 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n656 0.041
R374 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n999 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n998 0.041
R375 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n710 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n709 0.041
R376 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n961 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n960 0.041
R377 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n940 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n939 0.041
R378 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n604 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n603 0.041
R379 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n923 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n922 0.041
R380 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n902 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n901 0.041
R381 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n978 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n977 0.041
R382 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n763 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n762 0.041
R383 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n188 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n187 0.041
R384 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n235 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n222 0.041
R385 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n423 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n422 0.041
R386 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n136 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n135 0.041
R387 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n183 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n170 0.041
R388 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n370 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n369 0.041
R389 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n476 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n475 0.041
R390 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n287 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n274 0.041
R391 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n240 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n239 0.041
R392 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n596 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n595 0.039
R393 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n59 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n58 0.039
R394 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n991 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n990 0.039
R395 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n953 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n952 0.039
R396 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n915 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n914 0.039
R397 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n128 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n127 0.039
R398 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n215 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n213 0.039
R399 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n231 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n230 0.039
R400 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n163 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n161 0.039
R401 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n179 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n178 0.039
R402 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n267 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n265 0.039
R403 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n283 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n282 0.039
R404 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n360 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n359 0.039
R405 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n894 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n893 0.039
R406 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n698 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n692 0.038
R407 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n751 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n745 0.038
R408 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n645 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n639 0.038
R409 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n804 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n798 0.038
R410 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n515 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n509 0.038
R411 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n462 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n456 0.038
R412 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n409 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n403 0.038
R413 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n42 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n40 0.038
R414 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n705 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n691 0.038
R415 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n706 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n673 0.038
R416 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n758 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n744 0.038
R417 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n759 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n726 0.038
R418 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n974 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n973 0.038
R419 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n653 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n620 0.038
R420 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n652 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n638 0.038
R421 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n936 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n935 0.038
R422 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1012 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1011 0.038
R423 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n811 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n797 0.038
R424 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n812 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n779 0.038
R425 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n522 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n508 0.038
R426 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n236 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n204 0.038
R427 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n469 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n455 0.038
R428 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n470 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n437 0.038
R429 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n184 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n152 0.038
R430 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n416 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n402 0.038
R431 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n417 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n384 0.038
R432 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n523 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n490 0.038
R433 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n288 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n256 0.038
R434 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n598 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n586 0.037
R435 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n70 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n69 0.037
R436 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n130 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n118 0.037
R437 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n362 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n350 0.037
R438 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n896 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n884 0.037
R439 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n684 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n682 0.036
R440 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n701 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n700 0.036
R441 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n669 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n668 0.036
R442 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n737 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n735 0.036
R443 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n754 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n753 0.036
R444 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n722 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n721 0.036
R445 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n941 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n940 0.036
R446 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n616 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n615 0.036
R447 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n631 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n629 0.036
R448 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n648 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n647 0.036
R449 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n903 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n902 0.036
R450 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n979 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n978 0.036
R451 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n790 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n788 0.036
R452 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n807 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n806 0.036
R453 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n775 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n774 0.036
R454 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n501 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n499 0.036
R455 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n518 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n517 0.036
R456 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n200 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n199 0.036
R457 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n448 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n446 0.036
R458 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n465 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n464 0.036
R459 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n433 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n432 0.036
R460 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n148 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n147 0.036
R461 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n395 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n393 0.036
R462 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n412 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n411 0.036
R463 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n380 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n379 0.036
R464 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n486 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n485 0.036
R465 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n252 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n251 0.036
R466 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/DRAIN vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1038 0.036
R467 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n993 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n983 0.035
R468 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n955 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n945 0.035
R469 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n917 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n907 0.035
R470 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1028 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1027 0.035
R471 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n852 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n851 0.035
R472 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n554 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n553 0.035
R473 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n319 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n318 0.035
R474 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n208 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n207 0.034
R475 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n156 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n155 0.034
R476 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n260 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n259 0.034
R477 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n132 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n131 0.034
R478 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n364 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n363 0.034
R479 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n600 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n599 0.034
R480 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n898 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n897 0.034
R481 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n17 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n14 0.033
R482 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n27 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n25 0.033
R483 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1023 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1022 0.033
R484 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1019 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1018 0.033
R485 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1015 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1014 0.033
R486 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n957 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n938 0.032
R487 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n919 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n900 0.032
R488 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n995 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n976 0.032
R489 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n588 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n587 0.032
R490 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n659 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n658 0.032
R491 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n712 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n711 0.032
R492 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n606 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n605 0.032
R493 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n765 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n764 0.032
R494 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n120 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n119 0.032
R495 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n190 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n189 0.032
R496 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n425 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n424 0.032
R497 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n138 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n137 0.032
R498 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n372 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n371 0.032
R499 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n478 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n477 0.032
R500 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n242 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n241 0.032
R501 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n354 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n353 0.032
R502 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n886 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n885 0.032
R503 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n677 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n676 0.031
R504 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n665 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n664 0.031
R505 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n730 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n729 0.031
R506 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n718 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n717 0.031
R507 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n612 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n611 0.031
R508 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n624 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n623 0.031
R509 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n783 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n782 0.031
R510 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n771 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n770 0.031
R511 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n494 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n493 0.031
R512 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n196 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n195 0.031
R513 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n441 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n440 0.031
R514 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n420 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n419 0.031
R515 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n144 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n143 0.031
R516 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n388 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n387 0.031
R517 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n367 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n366 0.031
R518 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n473 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n472 0.031
R519 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n248 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n247 0.031
R520 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n593 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n590 0.03
R521 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n569 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n568 0.03
R522 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n125 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n122 0.03
R523 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n101 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n100 0.03
R524 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n357 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n356 0.03
R525 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n333 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n332 0.03
R526 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n891 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n888 0.03
R527 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n867 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n866 0.03
R528 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n568 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n567 0.029
R529 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n58 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n57 0.029
R530 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n100 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n99 0.029
R531 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n332 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n331 0.029
R532 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n866 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n865 0.029
R533 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n109 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n108 0.029
R534 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n105 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n104 0.029
R535 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n341 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n340 0.029
R536 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n337 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n336 0.029
R537 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n577 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n576 0.029
R538 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n573 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n572 0.029
R539 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n875 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n874 0.029
R540 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n871 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n870 0.029
R541 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n13 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n11 0.028
R542 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n31 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n28 0.028
R543 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n595 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n593 0.028
R544 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n65 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n63 0.028
R545 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n127 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n125 0.028
R546 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n359 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n357 0.028
R547 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n893 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n891 0.028
R548 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1033 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n90 0.026
R549 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n0 0.026
R550 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n20 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n18 0.026
R551 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n222 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n220 0.026
R552 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n170 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n168 0.026
R553 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n274 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n272 0.026
R554 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n60 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n59 0.026
R555 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n7 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n2 0.024
R556 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n47 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n45 0.024
R557 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n691 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n689 0.024
R558 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n990 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n988 0.024
R559 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n744 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n742 0.024
R560 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n952 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n950 0.024
R561 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n638 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n636 0.024
R562 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n914 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n913 0.024
R563 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n797 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n795 0.024
R564 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n508 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n506 0.024
R565 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n217 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n215 0.024
R566 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n455 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n453 0.024
R567 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n165 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n163 0.024
R568 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n402 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n400 0.024
R569 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n269 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n267 0.024
R570 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n21 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n9 0.023
R571 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1006 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1005 0.022
R572 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n968 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n967 0.022
R573 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n930 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n929 0.022
R574 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n686 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n684 0.022
R575 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n739 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n737 0.022
R576 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n633 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n631 0.022
R577 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n792 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n790 0.022
R578 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n503 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n501 0.022
R579 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n450 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n448 0.022
R580 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n397 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n395 0.022
R581 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n229 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n228 0.021
R582 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n177 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n176 0.021
R583 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n281 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n280 0.021
R584 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n66 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n65 0.02
R585 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n60 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n51 0.019
R586 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n699 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n698 0.019
R587 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n752 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n751 0.019
R588 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n646 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n645 0.019
R589 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n805 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n804 0.019
R590 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n516 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n515 0.019
R591 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n463 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n462 0.019
R592 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n410 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n409 0.019
R593 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1024 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1023 0.017
R594 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1022 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1021 0.017
R595 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1020 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1019 0.017
R596 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1018 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1017 0.017
R597 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1016 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1015 0.017
R598 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n821 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n820 0.017
R599 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n830 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n829 0.017
R600 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n839 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n838 0.017
R601 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n848 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n847 0.017
R602 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n550 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n549 0.017
R603 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n541 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n540 0.017
R604 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n532 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n531 0.017
R605 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n297 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n296 0.017
R606 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n306 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n305 0.017
R607 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n315 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n314 0.017
R608 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n32 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n31 0.016
R609 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n818 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n817 0.016
R610 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n816 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n815 0.016
R611 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n827 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n826 0.016
R612 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n825 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n824 0.016
R613 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n836 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n835 0.016
R614 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n834 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n833 0.016
R615 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n845 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n844 0.016
R616 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n843 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n842 0.016
R617 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n547 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n546 0.016
R618 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n545 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n544 0.016
R619 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n538 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n537 0.016
R620 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n536 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n535 0.016
R621 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n529 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n528 0.016
R622 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n527 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n526 0.016
R623 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n294 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n293 0.016
R624 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n292 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n291 0.016
R625 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n303 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n302 0.016
R626 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n301 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n300 0.016
R627 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n312 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n311 0.016
R628 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n310 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n309 0.016
R629 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1029 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1028 0.015
R630 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n819 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n818 0.015
R631 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n828 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n827 0.015
R632 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n823 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n822 0.015
R633 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n837 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n836 0.015
R634 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n832 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n831 0.015
R635 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n846 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n845 0.015
R636 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n841 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n840 0.015
R637 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n853 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n852 0.015
R638 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n555 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n554 0.015
R639 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n548 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n547 0.015
R640 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n543 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n542 0.015
R641 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n539 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n538 0.015
R642 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n534 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n533 0.015
R643 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n530 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n529 0.015
R644 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n295 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n294 0.015
R645 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n304 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n303 0.015
R646 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n299 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n298 0.015
R647 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n313 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n312 0.015
R648 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n308 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n307 0.015
R649 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n320 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n319 0.015
R650 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n92 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n91 0.015
R651 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n324 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n323 0.015
R652 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n560 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n559 0.015
R653 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n858 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n857 0.015
R654 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1026 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1025 0.013
R655 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n850 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n849 0.013
R656 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n552 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n551 0.013
R657 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n317 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n316 0.013
R658 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n24 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n23 0.013
R659 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n38 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n37 0.013
R660 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n2 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1 0.012
R661 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n20 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n13 0.012
R662 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n34 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n27 0.012
R663 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n34 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n32 0.012
R664 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n93 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n92 0.012
R665 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n325 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n324 0.012
R666 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n561 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n560 0.012
R667 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n859 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n858 0.012
R668 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n79 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n78 0.011
R669 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n74 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n73 0.011
R670 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n992 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n991 0.011
R671 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n954 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n953 0.011
R672 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n916 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n915 0.011
R673 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n942 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n941 0.01
R674 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n904 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n903 0.01
R675 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n980 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n979 0.01
R676 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n108 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n107 0.01
R677 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n340 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n339 0.01
R678 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n576 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n575 0.01
R679 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n874 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n873 0.01
R680 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n35 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n24 0.01
R681 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n37 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n36 0.01
R682 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n39 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n38 0.01
R683 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n49 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n48 0.01
R684 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1038 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1037 0.01
R685 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n89 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n88 0.01
R686 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n43 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n42 0.009
R687 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n570 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n569 0.009
R688 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n102 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n101 0.009
R689 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n334 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n333 0.009
R690 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n868 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n867 0.009
R691 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n103 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n93 0.008
R692 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n335 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n325 0.008
R693 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n571 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n561 0.008
R694 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n869 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n859 0.008
R695 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n23 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n22 0.008
R696 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n73 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n72 0.008
R697 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n47 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n43 0.007
R698 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n213 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n212 0.007
R699 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n230 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n229 0.007
R700 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n161 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n160 0.007
R701 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n178 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n177 0.007
R702 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n265 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n264 0.007
R703 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n282 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n281 0.007
R704 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n682 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n681 0.006
R705 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n700 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n699 0.006
R706 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n660 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n659 0.006
R707 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n735 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n734 0.006
R708 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n753 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n752 0.006
R709 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n713 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n712 0.006
R710 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n607 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n606 0.006
R711 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n629 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n628 0.006
R712 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n647 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n646 0.006
R713 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n788 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n787 0.006
R714 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n806 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n805 0.006
R715 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n766 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n765 0.006
R716 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n499 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n498 0.006
R717 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n517 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n516 0.006
R718 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n191 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n190 0.006
R719 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n446 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n445 0.006
R720 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n464 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n463 0.006
R721 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n426 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n425 0.006
R722 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n139 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n138 0.006
R723 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n393 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n392 0.006
R724 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n411 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n410 0.006
R725 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n373 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n372 0.006
R726 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n479 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n478 0.006
R727 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n243 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n242 0.006
R728 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n110 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n109 0.006
R729 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n104 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n103 0.006
R730 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n342 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n341 0.006
R731 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n336 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n335 0.006
R732 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n578 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n577 0.006
R733 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n572 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n571 0.006
R734 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n876 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n875 0.006
R735 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n870 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n869 0.006
R736 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n9 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n8 0.006
R737 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n22 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n21 0.006
R738 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1035 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1034 0.005
R739 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1036 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1035 0.005
R740 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n586 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n585 0.005
R741 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n598 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n597 0.005
R742 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n590 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n588 0.005
R743 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n692 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/GATE 0.005
R744 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n745 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/GATE 0.005
R745 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n639 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE 0.005
R746 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n798 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/GATE 0.005
R747 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n118 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n117 0.005
R748 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n130 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n129 0.005
R749 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n122 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n120 0.005
R750 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n509 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE 0.005
R751 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n456 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/GATE 0.005
R752 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n403 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/GATE 0.005
R753 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n133 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n132 0.005
R754 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n131 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n111 0.005
R755 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n106 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n105 0.005
R756 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n350 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n349 0.005
R757 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n362 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n361 0.005
R758 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n356 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n354 0.005
R759 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n365 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n364 0.005
R760 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n363 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n343 0.005
R761 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n338 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n337 0.005
R762 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n601 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n600 0.005
R763 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n599 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n579 0.005
R764 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n574 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n573 0.005
R765 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n884 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n883 0.005
R766 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n896 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n895 0.005
R767 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n888 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n886 0.005
R768 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n899 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n898 0.005
R769 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n897 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n877 0.005
R770 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n872 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n871 0.005
R771 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n90 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n86 0.005
R772 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n72 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n71 0.005
R773 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n88 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n87 0.004
R774 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n76 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n75 0.004
R775 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1027 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1026 0.004
R776 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n851 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n850 0.004
R777 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n553 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n552 0.004
R778 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n318 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n317 0.004
R779 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n84 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n83 0.004
R780 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/DRAIN vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n49 0.004
R781 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n969 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n968 0.004
R782 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n931 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n930 0.004
R783 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1007 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1006 0.004
R784 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n689 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n686 0.003
R785 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n658 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n657 0.003
R786 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n656 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n655 0.003
R787 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n668 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n667 0.003
R788 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n988 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n987 0.003
R789 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n742 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n739 0.003
R790 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n711 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n710 0.003
R791 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n709 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n708 0.003
R792 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n721 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n720 0.003
R793 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n950 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n949 0.003
R794 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n605 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n604 0.003
R795 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n603 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n602 0.003
R796 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n615 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n614 0.003
R797 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n636 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n633 0.003
R798 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n913 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n912 0.003
R799 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1030 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1029 0.003
R800 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n795 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n792 0.003
R801 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n764 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n763 0.003
R802 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n762 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n761 0.003
R803 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n774 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n773 0.003
R804 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n854 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n853 0.003
R805 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n506 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n503 0.003
R806 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n189 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n188 0.003
R807 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n187 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n186 0.003
R808 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n199 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n198 0.003
R809 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n220 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n217 0.003
R810 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n453 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n450 0.003
R811 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n424 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n423 0.003
R812 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n422 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n421 0.003
R813 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n432 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n431 0.003
R814 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n137 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n136 0.003
R815 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n135 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n134 0.003
R816 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n147 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n146 0.003
R817 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n168 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n165 0.003
R818 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n400 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n397 0.003
R819 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n371 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n370 0.003
R820 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n369 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n368 0.003
R821 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n379 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n378 0.003
R822 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n556 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n555 0.003
R823 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n477 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n476 0.003
R824 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n475 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n474 0.003
R825 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n485 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n484 0.003
R826 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n272 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n269 0.003
R827 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n241 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n240 0.003
R828 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n239 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n238 0.003
R829 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n251 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n250 0.003
R830 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n321 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n320 0.003
R831 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n78 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n77 0.003
R832 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n18 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n17 0.002
R833 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n75 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n74 0.002
R834 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n77 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n76 0.002
R835 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n36 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n35 0.002
R836 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1037 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1036 0.002
R837 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n772 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n769 0.002
R838 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n813 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n778 0.002
R839 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n719 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n716 0.002
R840 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n760 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n725 0.002
R841 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n666 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n663 0.002
R842 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n707 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n672 0.002
R843 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n654 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n619 0.002
R844 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n613 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n610 0.002
R845 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n418 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n383 0.002
R846 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n471 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n436 0.002
R847 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n524 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n489 0.002
R848 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n249 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n246 0.002
R849 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n289 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n255 0.002
R850 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n237 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n203 0.002
R851 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n197 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n194 0.002
R852 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n185 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n151 0.002
R853 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n145 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n142 0.002
R854 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n937 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n936 0.002
R855 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n975 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n974 0.002
R856 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1013 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1012 0.002
R857 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n430 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n429 0.001
R858 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n377 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n376 0.001
R859 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n483 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n482 0.001
R860 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n937 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n934 0.001
R861 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n975 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n972 0.001
R862 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1013 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1010 0.001
R863 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n597 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n596 0.001
R864 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n678 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n677 0.001
R865 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n679 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n678 0.001
R866 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n680 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n679 0.001
R867 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n681 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n680 0.001
R868 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n705 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n704 0.001
R869 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n704 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n703 0.001
R870 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n703 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n702 0.001
R871 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n702 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n701 0.001
R872 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n663 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n662 0.001
R873 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n662 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n661 0.001
R874 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n661 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n660 0.001
R875 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n672 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n671 0.001
R876 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n671 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n670 0.001
R877 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n670 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n669 0.001
R878 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n993 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n992 0.001
R879 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1009 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n999 0.001
R880 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1009 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1008 0.001
R881 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n731 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n730 0.001
R882 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n732 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n731 0.001
R883 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n733 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n732 0.001
R884 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n734 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n733 0.001
R885 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n758 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n757 0.001
R886 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n757 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n756 0.001
R887 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n756 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n755 0.001
R888 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n755 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n754 0.001
R889 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n716 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n715 0.001
R890 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n715 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n714 0.001
R891 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n714 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n713 0.001
R892 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n725 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n724 0.001
R893 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n724 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n723 0.001
R894 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n723 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n722 0.001
R895 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n955 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n954 0.001
R896 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n971 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n961 0.001
R897 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n971 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n970 0.001
R898 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n956 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n942 0.001
R899 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n972 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n958 0.001
R900 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n610 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n609 0.001
R901 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n609 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n608 0.001
R902 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n608 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n607 0.001
R903 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n619 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n618 0.001
R904 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n618 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n617 0.001
R905 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n617 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n616 0.001
R906 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n625 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n624 0.001
R907 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n626 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n625 0.001
R908 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n627 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n626 0.001
R909 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n628 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n627 0.001
R910 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n652 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n651 0.001
R911 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n651 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n650 0.001
R912 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n650 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n649 0.001
R913 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n649 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n648 0.001
R914 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n917 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n916 0.001
R915 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n933 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n923 0.001
R916 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n933 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n932 0.001
R917 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n918 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n904 0.001
R918 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n934 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n920 0.001
R919 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n994 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n980 0.001
R920 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1010 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n996 0.001
R921 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n784 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n783 0.001
R922 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n785 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n784 0.001
R923 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n786 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n785 0.001
R924 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n787 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n786 0.001
R925 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n811 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n810 0.001
R926 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n810 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n809 0.001
R927 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n809 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n808 0.001
R928 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n808 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n807 0.001
R929 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n769 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n768 0.001
R930 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n768 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n767 0.001
R931 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n767 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n766 0.001
R932 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n778 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n777 0.001
R933 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n777 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n776 0.001
R934 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n776 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n775 0.001
R935 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n820 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n819 0.001
R936 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n817 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n816 0.001
R937 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n815 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n814 0.001
R938 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n829 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n828 0.001
R939 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n826 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n825 0.001
R940 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n824 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n823 0.001
R941 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n838 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n837 0.001
R942 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n835 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n834 0.001
R943 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n833 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n832 0.001
R944 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n847 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n846 0.001
R945 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n844 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n843 0.001
R946 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n842 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n841 0.001
R947 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n129 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n128 0.001
R948 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n495 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n494 0.001
R949 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n496 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n495 0.001
R950 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n497 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n496 0.001
R951 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n498 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n497 0.001
R952 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n522 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n521 0.001
R953 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n521 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n520 0.001
R954 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n520 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n519 0.001
R955 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n519 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n518 0.001
R956 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n194 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n193 0.001
R957 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n193 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n192 0.001
R958 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n192 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n191 0.001
R959 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n203 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n202 0.001
R960 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n202 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n201 0.001
R961 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n201 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n200 0.001
R962 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n209 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n208 0.001
R963 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n210 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n209 0.001
R964 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n211 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n210 0.001
R965 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n212 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n211 0.001
R966 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n235 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n234 0.001
R967 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n234 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n233 0.001
R968 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n233 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n232 0.001
R969 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n232 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n231 0.001
R970 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n442 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n441 0.001
R971 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n443 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n442 0.001
R972 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n444 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n443 0.001
R973 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n445 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n444 0.001
R974 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n469 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n468 0.001
R975 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n468 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n467 0.001
R976 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n467 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n466 0.001
R977 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n466 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n465 0.001
R978 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n429 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n428 0.001
R979 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n428 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n427 0.001
R980 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n427 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n426 0.001
R981 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n436 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n435 0.001
R982 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n435 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n434 0.001
R983 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n434 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n433 0.001
R984 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n142 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n141 0.001
R985 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n141 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n140 0.001
R986 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n140 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n139 0.001
R987 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n151 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n150 0.001
R988 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n150 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n149 0.001
R989 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n149 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n148 0.001
R990 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n157 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n156 0.001
R991 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n158 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n157 0.001
R992 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n159 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n158 0.001
R993 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n160 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n159 0.001
R994 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n183 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n182 0.001
R995 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n182 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n181 0.001
R996 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n181 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n180 0.001
R997 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n180 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n179 0.001
R998 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n389 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n388 0.001
R999 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n390 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n389 0.001
R1000 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n391 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n390 0.001
R1001 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n392 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n391 0.001
R1002 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n416 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n415 0.001
R1003 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n415 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n414 0.001
R1004 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n414 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n413 0.001
R1005 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n413 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n412 0.001
R1006 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n376 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n375 0.001
R1007 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n375 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n374 0.001
R1008 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n374 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n373 0.001
R1009 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n383 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n382 0.001
R1010 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n382 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n381 0.001
R1011 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n381 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n380 0.001
R1012 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n549 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n548 0.001
R1013 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n546 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n545 0.001
R1014 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n544 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n543 0.001
R1015 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n540 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n539 0.001
R1016 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n537 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n536 0.001
R1017 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n535 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n534 0.001
R1018 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n531 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n530 0.001
R1019 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n528 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n527 0.001
R1020 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n526 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n525 0.001
R1021 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n482 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n481 0.001
R1022 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n481 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n480 0.001
R1023 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n480 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n479 0.001
R1024 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n489 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n488 0.001
R1025 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n488 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n487 0.001
R1026 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n487 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n486 0.001
R1027 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n261 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n260 0.001
R1028 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n262 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n261 0.001
R1029 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n263 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n262 0.001
R1030 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n264 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n263 0.001
R1031 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n287 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n286 0.001
R1032 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n286 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n285 0.001
R1033 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n285 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n284 0.001
R1034 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n284 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n283 0.001
R1035 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n246 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n245 0.001
R1036 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n245 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n244 0.001
R1037 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n244 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n243 0.001
R1038 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n255 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n254 0.001
R1039 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n254 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n253 0.001
R1040 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n253 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n252 0.001
R1041 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n296 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n295 0.001
R1042 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n293 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n292 0.001
R1043 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n291 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n290 0.001
R1044 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n305 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n304 0.001
R1045 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n302 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n301 0.001
R1046 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n300 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n299 0.001
R1047 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n314 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n313 0.001
R1048 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n311 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n310 0.001
R1049 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n309 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n308 0.001
R1050 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n111 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n110 0.001
R1051 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n361 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n360 0.001
R1052 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n343 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n342 0.001
R1053 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n579 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n578 0.001
R1054 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n895 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n894 0.001
R1055 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n877 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n876 0.001
R1056 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n86 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n85 0.001
R1057 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n85 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n84 0.001
R1058 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n83 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n82 0.001
R1059 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n82 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n81 0.001
R1060 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n81 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n80 0.001
R1061 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n48 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n39 0.001
R1062 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n813 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n812 0.001
R1063 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n772 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n771 0.001
R1064 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n719 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n718 0.001
R1065 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n760 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n759 0.001
R1066 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n707 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n706 0.001
R1067 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n666 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n665 0.001
R1068 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n613 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n612 0.001
R1069 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n654 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n653 0.001
R1070 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n418 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n417 0.001
R1071 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n471 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n470 0.001
R1072 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n524 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n523 0.001
R1073 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n289 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n288 0.001
R1074 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n249 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n248 0.001
R1075 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n197 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n196 0.001
R1076 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n237 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n236 0.001
R1077 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n145 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n144 0.001
R1078 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n185 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n184 0.001
R1079 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n377 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n367 0.001
R1080 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n430 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n420 0.001
R1081 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n483 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n473 0.001
R1082 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n919 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n918 0.001
R1083 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n957 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n956 0.001
R1084 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n995 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n994 0.001
R1085 VDD.n3076 VDD.t37 535.019
R1086 VDD.n2858 VDD.t9 535.019
R1087 VDD.n1859 VDD.t17 535.019
R1088 VDD.n1847 VDD.t12 535.019
R1089 VDD.n2417 VDD.t5 535.019
R1090 VDD.n3431 VDD.t0 535.019
R1091 VDD.n1614 VDD.t34 535.019
R1092 VDD.n1621 VDD.t21 535.019
R1093 VDD.n1907 VDD.t25 535.019
R1094 VDD.n3620 VDD.t30 535.019
R1095 VDD.n1878 VDD.n1876 82.758
R1096 VDD.n1506 VDD.n1505 82.758
R1097 VDD.n1896 VDD.n1894 70.344
R1098 VDD.n660 VDD.n659 70.344
R1099 VDD.n2204 VDD.n2202 57.931
R1100 VDD.n2373 VDD.n2372 57.931
R1101 VDD.n3612 VDD.n3610 45.517
R1102 VDD.n2391 VDD.n2390 45.517
R1103 VDD.n3134 VDD.n3133 33.103
R1104 VDD.n3247 VDD.n3246 33.103
R1105 VDD.n731 VDD.n730 33.103
R1106 VDD.n2303 VDD.n2302 33.103
R1107 VDD.n2066 VDD.n2065 33.103
R1108 VDD.n1966 VDD.n1965 33.103
R1109 VDD.n324 VDD.n323 33.103
R1110 VDD.n3509 VDD.n3508 33.103
R1111 VDD.n373 VDD.n372 33.103
R1112 VDD.n377 VDD.n376 33.103
R1113 VDD.n597 VDD.n596 33.103
R1114 VDD.n606 VDD.n605 33.103
R1115 VDD.n1155 VDD.n1154 33.103
R1116 VDD.n1563 VDD.n1562 33.103
R1117 VDD.n1555 VDD.n1554 33.103
R1118 VDD.n3588 VDD.n3586 33.103
R1119 VDD.n3048 VDD.n3047 33.103
R1120 VDD.n3361 VDD.n3360 33.103
R1121 VDD.n3370 VDD.n3369 33.103
R1122 VDD.n2409 VDD.n2408 33.103
R1123 VDD.n1784 VDD.n1783 33.103
R1124 VDD.n1407 VDD.n1406 33.103
R1125 VDD.n376 VDD.n375 31.001
R1126 VDD.n605 VDD.n604 31.001
R1127 VDD.n1554 VDD.n1553 31.001
R1128 VDD.n3369 VDD.n3368 31.001
R1129 VDD.n3067 VDD.n3066 30.117
R1130 VDD.n3423 VDD.n3421 30.117
R1131 VDD.n3122 VDD.n3121 28.965
R1132 VDD.n3259 VDD.n3258 28.965
R1133 VDD.n674 VDD.n673 28.965
R1134 VDD.n2291 VDD.n2290 28.965
R1135 VDD.n2054 VDD.n2053 28.965
R1136 VDD.n1978 VDD.n1977 28.965
R1137 VDD.n268 VDD.n267 28.965
R1138 VDD.n3521 VDD.n3520 28.965
R1139 VDD.n1095 VDD.n1094 28.965
R1140 VDD.n2991 VDD.n2990 28.965
R1141 VDD.n1796 VDD.n1795 28.965
R1142 VDD.n1395 VDD.n1394 28.965
R1143 VDD.n2231 VDD.n2226 26.352
R1144 VDD.n3583 VDD.n3582 26.352
R1145 VDD.n433 VDD.n428 26.352
R1146 VDD.n1173 VDD.n1168 26.352
R1147 VDD.n3061 VDD.n2979 26.352
R1148 VDD.n3110 VDD.n3109 24.827
R1149 VDD.n3271 VDD.n3270 24.827
R1150 VDD.n740 VDD.n739 24.827
R1151 VDD.n2279 VDD.n2278 24.827
R1152 VDD.n2042 VDD.n2041 24.827
R1153 VDD.n1990 VDD.n1989 24.827
R1154 VDD.n333 VDD.n332 24.827
R1155 VDD.n3533 VDD.n3532 24.827
R1156 VDD.n354 VDD.n353 24.827
R1157 VDD.n396 VDD.n395 24.827
R1158 VDD.n572 VDD.n571 24.827
R1159 VDD.n631 VDD.n630 24.827
R1160 VDD.n1164 VDD.n1163 24.827
R1161 VDD.n1587 VDD.n1586 24.827
R1162 VDD.n1530 VDD.n1529 24.827
R1163 VDD.n3057 VDD.n3056 24.827
R1164 VDD.n3336 VDD.n3335 24.827
R1165 VDD.n3395 VDD.n3394 24.827
R1166 VDD.n1808 VDD.n1807 24.827
R1167 VDD.n1383 VDD.n1382 24.827
R1168 VDD.n3077 VDD.n3076 24.127
R1169 VDD.n2859 VDD.n2858 24.127
R1170 VDD.n2682 VDD.n2681 24.127
R1171 VDD.n2947 VDD.n2946 24.127
R1172 VDD.n1723 VDD.n1722 24.127
R1173 VDD.n1268 VDD.n1267 24.127
R1174 VDD.n1848 VDD.n1847 24.127
R1175 VDD.n1860 VDD.n1859 24.127
R1176 VDD.n3432 VDD.n3431 24.127
R1177 VDD.n2418 VDD.n2417 24.127
R1178 VDD.n3301 VDD.n3300 24.127
R1179 VDD.n3308 VDD.n3307 24.127
R1180 VDD.n1473 VDD.n1472 24.127
R1181 VDD.n1483 VDD.n1482 24.127
R1182 VDD.n1622 VDD.n1621 24.127
R1183 VDD.n1615 VDD.n1614 24.127
R1184 VDD.n1908 VDD.n1907 24.127
R1185 VDD.n3621 VDD.n3620 24.127
R1186 VDD.n2122 VDD.n2121 24.127
R1187 VDD.n542 VDD.n541 24.127
R1188 VDD.n3098 VDD.n3097 20.689
R1189 VDD.n3283 VDD.n3282 20.689
R1190 VDD.n3202 VDD.n3201 20.689
R1191 VDD.n665 VDD.n664 20.689
R1192 VDD.n2267 VDD.n2266 20.689
R1193 VDD.n2347 VDD.n2346 20.689
R1194 VDD.n2030 VDD.n2029 20.689
R1195 VDD.n2002 VDD.n2001 20.689
R1196 VDD.n1923 VDD.n1922 20.689
R1197 VDD.n259 VDD.n258 20.689
R1198 VDD.n3545 VDD.n3544 20.689
R1199 VDD.n3465 VDD.n3464 20.689
R1200 VDD.n1086 VDD.n1085 20.689
R1201 VDD.n2676 VDD.n2674 20.689
R1202 VDD.n2982 VDD.n2981 20.689
R1203 VDD.n3441 VDD.n3440 20.689
R1204 VDD.n1371 VDD.n1370 20.689
R1205 VDD.n1841 VDD.t13 19.133
R1206 VDD.n1889 VDD.t59 19.133
R1207 VDD.n1865 VDD.t18 16.263
R1208 VDD.n1881 VDD.t50 16.263
R1209 VDD.n2212 VDD.t43 16.263
R1210 VDD.n3143 VDD.n3142 15.193
R1211 VDD.n3240 VDD.n3239 15.193
R1212 VDD.n717 VDD.n716 15.193
R1213 VDD.n2312 VDD.n2311 15.193
R1214 VDD.n2075 VDD.n2074 15.193
R1215 VDD.n1959 VDD.n1958 15.193
R1216 VDD.n310 VDD.n309 15.193
R1217 VDD.n3502 VDD.n3501 15.193
R1218 VDD.n309 VDD.n308 15.193
R1219 VDD.n3501 VDD.n3500 15.193
R1220 VDD.n2074 VDD.n2073 15.193
R1221 VDD.n1958 VDD.n1957 15.193
R1222 VDD.n716 VDD.n715 15.193
R1223 VDD.n2311 VDD.n2310 15.193
R1224 VDD.n1141 VDD.n1140 15.193
R1225 VDD.n1140 VDD.n1139 15.193
R1226 VDD.n3034 VDD.n3033 15.193
R1227 VDD.n1777 VDD.n1776 15.193
R1228 VDD.n1416 VDD.n1415 15.193
R1229 VDD.n1415 VDD.n1414 15.193
R1230 VDD.n1776 VDD.n1775 15.193
R1231 VDD.n3142 VDD.n3141 15.193
R1232 VDD.n3239 VDD.n3238 15.193
R1233 VDD.n3033 VDD.n3032 15.193
R1234 VDD.n1879 VDD.n1875 15.058
R1235 VDD.n1507 VDD.n1504 15.058
R1236 VDD.n3180 VDD.n3179 14.482
R1237 VDD.n702 VDD.n696 14.482
R1238 VDD.n2348 VDD.n2347 14.482
R1239 VDD.n2112 VDD.n2111 14.482
R1240 VDD.n1924 VDD.n1923 14.482
R1241 VDD.n295 VDD.n289 14.482
R1242 VDD.n3466 VDD.n3465 14.482
R1243 VDD.n346 VDD.n345 14.482
R1244 VDD.n412 VDD.n406 14.482
R1245 VDD.n562 VDD.n561 14.482
R1246 VDD.n645 VDD.n644 14.482
R1247 VDD.n1114 VDD.n1108 14.482
R1248 VDD.n1601 VDD.n1600 14.482
R1249 VDD.n1520 VDD.n1519 14.482
R1250 VDD.n3010 VDD.n3004 14.482
R1251 VDD.n3326 VDD.n3325 14.482
R1252 VDD.n3409 VDD.n3408 14.482
R1253 VDD.n1822 VDD.n1821 14.482
R1254 VDD.n1742 VDD.n1741 14.482
R1255 VDD.n1453 VDD.n1452 14.482
R1256 VDD.n3155 VDD.n3154 13.432
R1257 VDD.n3228 VDD.n3227 13.432
R1258 VDD.n678 VDD.n677 13.432
R1259 VDD.n2324 VDD.n2323 13.432
R1260 VDD.n2087 VDD.n2086 13.432
R1261 VDD.n1947 VDD.n1946 13.432
R1262 VDD.n272 VDD.n271 13.432
R1263 VDD.n3490 VDD.n3489 13.432
R1264 VDD.n271 VDD.n270 13.432
R1265 VDD.n3489 VDD.n3488 13.432
R1266 VDD.n2086 VDD.n2085 13.432
R1267 VDD.n1946 VDD.n1945 13.432
R1268 VDD.n677 VDD.n676 13.432
R1269 VDD.n2323 VDD.n2322 13.432
R1270 VDD.n358 VDD.n357 13.432
R1271 VDD.n386 VDD.n385 13.432
R1272 VDD.n585 VDD.n584 13.432
R1273 VDD.n618 VDD.n617 13.432
R1274 VDD.n619 VDD.n618 13.432
R1275 VDD.n387 VDD.n386 13.432
R1276 VDD.n357 VDD.n356 13.432
R1277 VDD.n584 VDD.n583 13.432
R1278 VDD.n1099 VDD.n1098 13.432
R1279 VDD.n1576 VDD.n1575 13.432
R1280 VDD.n1542 VDD.n1541 13.432
R1281 VDD.n1098 VDD.n1097 13.432
R1282 VDD.n1543 VDD.n1542 13.432
R1283 VDD.n1575 VDD.n1574 13.432
R1284 VDD.n2995 VDD.n2994 13.432
R1285 VDD.n3349 VDD.n3348 13.432
R1286 VDD.n3382 VDD.n3381 13.432
R1287 VDD.n1765 VDD.n1764 13.432
R1288 VDD.n1428 VDD.n1427 13.432
R1289 VDD.n1427 VDD.n1426 13.432
R1290 VDD.n1764 VDD.n1763 13.432
R1291 VDD.n3154 VDD.n3153 13.432
R1292 VDD.n3227 VDD.n3226 13.432
R1293 VDD.n2994 VDD.n2993 13.432
R1294 VDD.n3383 VDD.n3382 13.432
R1295 VDD.n3348 VDD.n3347 13.432
R1296 VDD.n2216 VDD.t53 13.393
R1297 VDD.n3623 VDD.t31 13.393
R1298 VDD.n3099 VDD.n3098 12.833
R1299 VDD.n3284 VDD.n3283 12.833
R1300 VDD.n3203 VDD.n3202 12.833
R1301 VDD.n666 VDD.n665 12.833
R1302 VDD.n2268 VDD.n2267 12.833
R1303 VDD.n2031 VDD.n2030 12.833
R1304 VDD.n2003 VDD.n2002 12.833
R1305 VDD.n260 VDD.n259 12.833
R1306 VDD.n3546 VDD.n3545 12.833
R1307 VDD.n1087 VDD.n1086 12.833
R1308 VDD.n2983 VDD.n2982 12.833
R1309 VDD.n1372 VDD.n1371 12.833
R1310 VDD.n1897 VDD.n1893 12.8
R1311 VDD.n661 VDD.n658 12.8
R1312 VDD.n3167 VDD.n3166 11.633
R1313 VDD.n3215 VDD.n3214 11.633
R1314 VDD.n708 VDD.n707 11.633
R1315 VDD.n2336 VDD.n2335 11.633
R1316 VDD.n2099 VDD.n2098 11.633
R1317 VDD.n1935 VDD.n1934 11.633
R1318 VDD.n301 VDD.n300 11.633
R1319 VDD.n3477 VDD.n3476 11.633
R1320 VDD.n300 VDD.n299 11.633
R1321 VDD.n3476 VDD.n3475 11.633
R1322 VDD.n2098 VDD.n2097 11.633
R1323 VDD.n1934 VDD.n1933 11.633
R1324 VDD.n707 VDD.n706 11.633
R1325 VDD.n2335 VDD.n2334 11.633
R1326 VDD.n1132 VDD.n1131 11.633
R1327 VDD.n1131 VDD.n1130 11.633
R1328 VDD.n3025 VDD.n3024 11.633
R1329 VDD.n1753 VDD.n1752 11.633
R1330 VDD.n1440 VDD.n1439 11.633
R1331 VDD.n1439 VDD.n1438 11.633
R1332 VDD.n1752 VDD.n1751 11.633
R1333 VDD.n3166 VDD.n3165 11.633
R1334 VDD.n3214 VDD.n3213 11.633
R1335 VDD.n3024 VDD.n3023 11.633
R1336 VDD.n2206 VDD.n2205 10.541
R1337 VDD.n2374 VDD.n2371 10.541
R1338 VDD.n1909 VDD.t26 10.523
R1339 VDD.n3596 VDD.t41 10.523
R1340 VDD.n3168 VDD.n3167 10.344
R1341 VDD.n3217 VDD.n3215 10.344
R1342 VDD.n714 VDD.n708 10.344
R1343 VDD.n2337 VDD.n2336 10.344
R1344 VDD.n2100 VDD.n2099 10.344
R1345 VDD.n1936 VDD.n1935 10.344
R1346 VDD.n307 VDD.n301 10.344
R1347 VDD.n3479 VDD.n3477 10.344
R1348 VDD.n1138 VDD.n1132 10.344
R1349 VDD.n3031 VDD.n3025 10.344
R1350 VDD.n1754 VDD.n1753 10.344
R1351 VDD.n1441 VDD.n1440 10.344
R1352 VDD.n3179 VDD.n3178 9.797
R1353 VDD.n696 VDD.n695 9.797
R1354 VDD.n2111 VDD.n2110 9.797
R1355 VDD.n289 VDD.n288 9.797
R1356 VDD.n288 VDD.n287 9.797
R1357 VDD.n2110 VDD.n2109 9.797
R1358 VDD.n695 VDD.n694 9.797
R1359 VDD.n345 VDD.n344 9.797
R1360 VDD.n405 VDD.n404 9.797
R1361 VDD.n561 VDD.n560 9.797
R1362 VDD.n643 VDD.n642 9.797
R1363 VDD.n644 VDD.n643 9.797
R1364 VDD.n406 VDD.n405 9.797
R1365 VDD.n344 VDD.n343 9.797
R1366 VDD.n560 VDD.n559 9.797
R1367 VDD.n1108 VDD.n1107 9.797
R1368 VDD.n1600 VDD.n1599 9.797
R1369 VDD.n1518 VDD.n1517 9.797
R1370 VDD.n1107 VDD.n1106 9.797
R1371 VDD.n1599 VDD.n1598 9.797
R1372 VDD.n1519 VDD.n1518 9.797
R1373 VDD.n3004 VDD.n3003 9.797
R1374 VDD.n3325 VDD.n3324 9.797
R1375 VDD.n3407 VDD.n3406 9.797
R1376 VDD.n1820 VDD.n1819 9.797
R1377 VDD.n1741 VDD.n1740 9.797
R1378 VDD.n1452 VDD.n1451 9.797
R1379 VDD.n1451 VDD.n1450 9.797
R1380 VDD.n1740 VDD.n1739 9.797
R1381 VDD.n1821 VDD.n1820 9.797
R1382 VDD.n3178 VDD.n3177 9.797
R1383 VDD.n3003 VDD.n3002 9.797
R1384 VDD.n3408 VDD.n3407 9.797
R1385 VDD.n3324 VDD.n3323 9.797
R1386 VDD.n2812 VDD.n2811 9.411
R1387 VDD.n1238 VDD.n1237 9.411
R1388 VDD.n802 VDD.n801 9.411
R1389 VDD.n2545 VDD.n2544 9.411
R1390 VDD.n2605 VDD.n2604 9.411
R1391 VDD.n2453 VDD.n2452 9.411
R1392 VDD.n984 VDD.n983 9.411
R1393 VDD.n1335 VDD.n1334 9.411
R1394 VDD.n1045 VDD.n1044 9.411
R1395 VDD.n217 VDD.n216 9.411
R1396 VDD.n2156 VDD.n2155 9.411
R1397 VDD.n512 VDD.n511 9.411
R1398 VDD.n1693 VDD.n1692 9.411
R1399 VDD.n2716 VDD.n2715 9.411
R1400 VDD.n2917 VDD.n2916 9.411
R1401 VDD.n3111 VDD.n3110 9.352
R1402 VDD.n3272 VDD.n3271 9.352
R1403 VDD.n741 VDD.n740 9.352
R1404 VDD.n2280 VDD.n2279 9.352
R1405 VDD.n2043 VDD.n2042 9.352
R1406 VDD.n1991 VDD.n1990 9.352
R1407 VDD.n334 VDD.n333 9.352
R1408 VDD.n3534 VDD.n3533 9.352
R1409 VDD.n403 VDD.n396 9.352
R1410 VDD.n632 VDD.n631 9.352
R1411 VDD.n573 VDD.n572 9.352
R1412 VDD.n355 VDD.n354 9.352
R1413 VDD.n1165 VDD.n1164 9.352
R1414 VDD.n1531 VDD.n1530 9.352
R1415 VDD.n1588 VDD.n1587 9.352
R1416 VDD.n3058 VDD.n3057 9.352
R1417 VDD.n3396 VDD.n3395 9.352
R1418 VDD.n1809 VDD.n1808 9.352
R1419 VDD.n1384 VDD.n1383 9.352
R1420 VDD.n3337 VDD.n3336 9.352
R1421 VDD.n2789 VDD.n2788 9.3
R1422 VDD.n2777 VDD.n2776 9.3
R1423 VDD.n2836 VDD.n2835 9.3
R1424 VDD.n2831 VDD.n2830 9.3
R1425 VDD.n2824 VDD.n2823 9.3
R1426 VDD.n2817 VDD.n2816 9.3
R1427 VDD.n2834 VDD.n2833 9.3
R1428 VDD.n2829 VDD.n2828 9.3
R1429 VDD.n2827 VDD.n2826 9.3
R1430 VDD.n2822 VDD.n2821 9.3
R1431 VDD.n2820 VDD.n2819 9.3
R1432 VDD.n2815 VDD.n2814 9.3
R1433 VDD.n2782 VDD.n2781 9.3
R1434 VDD.n2787 VDD.n2786 9.3
R1435 VDD.n2794 VDD.n2793 9.3
R1436 VDD.n2810 VDD.n2809 9.3
R1437 VDD.n2813 VDD.n2812 9.3
R1438 VDD.n2838 VDD.n2837 9.3
R1439 VDD.n2842 VDD.n2841 9.3
R1440 VDD.n2768 VDD.n2767 9.3
R1441 VDD.n2764 VDD.n2763 9.3
R1442 VDD.n2773 VDD.n2772 9.3
R1443 VDD.n779 VDD.n778 9.3
R1444 VDD.n767 VDD.n766 9.3
R1445 VDD.n826 VDD.n825 9.3
R1446 VDD.n821 VDD.n820 9.3
R1447 VDD.n814 VDD.n813 9.3
R1448 VDD.n807 VDD.n806 9.3
R1449 VDD.n824 VDD.n823 9.3
R1450 VDD.n819 VDD.n818 9.3
R1451 VDD.n817 VDD.n816 9.3
R1452 VDD.n812 VDD.n811 9.3
R1453 VDD.n810 VDD.n809 9.3
R1454 VDD.n805 VDD.n804 9.3
R1455 VDD.n772 VDD.n771 9.3
R1456 VDD.n777 VDD.n776 9.3
R1457 VDD.n784 VDD.n783 9.3
R1458 VDD.n800 VDD.n799 9.3
R1459 VDD.n803 VDD.n802 9.3
R1460 VDD.n828 VDD.n827 9.3
R1461 VDD.n831 VDD.n830 9.3
R1462 VDD.n758 VDD.n757 9.3
R1463 VDD.n754 VDD.n753 9.3
R1464 VDD.n763 VDD.n762 9.3
R1465 VDD.n2571 VDD.n2570 9.3
R1466 VDD.n2564 VDD.n2563 9.3
R1467 VDD.n2557 VDD.n2556 9.3
R1468 VDD.n2550 VDD.n2549 9.3
R1469 VDD.n2546 VDD.n2545 9.3
R1470 VDD.n2526 VDD.n2525 9.3
R1471 VDD.n2543 VDD.n2542 9.3
R1472 VDD.n2548 VDD.n2547 9.3
R1473 VDD.n2553 VDD.n2552 9.3
R1474 VDD.n2555 VDD.n2554 9.3
R1475 VDD.n2560 VDD.n2559 9.3
R1476 VDD.n2562 VDD.n2561 9.3
R1477 VDD.n2567 VDD.n2566 9.3
R1478 VDD.n2569 VDD.n2568 9.3
R1479 VDD.n2574 VDD.n2573 9.3
R1480 VDD.n2510 VDD.n2509 9.3
R1481 VDD.n2506 VDD.n2505 9.3
R1482 VDD.n2501 VDD.n2500 9.3
R1483 VDD.n2497 VDD.n2496 9.3
R1484 VDD.n2515 VDD.n2514 9.3
R1485 VDD.n2519 VDD.n2518 9.3
R1486 VDD.n2521 VDD.n2520 9.3
R1487 VDD.n2454 VDD.n2453 9.3
R1488 VDD.n2460 VDD.n2459 9.3
R1489 VDD.n2484 VDD.n2483 9.3
R1490 VDD.n2480 VDD.n2479 9.3
R1491 VDD.n2475 VDD.n2474 9.3
R1492 VDD.n2471 VDD.n2470 9.3
R1493 VDD.n2466 VDD.n2465 9.3
R1494 VDD.n2464 VDD.n2463 9.3
R1495 VDD.n2490 VDD.n2489 9.3
R1496 VDD.n2430 VDD.n2429 9.3
R1497 VDD.n2435 VDD.n2434 9.3
R1498 VDD.n2442 VDD.n2441 9.3
R1499 VDD.n2451 VDD.n2450 9.3
R1500 VDD.n2433 VDD.n2432 9.3
R1501 VDD.n2437 VDD.n2436 9.3
R1502 VDD.n2440 VDD.n2439 9.3
R1503 VDD.n2444 VDD.n2443 9.3
R1504 VDD.n2447 VDD.n2446 9.3
R1505 VDD.n2449 VDD.n2448 9.3
R1506 VDD.n2428 VDD.n2427 9.3
R1507 VDD.n2426 VDD.n2425 9.3
R1508 VDD.n2456 VDD.n2455 9.3
R1509 VDD.n2606 VDD.n2605 9.3
R1510 VDD.n2612 VDD.n2611 9.3
R1511 VDD.n2616 VDD.n2615 9.3
R1512 VDD.n2618 VDD.n2617 9.3
R1513 VDD.n2623 VDD.n2622 9.3
R1514 VDD.n2627 VDD.n2626 9.3
R1515 VDD.n2632 VDD.n2631 9.3
R1516 VDD.n2636 VDD.n2635 9.3
R1517 VDD.n2656 VDD.n2655 9.3
R1518 VDD.n2582 VDD.n2581 9.3
R1519 VDD.n2587 VDD.n2586 9.3
R1520 VDD.n2594 VDD.n2593 9.3
R1521 VDD.n2603 VDD.n2602 9.3
R1522 VDD.n2585 VDD.n2584 9.3
R1523 VDD.n2589 VDD.n2588 9.3
R1524 VDD.n2592 VDD.n2591 9.3
R1525 VDD.n2596 VDD.n2595 9.3
R1526 VDD.n2599 VDD.n2598 9.3
R1527 VDD.n2601 VDD.n2600 9.3
R1528 VDD.n2580 VDD.n2579 9.3
R1529 VDD.n2416 VDD.n2415 9.3
R1530 VDD.n2608 VDD.n2607 9.3
R1531 VDD.n3303 VDD.n3302 9.3
R1532 VDD.n3299 VDD.n3298 9.3
R1533 VDD.n3310 VDD.n3309 9.3
R1534 VDD.n3312 VDD.n3311 9.3
R1535 VDD.n961 VDD.n960 9.3
R1536 VDD.n949 VDD.n948 9.3
R1537 VDD.n1008 VDD.n1007 9.3
R1538 VDD.n1003 VDD.n1002 9.3
R1539 VDD.n996 VDD.n995 9.3
R1540 VDD.n989 VDD.n988 9.3
R1541 VDD.n1006 VDD.n1005 9.3
R1542 VDD.n1001 VDD.n1000 9.3
R1543 VDD.n999 VDD.n998 9.3
R1544 VDD.n994 VDD.n993 9.3
R1545 VDD.n992 VDD.n991 9.3
R1546 VDD.n987 VDD.n986 9.3
R1547 VDD.n954 VDD.n953 9.3
R1548 VDD.n959 VDD.n958 9.3
R1549 VDD.n966 VDD.n965 9.3
R1550 VDD.n982 VDD.n981 9.3
R1551 VDD.n985 VDD.n984 9.3
R1552 VDD.n1010 VDD.n1009 9.3
R1553 VDD.n1013 VDD.n1012 9.3
R1554 VDD.n940 VDD.n939 9.3
R1555 VDD.n936 VDD.n935 9.3
R1556 VDD.n945 VDD.n944 9.3
R1557 VDD.n1020 VDD.n1019 9.3
R1558 VDD.n1027 VDD.n1026 9.3
R1559 VDD.n1034 VDD.n1033 9.3
R1560 VDD.n1041 VDD.n1040 9.3
R1561 VDD.n1046 VDD.n1045 9.3
R1562 VDD.n1056 VDD.n1055 9.3
R1563 VDD.n1063 VDD.n1062 9.3
R1564 VDD.n1052 VDD.n1051 9.3
R1565 VDD.n1076 VDD.n1075 9.3
R1566 VDD.n1072 VDD.n1071 9.3
R1567 VDD.n1067 VDD.n1066 9.3
R1568 VDD.n1082 VDD.n1081 9.3
R1569 VDD.n1048 VDD.n1047 9.3
R1570 VDD.n1043 VDD.n1042 9.3
R1571 VDD.n1039 VDD.n1038 9.3
R1572 VDD.n1036 VDD.n1035 9.3
R1573 VDD.n1032 VDD.n1031 9.3
R1574 VDD.n1029 VDD.n1028 9.3
R1575 VDD.n1025 VDD.n1024 9.3
R1576 VDD.n1022 VDD.n1021 9.3
R1577 VDD.n1018 VDD.n1017 9.3
R1578 VDD.n1058 VDD.n1057 9.3
R1579 VDD.n1336 VDD.n1335 9.3
R1580 VDD.n1329 VDD.n1328 9.3
R1581 VDD.n1302 VDD.n1301 9.3
R1582 VDD.n1324 VDD.n1323 9.3
R1583 VDD.n1307 VDD.n1306 9.3
R1584 VDD.n1312 VDD.n1311 9.3
R1585 VDD.n1317 VDD.n1316 9.3
R1586 VDD.n1322 VDD.n1321 9.3
R1587 VDD.n1283 VDD.n1282 9.3
R1588 VDD.n1359 VDD.n1358 9.3
R1589 VDD.n1354 VDD.n1353 9.3
R1590 VDD.n1347 VDD.n1346 9.3
R1591 VDD.n1338 VDD.n1337 9.3
R1592 VDD.n1357 VDD.n1356 9.3
R1593 VDD.n1352 VDD.n1351 9.3
R1594 VDD.n1350 VDD.n1349 9.3
R1595 VDD.n1345 VDD.n1344 9.3
R1596 VDD.n1343 VDD.n1342 9.3
R1597 VDD.n1340 VDD.n1339 9.3
R1598 VDD.n1361 VDD.n1360 9.3
R1599 VDD.n1363 VDD.n1362 9.3
R1600 VDD.n1333 VDD.n1332 9.3
R1601 VDD.n1613 VDD.n1612 9.3
R1602 VDD.n1626 VDD.n1625 9.3
R1603 VDD.n1624 VDD.n1623 9.3
R1604 VDD.n1617 VDD.n1616 9.3
R1605 VDD.n1471 VDD.n1470 9.3
R1606 VDD.n1475 VDD.n1474 9.3
R1607 VDD.n1485 VDD.n1484 9.3
R1608 VDD.n1487 VDD.n1486 9.3
R1609 VDD.n1919 VDD.n1918 9.3
R1610 VDD.n1930 VDD.n1929 9.3
R1611 VDD.n1942 VDD.n1941 9.3
R1612 VDD.n1954 VDD.n1953 9.3
R1613 VDD.n1972 VDD.n1971 9.3
R1614 VDD.n1984 VDD.n1983 9.3
R1615 VDD.n1996 VDD.n1995 9.3
R1616 VDD.n2008 VDD.n2007 9.3
R1617 VDD.n2010 VDD.n2009 9.3
R1618 VDD.n1998 VDD.n1997 9.3
R1619 VDD.n1986 VDD.n1985 9.3
R1620 VDD.n1974 VDD.n1973 9.3
R1621 VDD.n1952 VDD.n1951 9.3
R1622 VDD.n1940 VDD.n1939 9.3
R1623 VDD.n1928 VDD.n1927 9.3
R1624 VDD.n1917 VDD.n1916 9.3
R1625 VDD.n2006 VDD.n2005 9.3
R1626 VDD.n2005 VDD.n2004 9.3
R1627 VDD.n1994 VDD.n1993 9.3
R1628 VDD.n1993 VDD.n1992 9.3
R1629 VDD.n1982 VDD.n1981 9.3
R1630 VDD.n1981 VDD.n1980 9.3
R1631 VDD.n1970 VDD.n1969 9.3
R1632 VDD.n1969 VDD.n1968 9.3
R1633 VDD.n1962 VDD.n1961 9.3
R1634 VDD.n1961 VDD.n1960 9.3
R1635 VDD.n1950 VDD.n1949 9.3
R1636 VDD.n1949 VDD.n1948 9.3
R1637 VDD.n1938 VDD.n1937 9.3
R1638 VDD.n1937 VDD.n1936 9.3
R1639 VDD.n1926 VDD.n1925 9.3
R1640 VDD.n1925 VDD.n1924 9.3
R1641 VDD.n556 VDD.n555 9.3
R1642 VDD.n568 VDD.n567 9.3
R1643 VDD.n580 VDD.n579 9.3
R1644 VDD.n593 VDD.n592 9.3
R1645 VDD.n612 VDD.n611 9.3
R1646 VDD.n625 VDD.n624 9.3
R1647 VDD.n637 VDD.n636 9.3
R1648 VDD.n649 VDD.n648 9.3
R1649 VDD.n412 VDD.n411 9.3
R1650 VDD.n434 VDD.n433 9.3
R1651 VDD.n402 VDD.n401 9.3
R1652 VDD.n393 VDD.n392 9.3
R1653 VDD.n383 VDD.n382 9.3
R1654 VDD.n371 VDD.n370 9.3
R1655 VDD.n364 VDD.n363 9.3
R1656 VDD.n352 VDD.n351 9.3
R1657 VDD.n651 VDD.n650 9.3
R1658 VDD.n647 VDD.n646 9.3
R1659 VDD.n646 VDD.n645 9.3
R1660 VDD.n639 VDD.n638 9.3
R1661 VDD.n635 VDD.n634 9.3
R1662 VDD.n634 VDD.n633 9.3
R1663 VDD.n627 VDD.n626 9.3
R1664 VDD.n623 VDD.n622 9.3
R1665 VDD.n622 VDD.n621 9.3
R1666 VDD.n614 VDD.n613 9.3
R1667 VDD.n610 VDD.n609 9.3
R1668 VDD.n609 VDD.n608 9.3
R1669 VDD.n601 VDD.n600 9.3
R1670 VDD.n600 VDD.n599 9.3
R1671 VDD.n591 VDD.n590 9.3
R1672 VDD.n589 VDD.n588 9.3
R1673 VDD.n588 VDD.n587 9.3
R1674 VDD.n578 VDD.n577 9.3
R1675 VDD.n576 VDD.n575 9.3
R1676 VDD.n575 VDD.n574 9.3
R1677 VDD.n566 VDD.n565 9.3
R1678 VDD.n564 VDD.n563 9.3
R1679 VDD.n563 VDD.n562 9.3
R1680 VDD.n554 VDD.n553 9.3
R1681 VDD.n194 VDD.n193 9.3
R1682 VDD.n182 VDD.n181 9.3
R1683 VDD.n241 VDD.n240 9.3
R1684 VDD.n236 VDD.n235 9.3
R1685 VDD.n229 VDD.n228 9.3
R1686 VDD.n222 VDD.n221 9.3
R1687 VDD.n239 VDD.n238 9.3
R1688 VDD.n234 VDD.n233 9.3
R1689 VDD.n232 VDD.n231 9.3
R1690 VDD.n227 VDD.n226 9.3
R1691 VDD.n225 VDD.n224 9.3
R1692 VDD.n220 VDD.n219 9.3
R1693 VDD.n187 VDD.n186 9.3
R1694 VDD.n192 VDD.n191 9.3
R1695 VDD.n199 VDD.n198 9.3
R1696 VDD.n215 VDD.n214 9.3
R1697 VDD.n218 VDD.n217 9.3
R1698 VDD.n243 VDD.n242 9.3
R1699 VDD.n247 VDD.n246 9.3
R1700 VDD.n173 VDD.n172 9.3
R1701 VDD.n169 VDD.n168 9.3
R1702 VDD.n178 VDD.n177 9.3
R1703 VDD.n2157 VDD.n2156 9.3
R1704 VDD.n2163 VDD.n2162 9.3
R1705 VDD.n2188 VDD.n2187 9.3
R1706 VDD.n2167 VDD.n2166 9.3
R1707 VDD.n2184 VDD.n2183 9.3
R1708 VDD.n2178 VDD.n2177 9.3
R1709 VDD.n2174 VDD.n2173 9.3
R1710 VDD.n2169 VDD.n2168 9.3
R1711 VDD.n2194 VDD.n2193 9.3
R1712 VDD.n2133 VDD.n2132 9.3
R1713 VDD.n2138 VDD.n2137 9.3
R1714 VDD.n2145 VDD.n2144 9.3
R1715 VDD.n2154 VDD.n2153 9.3
R1716 VDD.n2136 VDD.n2135 9.3
R1717 VDD.n2140 VDD.n2139 9.3
R1718 VDD.n2143 VDD.n2142 9.3
R1719 VDD.n2147 VDD.n2146 9.3
R1720 VDD.n2150 VDD.n2149 9.3
R1721 VDD.n2152 VDD.n2151 9.3
R1722 VDD.n2131 VDD.n2130 9.3
R1723 VDD.n2129 VDD.n2128 9.3
R1724 VDD.n2159 VDD.n2158 9.3
R1725 VDD.n538 VDD.n537 9.3
R1726 VDD.n531 VDD.n530 9.3
R1727 VDD.n524 VDD.n523 9.3
R1728 VDD.n517 VDD.n516 9.3
R1729 VDD.n513 VDD.n512 9.3
R1730 VDD.n501 VDD.n500 9.3
R1731 VDD.n494 VDD.n493 9.3
R1732 VDD.n506 VDD.n505 9.3
R1733 VDD.n479 VDD.n478 9.3
R1734 VDD.n484 VDD.n483 9.3
R1735 VDD.n489 VDD.n488 9.3
R1736 VDD.n460 VDD.n459 9.3
R1737 VDD.n510 VDD.n509 9.3
R1738 VDD.n515 VDD.n514 9.3
R1739 VDD.n520 VDD.n519 9.3
R1740 VDD.n522 VDD.n521 9.3
R1741 VDD.n527 VDD.n526 9.3
R1742 VDD.n529 VDD.n528 9.3
R1743 VDD.n534 VDD.n533 9.3
R1744 VDD.n536 VDD.n535 9.3
R1745 VDD.n540 VDD.n539 9.3
R1746 VDD.n499 VDD.n498 9.3
R1747 VDD.n2126 VDD.n2125 9.3
R1748 VDD.n546 VDD.n545 9.3
R1749 VDD.n544 VDD.n543 9.3
R1750 VDD.n2124 VDD.n2123 9.3
R1751 VDD.n2116 VDD.n2115 9.3
R1752 VDD.n2104 VDD.n2103 9.3
R1753 VDD.n2092 VDD.n2091 9.3
R1754 VDD.n2080 VDD.n2079 9.3
R1755 VDD.n2062 VDD.n2061 9.3
R1756 VDD.n2050 VDD.n2049 9.3
R1757 VDD.n2038 VDD.n2037 9.3
R1758 VDD.n2024 VDD.n2023 9.3
R1759 VDD.n2118 VDD.n2117 9.3
R1760 VDD.n2114 VDD.n2113 9.3
R1761 VDD.n2113 VDD.n2112 9.3
R1762 VDD.n2106 VDD.n2105 9.3
R1763 VDD.n2102 VDD.n2101 9.3
R1764 VDD.n2101 VDD.n2100 9.3
R1765 VDD.n2094 VDD.n2093 9.3
R1766 VDD.n2090 VDD.n2089 9.3
R1767 VDD.n2089 VDD.n2088 9.3
R1768 VDD.n2082 VDD.n2081 9.3
R1769 VDD.n2078 VDD.n2077 9.3
R1770 VDD.n2077 VDD.n2076 9.3
R1771 VDD.n2070 VDD.n2069 9.3
R1772 VDD.n2069 VDD.n2068 9.3
R1773 VDD.n2060 VDD.n2059 9.3
R1774 VDD.n2058 VDD.n2057 9.3
R1775 VDD.n2057 VDD.n2056 9.3
R1776 VDD.n2048 VDD.n2047 9.3
R1777 VDD.n2046 VDD.n2045 9.3
R1778 VDD.n2045 VDD.n2044 9.3
R1779 VDD.n2036 VDD.n2035 9.3
R1780 VDD.n2034 VDD.n2033 9.3
R1781 VDD.n2033 VDD.n2032 9.3
R1782 VDD.n2026 VDD.n2025 9.3
R1783 VDD.n3461 VDD.n3460 9.3
R1784 VDD.n3472 VDD.n3471 9.3
R1785 VDD.n3485 VDD.n3484 9.3
R1786 VDD.n3497 VDD.n3496 9.3
R1787 VDD.n3515 VDD.n3514 9.3
R1788 VDD.n3527 VDD.n3526 9.3
R1789 VDD.n3539 VDD.n3538 9.3
R1790 VDD.n3551 VDD.n3550 9.3
R1791 VDD.n3582 VDD.n3581 9.3
R1792 VDD.n331 VDD.n330 9.3
R1793 VDD.n266 VDD.n265 9.3
R1794 VDD.n322 VDD.n321 9.3
R1795 VDD.n316 VDD.n315 9.3
R1796 VDD.n335 VDD.n316 9.3
R1797 VDD.n278 VDD.n277 9.3
R1798 VDD.n335 VDD.n278 9.3
R1799 VDD.n307 VDD.n306 9.3
R1800 VDD.n335 VDD.n307 9.3
R1801 VDD.n295 VDD.n294 9.3
R1802 VDD.n3553 VDD.n3552 9.3
R1803 VDD.n3549 VDD.n3548 9.3
R1804 VDD.n3548 VDD.n3547 9.3
R1805 VDD.n3541 VDD.n3540 9.3
R1806 VDD.n3537 VDD.n3536 9.3
R1807 VDD.n3536 VDD.n3535 9.3
R1808 VDD.n3529 VDD.n3528 9.3
R1809 VDD.n3525 VDD.n3524 9.3
R1810 VDD.n3524 VDD.n3523 9.3
R1811 VDD.n3517 VDD.n3516 9.3
R1812 VDD.n3513 VDD.n3512 9.3
R1813 VDD.n3512 VDD.n3511 9.3
R1814 VDD.n3505 VDD.n3504 9.3
R1815 VDD.n3504 VDD.n3503 9.3
R1816 VDD.n3495 VDD.n3494 9.3
R1817 VDD.n3493 VDD.n3492 9.3
R1818 VDD.n3492 VDD.n3491 9.3
R1819 VDD.n3483 VDD.n3482 9.3
R1820 VDD.n3481 VDD.n3480 9.3
R1821 VDD.n3480 VDD.n3479 9.3
R1822 VDD.n3470 VDD.n3469 9.3
R1823 VDD.n3459 VDD.n3458 9.3
R1824 VDD.n3468 VDD.n3467 9.3
R1825 VDD.n3467 VDD.n3466 9.3
R1826 VDD.n2352 VDD.n2351 9.3
R1827 VDD.n2341 VDD.n2340 9.3
R1828 VDD.n2329 VDD.n2328 9.3
R1829 VDD.n2317 VDD.n2316 9.3
R1830 VDD.n2299 VDD.n2298 9.3
R1831 VDD.n2287 VDD.n2286 9.3
R1832 VDD.n2275 VDD.n2274 9.3
R1833 VDD.n2263 VDD.n2262 9.3
R1834 VDD.n2232 VDD.n2231 9.3
R1835 VDD.n738 VDD.n737 9.3
R1836 VDD.n672 VDD.n671 9.3
R1837 VDD.n729 VDD.n728 9.3
R1838 VDD.n723 VDD.n722 9.3
R1839 VDD.n742 VDD.n723 9.3
R1840 VDD.n684 VDD.n683 9.3
R1841 VDD.n742 VDD.n684 9.3
R1842 VDD.n714 VDD.n713 9.3
R1843 VDD.n742 VDD.n714 9.3
R1844 VDD.n702 VDD.n701 9.3
R1845 VDD.n2261 VDD.n2260 9.3
R1846 VDD.n2271 VDD.n2270 9.3
R1847 VDD.n2270 VDD.n2269 9.3
R1848 VDD.n2273 VDD.n2272 9.3
R1849 VDD.n2283 VDD.n2282 9.3
R1850 VDD.n2282 VDD.n2281 9.3
R1851 VDD.n2285 VDD.n2284 9.3
R1852 VDD.n2295 VDD.n2294 9.3
R1853 VDD.n2294 VDD.n2293 9.3
R1854 VDD.n2297 VDD.n2296 9.3
R1855 VDD.n2307 VDD.n2306 9.3
R1856 VDD.n2306 VDD.n2305 9.3
R1857 VDD.n2315 VDD.n2314 9.3
R1858 VDD.n2314 VDD.n2313 9.3
R1859 VDD.n2319 VDD.n2318 9.3
R1860 VDD.n2327 VDD.n2326 9.3
R1861 VDD.n2326 VDD.n2325 9.3
R1862 VDD.n2331 VDD.n2330 9.3
R1863 VDD.n2339 VDD.n2338 9.3
R1864 VDD.n2338 VDD.n2337 9.3
R1865 VDD.n2343 VDD.n2342 9.3
R1866 VDD.n2354 VDD.n2353 9.3
R1867 VDD.n2350 VDD.n2349 9.3
R1868 VDD.n2349 VDD.n2348 9.3
R1869 VDD.n1694 VDD.n1693 9.3
R1870 VDD.n1687 VDD.n1686 9.3
R1871 VDD.n1660 VDD.n1659 9.3
R1872 VDD.n1682 VDD.n1681 9.3
R1873 VDD.n1665 VDD.n1664 9.3
R1874 VDD.n1670 VDD.n1669 9.3
R1875 VDD.n1675 VDD.n1674 9.3
R1876 VDD.n1680 VDD.n1679 9.3
R1877 VDD.n1641 VDD.n1640 9.3
R1878 VDD.n1717 VDD.n1716 9.3
R1879 VDD.n1712 VDD.n1711 9.3
R1880 VDD.n1705 VDD.n1704 9.3
R1881 VDD.n1696 VDD.n1695 9.3
R1882 VDD.n1715 VDD.n1714 9.3
R1883 VDD.n1710 VDD.n1709 9.3
R1884 VDD.n1708 VDD.n1707 9.3
R1885 VDD.n1703 VDD.n1702 9.3
R1886 VDD.n1701 VDD.n1700 9.3
R1887 VDD.n1698 VDD.n1697 9.3
R1888 VDD.n1719 VDD.n1718 9.3
R1889 VDD.n1721 VDD.n1720 9.3
R1890 VDD.n1691 VDD.n1690 9.3
R1891 VDD.n1850 VDD.n1849 9.3
R1892 VDD.n1846 VDD.n1845 9.3
R1893 VDD.n1862 VDD.n1861 9.3
R1894 VDD.n1864 VDD.n1863 9.3
R1895 VDD.n1264 VDD.n1263 9.3
R1896 VDD.n1257 VDD.n1256 9.3
R1897 VDD.n1250 VDD.n1249 9.3
R1898 VDD.n1243 VDD.n1242 9.3
R1899 VDD.n1239 VDD.n1238 9.3
R1900 VDD.n1227 VDD.n1226 9.3
R1901 VDD.n1220 VDD.n1219 9.3
R1902 VDD.n1232 VDD.n1231 9.3
R1903 VDD.n1205 VDD.n1204 9.3
R1904 VDD.n1210 VDD.n1209 9.3
R1905 VDD.n1215 VDD.n1214 9.3
R1906 VDD.n1200 VDD.n1199 9.3
R1907 VDD.n1236 VDD.n1235 9.3
R1908 VDD.n1241 VDD.n1240 9.3
R1909 VDD.n1246 VDD.n1245 9.3
R1910 VDD.n1248 VDD.n1247 9.3
R1911 VDD.n1253 VDD.n1252 9.3
R1912 VDD.n1255 VDD.n1254 9.3
R1913 VDD.n1260 VDD.n1259 9.3
R1914 VDD.n1262 VDD.n1261 9.3
R1915 VDD.n1266 VDD.n1265 9.3
R1916 VDD.n1225 VDD.n1224 9.3
R1917 VDD.n1727 VDD.n1726 9.3
R1918 VDD.n1272 VDD.n1271 9.3
R1919 VDD.n1270 VDD.n1269 9.3
R1920 VDD.n1725 VDD.n1724 9.3
R1921 VDD.n1514 VDD.n1513 9.3
R1922 VDD.n1526 VDD.n1525 9.3
R1923 VDD.n1538 VDD.n1537 9.3
R1924 VDD.n1550 VDD.n1549 9.3
R1925 VDD.n1569 VDD.n1568 9.3
R1926 VDD.n1581 VDD.n1580 9.3
R1927 VDD.n1593 VDD.n1592 9.3
R1928 VDD.n1605 VDD.n1604 9.3
R1929 VDD.n1174 VDD.n1173 9.3
R1930 VDD.n1607 VDD.n1606 9.3
R1931 VDD.n1595 VDD.n1594 9.3
R1932 VDD.n1583 VDD.n1582 9.3
R1933 VDD.n1571 VDD.n1570 9.3
R1934 VDD.n1548 VDD.n1547 9.3
R1935 VDD.n1536 VDD.n1535 9.3
R1936 VDD.n1524 VDD.n1523 9.3
R1937 VDD.n1512 VDD.n1511 9.3
R1938 VDD.n1162 VDD.n1161 9.3
R1939 VDD.n1093 VDD.n1092 9.3
R1940 VDD.n1153 VDD.n1152 9.3
R1941 VDD.n1147 VDD.n1146 9.3
R1942 VDD.n1166 VDD.n1147 9.3
R1943 VDD.n1105 VDD.n1104 9.3
R1944 VDD.n1166 VDD.n1105 9.3
R1945 VDD.n1138 VDD.n1137 9.3
R1946 VDD.n1166 VDD.n1138 9.3
R1947 VDD.n1114 VDD.n1113 9.3
R1948 VDD.n1603 VDD.n1602 9.3
R1949 VDD.n1602 VDD.n1601 9.3
R1950 VDD.n1591 VDD.n1590 9.3
R1951 VDD.n1590 VDD.n1589 9.3
R1952 VDD.n1579 VDD.n1578 9.3
R1953 VDD.n1578 VDD.n1577 9.3
R1954 VDD.n1567 VDD.n1566 9.3
R1955 VDD.n1566 VDD.n1565 9.3
R1956 VDD.n1559 VDD.n1558 9.3
R1957 VDD.n1558 VDD.n1557 9.3
R1958 VDD.n1546 VDD.n1545 9.3
R1959 VDD.n1545 VDD.n1544 9.3
R1960 VDD.n1534 VDD.n1533 9.3
R1961 VDD.n1533 VDD.n1532 9.3
R1962 VDD.n1522 VDD.n1521 9.3
R1963 VDD.n1521 VDD.n1520 9.3
R1964 VDD.n1826 VDD.n1825 9.3
R1965 VDD.n1814 VDD.n1813 9.3
R1966 VDD.n1802 VDD.n1801 9.3
R1967 VDD.n1790 VDD.n1789 9.3
R1968 VDD.n1772 VDD.n1771 9.3
R1969 VDD.n1760 VDD.n1759 9.3
R1970 VDD.n1748 VDD.n1747 9.3
R1971 VDD.n1736 VDD.n1735 9.3
R1972 VDD.n1367 VDD.n1366 9.3
R1973 VDD.n1379 VDD.n1378 9.3
R1974 VDD.n1391 VDD.n1390 9.3
R1975 VDD.n1403 VDD.n1402 9.3
R1976 VDD.n1421 VDD.n1420 9.3
R1977 VDD.n1433 VDD.n1432 9.3
R1978 VDD.n1445 VDD.n1444 9.3
R1979 VDD.n1457 VDD.n1456 9.3
R1980 VDD.n1828 VDD.n1827 9.3
R1981 VDD.n1824 VDD.n1823 9.3
R1982 VDD.n1823 VDD.n1822 9.3
R1983 VDD.n1459 VDD.n1458 9.3
R1984 VDD.n1455 VDD.n1454 9.3
R1985 VDD.n1454 VDD.n1453 9.3
R1986 VDD.n1447 VDD.n1446 9.3
R1987 VDD.n1443 VDD.n1442 9.3
R1988 VDD.n1442 VDD.n1441 9.3
R1989 VDD.n1435 VDD.n1434 9.3
R1990 VDD.n1431 VDD.n1430 9.3
R1991 VDD.n1430 VDD.n1429 9.3
R1992 VDD.n1423 VDD.n1422 9.3
R1993 VDD.n1419 VDD.n1418 9.3
R1994 VDD.n1418 VDD.n1417 9.3
R1995 VDD.n1411 VDD.n1410 9.3
R1996 VDD.n1410 VDD.n1409 9.3
R1997 VDD.n1401 VDD.n1400 9.3
R1998 VDD.n1399 VDD.n1398 9.3
R1999 VDD.n1398 VDD.n1397 9.3
R2000 VDD.n1389 VDD.n1388 9.3
R2001 VDD.n1387 VDD.n1386 9.3
R2002 VDD.n1386 VDD.n1385 9.3
R2003 VDD.n1377 VDD.n1376 9.3
R2004 VDD.n1375 VDD.n1374 9.3
R2005 VDD.n1374 VDD.n1373 9.3
R2006 VDD.n1365 VDD.n1364 9.3
R2007 VDD.n1734 VDD.n1733 9.3
R2008 VDD.n1744 VDD.n1743 9.3
R2009 VDD.n1743 VDD.n1742 9.3
R2010 VDD.n1746 VDD.n1745 9.3
R2011 VDD.n1756 VDD.n1755 9.3
R2012 VDD.n1755 VDD.n1754 9.3
R2013 VDD.n1758 VDD.n1757 9.3
R2014 VDD.n1768 VDD.n1767 9.3
R2015 VDD.n1767 VDD.n1766 9.3
R2016 VDD.n1770 VDD.n1769 9.3
R2017 VDD.n1780 VDD.n1779 9.3
R2018 VDD.n1779 VDD.n1778 9.3
R2019 VDD.n1788 VDD.n1787 9.3
R2020 VDD.n1787 VDD.n1786 9.3
R2021 VDD.n1792 VDD.n1791 9.3
R2022 VDD.n1800 VDD.n1799 9.3
R2023 VDD.n1799 VDD.n1798 9.3
R2024 VDD.n1804 VDD.n1803 9.3
R2025 VDD.n1812 VDD.n1811 9.3
R2026 VDD.n1811 VDD.n1810 9.3
R2027 VDD.n1816 VDD.n1815 9.3
R2028 VDD.n3289 VDD.n3288 9.3
R2029 VDD.n3277 VDD.n3276 9.3
R2030 VDD.n3265 VDD.n3264 9.3
R2031 VDD.n3253 VDD.n3252 9.3
R2032 VDD.n3235 VDD.n3234 9.3
R2033 VDD.n3223 VDD.n3222 9.3
R2034 VDD.n3210 VDD.n3209 9.3
R2035 VDD.n3208 VDD.n3207 9.3
R2036 VDD.n3219 VDD.n3218 9.3
R2037 VDD.n3218 VDD.n3217 9.3
R2038 VDD.n3221 VDD.n3220 9.3
R2039 VDD.n3231 VDD.n3230 9.3
R2040 VDD.n3230 VDD.n3229 9.3
R2041 VDD.n3233 VDD.n3232 9.3
R2042 VDD.n3243 VDD.n3242 9.3
R2043 VDD.n3242 VDD.n3241 9.3
R2044 VDD.n3251 VDD.n3250 9.3
R2045 VDD.n3250 VDD.n3249 9.3
R2046 VDD.n3255 VDD.n3254 9.3
R2047 VDD.n3263 VDD.n3262 9.3
R2048 VDD.n3262 VDD.n3261 9.3
R2049 VDD.n3267 VDD.n3266 9.3
R2050 VDD.n3275 VDD.n3274 9.3
R2051 VDD.n3274 VDD.n3273 9.3
R2052 VDD.n3279 VDD.n3278 9.3
R2053 VDD.n3287 VDD.n3286 9.3
R2054 VDD.n3286 VDD.n3285 9.3
R2055 VDD.n3291 VDD.n3290 9.3
R2056 VDD.n3206 VDD.n3205 9.3
R2057 VDD.n3205 VDD.n3204 9.3
R2058 VDD.n3196 VDD.n3195 9.3
R2059 VDD.n3198 VDD.n3197 9.3
R2060 VDD.n3413 VDD.n3412 9.3
R2061 VDD.n3401 VDD.n3400 9.3
R2062 VDD.n3389 VDD.n3388 9.3
R2063 VDD.n3376 VDD.n3375 9.3
R2064 VDD.n3357 VDD.n3356 9.3
R2065 VDD.n3344 VDD.n3343 9.3
R2066 VDD.n3332 VDD.n3331 9.3
R2067 VDD.n3320 VDD.n3319 9.3
R2068 VDD.n2979 VDD.n2978 9.3
R2069 VDD.n3055 VDD.n3054 9.3
R2070 VDD.n2989 VDD.n2988 9.3
R2071 VDD.n3046 VDD.n3045 9.3
R2072 VDD.n3040 VDD.n3039 9.3
R2073 VDD.n3059 VDD.n3040 9.3
R2074 VDD.n3001 VDD.n3000 9.3
R2075 VDD.n3059 VDD.n3001 9.3
R2076 VDD.n3031 VDD.n3030 9.3
R2077 VDD.n3059 VDD.n3031 9.3
R2078 VDD.n3010 VDD.n3009 9.3
R2079 VDD.n3318 VDD.n3317 9.3
R2080 VDD.n3328 VDD.n3327 9.3
R2081 VDD.n3327 VDD.n3326 9.3
R2082 VDD.n3330 VDD.n3329 9.3
R2083 VDD.n3340 VDD.n3339 9.3
R2084 VDD.n3339 VDD.n3338 9.3
R2085 VDD.n3342 VDD.n3341 9.3
R2086 VDD.n3353 VDD.n3352 9.3
R2087 VDD.n3352 VDD.n3351 9.3
R2088 VDD.n3355 VDD.n3354 9.3
R2089 VDD.n3365 VDD.n3364 9.3
R2090 VDD.n3364 VDD.n3363 9.3
R2091 VDD.n3374 VDD.n3373 9.3
R2092 VDD.n3373 VDD.n3372 9.3
R2093 VDD.n3378 VDD.n3377 9.3
R2094 VDD.n3387 VDD.n3386 9.3
R2095 VDD.n3386 VDD.n3385 9.3
R2096 VDD.n3391 VDD.n3390 9.3
R2097 VDD.n3399 VDD.n3398 9.3
R2098 VDD.n3398 VDD.n3397 9.3
R2099 VDD.n3403 VDD.n3402 9.3
R2100 VDD.n3411 VDD.n3410 9.3
R2101 VDD.n3410 VDD.n3409 9.3
R2102 VDD.n3415 VDD.n3414 9.3
R2103 VDD.n2717 VDD.n2716 9.3
R2104 VDD.n2723 VDD.n2722 9.3
R2105 VDD.n2748 VDD.n2747 9.3
R2106 VDD.n2727 VDD.n2726 9.3
R2107 VDD.n2744 VDD.n2743 9.3
R2108 VDD.n2738 VDD.n2737 9.3
R2109 VDD.n2734 VDD.n2733 9.3
R2110 VDD.n2729 VDD.n2728 9.3
R2111 VDD.n2754 VDD.n2753 9.3
R2112 VDD.n2693 VDD.n2692 9.3
R2113 VDD.n2698 VDD.n2697 9.3
R2114 VDD.n2705 VDD.n2704 9.3
R2115 VDD.n2714 VDD.n2713 9.3
R2116 VDD.n2696 VDD.n2695 9.3
R2117 VDD.n2700 VDD.n2699 9.3
R2118 VDD.n2703 VDD.n2702 9.3
R2119 VDD.n2707 VDD.n2706 9.3
R2120 VDD.n2710 VDD.n2709 9.3
R2121 VDD.n2712 VDD.n2711 9.3
R2122 VDD.n2691 VDD.n2690 9.3
R2123 VDD.n2689 VDD.n2688 9.3
R2124 VDD.n2719 VDD.n2718 9.3
R2125 VDD.n2943 VDD.n2942 9.3
R2126 VDD.n2936 VDD.n2935 9.3
R2127 VDD.n2929 VDD.n2928 9.3
R2128 VDD.n2922 VDD.n2921 9.3
R2129 VDD.n2918 VDD.n2917 9.3
R2130 VDD.n2906 VDD.n2905 9.3
R2131 VDD.n2899 VDD.n2898 9.3
R2132 VDD.n2911 VDD.n2910 9.3
R2133 VDD.n2884 VDD.n2883 9.3
R2134 VDD.n2889 VDD.n2888 9.3
R2135 VDD.n2894 VDD.n2893 9.3
R2136 VDD.n2865 VDD.n2864 9.3
R2137 VDD.n2915 VDD.n2914 9.3
R2138 VDD.n2920 VDD.n2919 9.3
R2139 VDD.n2925 VDD.n2924 9.3
R2140 VDD.n2927 VDD.n2926 9.3
R2141 VDD.n2932 VDD.n2931 9.3
R2142 VDD.n2934 VDD.n2933 9.3
R2143 VDD.n2939 VDD.n2938 9.3
R2144 VDD.n2941 VDD.n2940 9.3
R2145 VDD.n2945 VDD.n2944 9.3
R2146 VDD.n2904 VDD.n2903 9.3
R2147 VDD.n2686 VDD.n2685 9.3
R2148 VDD.n2951 VDD.n2950 9.3
R2149 VDD.n2949 VDD.n2948 9.3
R2150 VDD.n2684 VDD.n2683 9.3
R2151 VDD.n3094 VDD.n3093 9.3
R2152 VDD.n3106 VDD.n3105 9.3
R2153 VDD.n3118 VDD.n3117 9.3
R2154 VDD.n3130 VDD.n3129 9.3
R2155 VDD.n3148 VDD.n3147 9.3
R2156 VDD.n3160 VDD.n3159 9.3
R2157 VDD.n3172 VDD.n3171 9.3
R2158 VDD.n3184 VDD.n3183 9.3
R2159 VDD.n3092 VDD.n3091 9.3
R2160 VDD.n3102 VDD.n3101 9.3
R2161 VDD.n3101 VDD.n3100 9.3
R2162 VDD.n3104 VDD.n3103 9.3
R2163 VDD.n3114 VDD.n3113 9.3
R2164 VDD.n3113 VDD.n3112 9.3
R2165 VDD.n3116 VDD.n3115 9.3
R2166 VDD.n3126 VDD.n3125 9.3
R2167 VDD.n3125 VDD.n3124 9.3
R2168 VDD.n3128 VDD.n3127 9.3
R2169 VDD.n3138 VDD.n3137 9.3
R2170 VDD.n3137 VDD.n3136 9.3
R2171 VDD.n3146 VDD.n3145 9.3
R2172 VDD.n3145 VDD.n3144 9.3
R2173 VDD.n3150 VDD.n3149 9.3
R2174 VDD.n3158 VDD.n3157 9.3
R2175 VDD.n3157 VDD.n3156 9.3
R2176 VDD.n3162 VDD.n3161 9.3
R2177 VDD.n3170 VDD.n3169 9.3
R2178 VDD.n3169 VDD.n3168 9.3
R2179 VDD.n3174 VDD.n3173 9.3
R2180 VDD.n3182 VDD.n3181 9.3
R2181 VDD.n3181 VDD.n3180 9.3
R2182 VDD.n3186 VDD.n3185 9.3
R2183 VDD.n3758 VDD.n3757 9.3
R2184 VDD.n3735 VDD.n3734 9.3
R2185 VDD.n3743 VDD.n3742 9.3
R2186 VDD.n3747 VDD.n3746 9.3
R2187 VDD.n3770 VDD.n3769 9.3
R2188 VDD.n3765 VDD.n3764 9.3
R2189 VDD.n3762 VDD.n3761 9.3
R2190 VDD.n3731 VDD.n3730 9.3
R2191 VDD.n3800 VDD.n3799 9.3
R2192 VDD.n3777 VDD.n3776 9.3
R2193 VDD.n3785 VDD.n3784 9.3
R2194 VDD.n3789 VDD.n3788 9.3
R2195 VDD.n3812 VDD.n3811 9.3
R2196 VDD.n3807 VDD.n3806 9.3
R2197 VDD.n3804 VDD.n3803 9.3
R2198 VDD.n3773 VDD.n3772 9.3
R2199 VDD.n3911 VDD.n3910 9.3
R2200 VDD.n3888 VDD.n3887 9.3
R2201 VDD.n3896 VDD.n3895 9.3
R2202 VDD.n3900 VDD.n3899 9.3
R2203 VDD.n3923 VDD.n3922 9.3
R2204 VDD.n3918 VDD.n3917 9.3
R2205 VDD.n3915 VDD.n3914 9.3
R2206 VDD.n3884 VDD.n3883 9.3
R2207 VDD.n3859 VDD.n3858 9.3
R2208 VDD.n3863 VDD.n3862 9.3
R2209 VDD.n3866 VDD.n3865 9.3
R2210 VDD.n3871 VDD.n3870 9.3
R2211 VDD.n3848 VDD.n3847 9.3
R2212 VDD.n3844 VDD.n3843 9.3
R2213 VDD.n3836 VDD.n3835 9.3
R2214 VDD.n3832 VDD.n3831 9.3
R2215 VDD.n4022 VDD.n4021 9.3
R2216 VDD.n3999 VDD.n3998 9.3
R2217 VDD.n4007 VDD.n4006 9.3
R2218 VDD.n4011 VDD.n4010 9.3
R2219 VDD.n4034 VDD.n4033 9.3
R2220 VDD.n4029 VDD.n4028 9.3
R2221 VDD.n4026 VDD.n4025 9.3
R2222 VDD.n3995 VDD.n3994 9.3
R2223 VDD.n3970 VDD.n3969 9.3
R2224 VDD.n3974 VDD.n3973 9.3
R2225 VDD.n3977 VDD.n3976 9.3
R2226 VDD.n3982 VDD.n3981 9.3
R2227 VDD.n3959 VDD.n3958 9.3
R2228 VDD.n3955 VDD.n3954 9.3
R2229 VDD.n3947 VDD.n3946 9.3
R2230 VDD.n3943 VDD.n3942 9.3
R2231 VDD.n4133 VDD.n4132 9.3
R2232 VDD.n4110 VDD.n4109 9.3
R2233 VDD.n4118 VDD.n4117 9.3
R2234 VDD.n4122 VDD.n4121 9.3
R2235 VDD.n4145 VDD.n4144 9.3
R2236 VDD.n4140 VDD.n4139 9.3
R2237 VDD.n4137 VDD.n4136 9.3
R2238 VDD.n4106 VDD.n4105 9.3
R2239 VDD.n4081 VDD.n4080 9.3
R2240 VDD.n4085 VDD.n4084 9.3
R2241 VDD.n4088 VDD.n4087 9.3
R2242 VDD.n4093 VDD.n4092 9.3
R2243 VDD.n4070 VDD.n4069 9.3
R2244 VDD.n4066 VDD.n4065 9.3
R2245 VDD.n4058 VDD.n4057 9.3
R2246 VDD.n4054 VDD.n4053 9.3
R2247 VDD.n4244 VDD.n4243 9.3
R2248 VDD.n4221 VDD.n4220 9.3
R2249 VDD.n4229 VDD.n4228 9.3
R2250 VDD.n4233 VDD.n4232 9.3
R2251 VDD.n4256 VDD.n4255 9.3
R2252 VDD.n4251 VDD.n4250 9.3
R2253 VDD.n4248 VDD.n4247 9.3
R2254 VDD.n4217 VDD.n4216 9.3
R2255 VDD.n4192 VDD.n4191 9.3
R2256 VDD.n4196 VDD.n4195 9.3
R2257 VDD.n4199 VDD.n4198 9.3
R2258 VDD.n4204 VDD.n4203 9.3
R2259 VDD.n4181 VDD.n4180 9.3
R2260 VDD.n4177 VDD.n4176 9.3
R2261 VDD.n4169 VDD.n4168 9.3
R2262 VDD.n4165 VDD.n4164 9.3
R2263 VDD.n4360 VDD.n4359 9.3
R2264 VDD.n4337 VDD.n4336 9.3
R2265 VDD.n4345 VDD.n4344 9.3
R2266 VDD.n4349 VDD.n4348 9.3
R2267 VDD.n4372 VDD.n4371 9.3
R2268 VDD.n4367 VDD.n4366 9.3
R2269 VDD.n4364 VDD.n4363 9.3
R2270 VDD.n4333 VDD.n4332 9.3
R2271 VDD.n4402 VDD.n4401 9.3
R2272 VDD.n4379 VDD.n4378 9.3
R2273 VDD.n4387 VDD.n4386 9.3
R2274 VDD.n4391 VDD.n4390 9.3
R2275 VDD.n4414 VDD.n4413 9.3
R2276 VDD.n4409 VDD.n4408 9.3
R2277 VDD.n4406 VDD.n4405 9.3
R2278 VDD.n4375 VDD.n4374 9.3
R2279 VDD.n4520 VDD.n4519 9.3
R2280 VDD.n4497 VDD.n4496 9.3
R2281 VDD.n4505 VDD.n4504 9.3
R2282 VDD.n4509 VDD.n4508 9.3
R2283 VDD.n4532 VDD.n4531 9.3
R2284 VDD.n4527 VDD.n4526 9.3
R2285 VDD.n4524 VDD.n4523 9.3
R2286 VDD.n4493 VDD.n4492 9.3
R2287 VDD.n4468 VDD.n4467 9.3
R2288 VDD.n4472 VDD.n4471 9.3
R2289 VDD.n4475 VDD.n4474 9.3
R2290 VDD.n4480 VDD.n4479 9.3
R2291 VDD.n4457 VDD.n4456 9.3
R2292 VDD.n4453 VDD.n4452 9.3
R2293 VDD.n4445 VDD.n4444 9.3
R2294 VDD.n4441 VDD.n4440 9.3
R2295 VDD.n4638 VDD.n4637 9.3
R2296 VDD.n4615 VDD.n4614 9.3
R2297 VDD.n4623 VDD.n4622 9.3
R2298 VDD.n4627 VDD.n4626 9.3
R2299 VDD.n4650 VDD.n4649 9.3
R2300 VDD.n4645 VDD.n4644 9.3
R2301 VDD.n4642 VDD.n4641 9.3
R2302 VDD.n4611 VDD.n4610 9.3
R2303 VDD.n4586 VDD.n4585 9.3
R2304 VDD.n4590 VDD.n4589 9.3
R2305 VDD.n4593 VDD.n4592 9.3
R2306 VDD.n4598 VDD.n4597 9.3
R2307 VDD.n4575 VDD.n4574 9.3
R2308 VDD.n4571 VDD.n4570 9.3
R2309 VDD.n4563 VDD.n4562 9.3
R2310 VDD.n4559 VDD.n4558 9.3
R2311 VDD.n4691 VDD.n4690 9.3
R2312 VDD.n4668 VDD.n4667 9.3
R2313 VDD.n4676 VDD.n4675 9.3
R2314 VDD.n4680 VDD.n4679 9.3
R2315 VDD.n4703 VDD.n4702 9.3
R2316 VDD.n4698 VDD.n4697 9.3
R2317 VDD.n4695 VDD.n4694 9.3
R2318 VDD.n4664 VDD.n4663 9.3
R2319 VDD.n28 VDD.n27 9.3
R2320 VDD.n32 VDD.n31 9.3
R2321 VDD.n35 VDD.n34 9.3
R2322 VDD.n40 VDD.n39 9.3
R2323 VDD.n17 VDD.n16 9.3
R2324 VDD.n13 VDD.n12 9.3
R2325 VDD.n5 VDD.n4 9.3
R2326 VDD.n1 VDD.n0 9.3
R2327 VDD.n2840 VDD.n2839 9.162
R2328 VDD.n2840 VDD.t10 9.162
R2329 VDD.n1198 VDD.t20 9.162
R2330 VDD.n829 VDD.t19 9.162
R2331 VDD.n2572 VDD.t7 9.162
R2332 VDD.n2654 VDD.n2653 9.162
R2333 VDD.n2488 VDD.t8 9.162
R2334 VDD.n1011 VDD.t35 9.162
R2335 VDD.n1281 VDD.n1280 9.162
R2336 VDD.n1080 VDD.t36 9.162
R2337 VDD.n245 VDD.n244 9.162
R2338 VDD.n245 VDD.t32 9.162
R2339 VDD.n458 VDD.t33 9.162
R2340 VDD.n1639 VDD.n1638 9.162
R2341 VDD.n2863 VDD.t11 9.162
R2342 VDD.n3751 VDD.t47 9.162
R2343 VDD.n3793 VDD.t56 9.162
R2344 VDD.n3904 VDD.t52 9.162
R2345 VDD.n3852 VDD.t64 9.162
R2346 VDD.n4015 VDD.t63 9.162
R2347 VDD.n3963 VDD.t66 9.162
R2348 VDD.n4126 VDD.t65 9.162
R2349 VDD.n4074 VDD.t44 9.162
R2350 VDD.n4237 VDD.t51 9.162
R2351 VDD.n4185 VDD.t61 9.162
R2352 VDD.n4353 VDD.t58 9.162
R2353 VDD.n4395 VDD.t62 9.162
R2354 VDD.n4513 VDD.t49 9.162
R2355 VDD.n4461 VDD.t42 9.162
R2356 VDD.n4631 VDD.t54 9.162
R2357 VDD.n4579 VDD.t45 9.162
R2358 VDD.n4684 VDD.t57 9.162
R2359 VDD.n21 VDD.t60 9.162
R2360 VDD.n2841 VDD.n2840 9.02
R2361 VDD.n830 VDD.n829 9.02
R2362 VDD.n2573 VDD.n2572 9.02
R2363 VDD.n1012 VDD.n1011 9.02
R2364 VDD.n246 VDD.n245 9.02
R2365 VDD.n2489 VDD.n2488 9.018
R2366 VDD.n2655 VDD.n2654 9.018
R2367 VDD.n1081 VDD.n1080 9.018
R2368 VDD.n1282 VDD.n1281 9.018
R2369 VDD.n2193 VDD.n2192 9.018
R2370 VDD.n459 VDD.n458 9.018
R2371 VDD.n1640 VDD.n1639 9.018
R2372 VDD.n1199 VDD.n1198 9.018
R2373 VDD.n2753 VDD.n2752 9.018
R2374 VDD.n2864 VDD.n2863 9.018
R2375 VDD.n2765 VDD.n2758 9
R2376 VDD.n2808 VDD.n2756 9
R2377 VDD.n2785 VDD.n2784 9
R2378 VDD.n2775 VDD.n2757 9
R2379 VDD.n755 VDD.n748 9
R2380 VDD.n798 VDD.n746 9
R2381 VDD.n775 VDD.n774 9
R2382 VDD.n765 VDD.n747 9
R2383 VDD.n2541 VDD.n2540 9
R2384 VDD.n2498 VDD.n2494 9
R2385 VDD.n2508 VDD.n2493 9
R2386 VDD.n2517 VDD.n2492 9
R2387 VDD.n2476 VDD.n2422 9
R2388 VDD.n2467 VDD.n2423 9
R2389 VDD.n2487 VDD.n2486 9
R2390 VDD.n2457 VDD.n2424 9
R2391 VDD.n2652 VDD.n2575 9
R2392 VDD.n2628 VDD.n2576 9
R2393 VDD.n2619 VDD.n2577 9
R2394 VDD.n2609 VDD.n2578 9
R2395 VDD.n937 VDD.n933 9
R2396 VDD.n980 VDD.n931 9
R2397 VDD.n957 VDD.n956 9
R2398 VDD.n947 VDD.n932 9
R2399 VDD.n1049 VDD.n1016 9
R2400 VDD.n1068 VDD.n1014 9
R2401 VDD.n1079 VDD.n1078 9
R2402 VDD.n1059 VDD.n1015 9
R2403 VDD.n1310 VDD.n1309 9
R2404 VDD.n1320 VDD.n1319 9
R2405 VDD.n1299 VDD.n1298 9
R2406 VDD.n1331 VDD.n1330 9
R2407 VDD.n170 VDD.n163 9
R2408 VDD.n213 VDD.n161 9
R2409 VDD.n190 VDD.n189 9
R2410 VDD.n180 VDD.n162 9
R2411 VDD.n2180 VDD.n2179 9
R2412 VDD.n2170 VDD.n1914 9
R2413 VDD.n2191 VDD.n2190 9
R2414 VDD.n2160 VDD.n1915 9
R2415 VDD.n508 VDD.n507 9
R2416 VDD.n487 VDD.n486 9
R2417 VDD.n476 VDD.n475 9
R2418 VDD.n497 VDD.n496 9
R2419 VDD.n1668 VDD.n1667 9
R2420 VDD.n1678 VDD.n1677 9
R2421 VDD.n1657 VDD.n1656 9
R2422 VDD.n1689 VDD.n1688 9
R2423 VDD.n1234 VDD.n1233 9
R2424 VDD.n1213 VDD.n1212 9
R2425 VDD.n1202 VDD.n1201 9
R2426 VDD.n1223 VDD.n1222 9
R2427 VDD.n2740 VDD.n2739 9
R2428 VDD.n2730 VDD.n2679 9
R2429 VDD.n2751 VDD.n2750 9
R2430 VDD.n2720 VDD.n2680 9
R2431 VDD.n2913 VDD.n2912 9
R2432 VDD.n2892 VDD.n2891 9
R2433 VDD.n2881 VDD.n2880 9
R2434 VDD.n2902 VDD.n2901 9
R2435 VDD.n3787 VDD.n3786 9
R2436 VDD.n3808 VDD.n3792 9
R2437 VDD.n3745 VDD.n3744 9
R2438 VDD.n3766 VDD.n3750 9
R2439 VDD.n3733 VDD.n3732 9
R2440 VDD.n3775 VDD.n3774 9
R2441 VDD.n3867 VDD.n3851 9
R2442 VDD.n3898 VDD.n3897 9
R2443 VDD.n3919 VDD.n3903 9
R2444 VDD.n3846 VDD.n3845 9
R2445 VDD.n3834 VDD.n3833 9
R2446 VDD.n3886 VDD.n3885 9
R2447 VDD.n3978 VDD.n3962 9
R2448 VDD.n4009 VDD.n4008 9
R2449 VDD.n4030 VDD.n4014 9
R2450 VDD.n3957 VDD.n3956 9
R2451 VDD.n3945 VDD.n3944 9
R2452 VDD.n3997 VDD.n3996 9
R2453 VDD.n4089 VDD.n4073 9
R2454 VDD.n4120 VDD.n4119 9
R2455 VDD.n4141 VDD.n4125 9
R2456 VDD.n4068 VDD.n4067 9
R2457 VDD.n4056 VDD.n4055 9
R2458 VDD.n4108 VDD.n4107 9
R2459 VDD.n4200 VDD.n4184 9
R2460 VDD.n4231 VDD.n4230 9
R2461 VDD.n4252 VDD.n4236 9
R2462 VDD.n4179 VDD.n4178 9
R2463 VDD.n4167 VDD.n4166 9
R2464 VDD.n4219 VDD.n4218 9
R2465 VDD.n4389 VDD.n4388 9
R2466 VDD.n4410 VDD.n4394 9
R2467 VDD.n4347 VDD.n4346 9
R2468 VDD.n4368 VDD.n4352 9
R2469 VDD.n4335 VDD.n4334 9
R2470 VDD.n4377 VDD.n4376 9
R2471 VDD.n4476 VDD.n4460 9
R2472 VDD.n4507 VDD.n4506 9
R2473 VDD.n4528 VDD.n4512 9
R2474 VDD.n4455 VDD.n4454 9
R2475 VDD.n4443 VDD.n4442 9
R2476 VDD.n4495 VDD.n4494 9
R2477 VDD.n4594 VDD.n4578 9
R2478 VDD.n4625 VDD.n4624 9
R2479 VDD.n4646 VDD.n4630 9
R2480 VDD.n4573 VDD.n4572 9
R2481 VDD.n4561 VDD.n4560 9
R2482 VDD.n4613 VDD.n4612 9
R2483 VDD.n36 VDD.n20 9
R2484 VDD.n4678 VDD.n4677 9
R2485 VDD.n4699 VDD.n4683 9
R2486 VDD.n15 VDD.n14 9
R2487 VDD.n3 VDD.n2 9
R2488 VDD.n4666 VDD.n4665 9
R2489 VDD.n342 VDD.n341 8.855
R2490 VDD.n656 VDD.n655 8.855
R2491 VDD.n2019 VDD.n2018 8.855
R2492 VDD.n2015 VDD.n2014 8.855
R2493 VDD.n2012 VDD.n2011 8.855
R2494 VDD.n2356 VDD.n2355 8.855
R2495 VDD.n422 VDD.n421 8.855
R2496 VDD.n419 VDD.n418 8.855
R2497 VDD.n417 VDD.n416 8.855
R2498 VDD.n428 VDD.n427 8.855
R2499 VDD.n653 VDD.n652 8.855
R2500 VDD.n414 VDD.n413 8.855
R2501 VDD.n2022 VDD.n2021 8.855
R2502 VDD.n1905 VDD.n1904 8.855
R2503 VDD.n1904 VDD.n1903 8.855
R2504 VDD.n297 VDD.n296 8.855
R2505 VDD.n283 VDD.n282 8.855
R2506 VDD.n285 VDD.n284 8.855
R2507 VDD.n281 VDD.n280 8.855
R2508 VDD.n335 VDD.n281 8.855
R2509 VDD.n3583 VDD.n336 8.855
R2510 VDD.n336 VDD.n335 8.855
R2511 VDD.n704 VDD.n703 8.855
R2512 VDD.n690 VDD.n689 8.855
R2513 VDD.n692 VDD.n691 8.855
R2514 VDD.n688 VDD.n687 8.855
R2515 VDD.n742 VDD.n688 8.855
R2516 VDD.n2226 VDD.n743 8.855
R2517 VDD.n743 VDD.n742 8.855
R2518 VDD.n1279 VDD.n1278 8.855
R2519 VDD.n1123 VDD.n1122 8.855
R2520 VDD.n1128 VDD.n1127 8.855
R2521 VDD.n1126 VDD.n1125 8.855
R2522 VDD.n1168 VDD.n1167 8.855
R2523 VDD.n1167 VDD.n1166 8.855
R2524 VDD.n1120 VDD.n1119 8.855
R2525 VDD.n1834 VDD.n1833 8.855
R2526 VDD.n1461 VDD.n1460 8.855
R2527 VDD.n928 VDD.n927 8.855
R2528 VDD.n1632 VDD.n1631 8.855
R2529 VDD.n1636 VDD.n1635 8.855
R2530 VDD.n1731 VDD.n1730 8.855
R2531 VDD.n1838 VDD.n1837 8.855
R2532 VDD.n1837 VDD.n1836 8.855
R2533 VDD.n1843 VDD.n1842 8.855
R2534 VDD.n1842 VDD.n1841 8.855
R2535 VDD.n1854 VDD.n1853 8.855
R2536 VDD.n1853 VDD.n1852 8.855
R2537 VDD.n1867 VDD.n1866 8.855
R2538 VDD.n1866 VDD.n1865 8.855
R2539 VDD.n1872 VDD.n1871 8.855
R2540 VDD.n1871 VDD.n1870 8.855
R2541 VDD.n1879 VDD.n1878 8.855
R2542 VDD.n1878 VDD.n1877 8.855
R2543 VDD.n1883 VDD.n1882 8.855
R2544 VDD.n1882 VDD.n1881 8.855
R2545 VDD.n1887 VDD.n1886 8.855
R2546 VDD.n1886 VDD.n1885 8.855
R2547 VDD.n1891 VDD.n1890 8.855
R2548 VDD.n1890 VDD.n1889 8.855
R2549 VDD.n1897 VDD.n1896 8.855
R2550 VDD.n1896 VDD.n1895 8.855
R2551 VDD.n2222 VDD.n2221 8.855
R2552 VDD.n2221 VDD.n2220 8.855
R2553 VDD.n2218 VDD.n2217 8.855
R2554 VDD.n2217 VDD.n2216 8.855
R2555 VDD.n2214 VDD.n2213 8.855
R2556 VDD.n2213 VDD.n2212 8.855
R2557 VDD.n2210 VDD.n2209 8.855
R2558 VDD.n2209 VDD.n2208 8.855
R2559 VDD.n2206 VDD.n2204 8.855
R2560 VDD.n2204 VDD.n2203 8.855
R2561 VDD.n2199 VDD.n2198 8.855
R2562 VDD.n2198 VDD.n2197 8.855
R2563 VDD.n1911 VDD.n1910 8.855
R2564 VDD.n1910 VDD.n1909 8.855
R2565 VDD.n3625 VDD.n3624 8.855
R2566 VDD.n3624 VDD.n3623 8.855
R2567 VDD.n3617 VDD.n3616 8.855
R2568 VDD.n3616 VDD.n3615 8.855
R2569 VDD.n3613 VDD.n3612 8.855
R2570 VDD.n3612 VDD.n3611 8.855
R2571 VDD.n3606 VDD.n3605 8.855
R2572 VDD.n3605 VDD.n3604 8.855
R2573 VDD.n3602 VDD.n3601 8.855
R2574 VDD.n3601 VDD.n3600 8.855
R2575 VDD.n3598 VDD.n3597 8.855
R2576 VDD.n3597 VDD.n3596 8.855
R2577 VDD.n3594 VDD.n3593 8.855
R2578 VDD.n3593 VDD.n3592 8.855
R2579 VDD.n3590 VDD.n3588 8.855
R2580 VDD.n3588 VDD.n3587 8.855
R2581 VDD.n255 VDD.n254 8.855
R2582 VDD.n254 VDD.n253 8.855
R2583 VDD.n2663 VDD.n2662 8.855
R2584 VDD.n2662 VDD.n2661 8.855
R2585 VDD.n2667 VDD.n2666 8.855
R2586 VDD.n2666 VDD.n2665 8.855
R2587 VDD.n2671 VDD.n2670 8.855
R2588 VDD.n2670 VDD.n2669 8.855
R2589 VDD.n3190 VDD.n3189 8.855
R2590 VDD.n3293 VDD.n3292 8.855
R2591 VDD.n3193 VDD.n3192 8.855
R2592 VDD.n2413 VDD.n2412 8.855
R2593 VDD.n1468 VDD.n1467 8.855
R2594 VDD.n1477 VDD.n1476 8.855
R2595 VDD.n1489 VDD.n1488 8.855
R2596 VDD.n1493 VDD.n1492 8.855
R2597 VDD.n1507 VDD.n1506 8.855
R2598 VDD.n1502 VDD.n1501 8.855
R2599 VDD.n1499 VDD.n1498 8.855
R2600 VDD.n1496 VDD.n1495 8.855
R2601 VDD.n661 VDD.n660 8.855
R2602 VDD.n2360 VDD.n2359 8.855
R2603 VDD.n2363 VDD.n2362 8.855
R2604 VDD.n2366 VDD.n2365 8.855
R2605 VDD.n2369 VDD.n2368 8.855
R2606 VDD.n2374 VDD.n2373 8.855
R2607 VDD.n2378 VDD.n2377 8.855
R2608 VDD.n2381 VDD.n2380 8.855
R2609 VDD.n2384 VDD.n2383 8.855
R2610 VDD.n2387 VDD.n2386 8.855
R2611 VDD.n2392 VDD.n2391 8.855
R2612 VDD.n2396 VDD.n2395 8.855
R2613 VDD.n2399 VDD.n2398 8.855
R2614 VDD.n2402 VDD.n2401 8.855
R2615 VDD.n2405 VDD.n2404 8.855
R2616 VDD.n2410 VDD.n2409 8.855
R2617 VDD.n3454 VDD.n3453 8.855
R2618 VDD.n3451 VDD.n3450 8.855
R2619 VDD.n3448 VDD.n3447 8.855
R2620 VDD.n3445 VDD.n3444 8.855
R2621 VDD.n3442 VDD.n3441 8.855
R2622 VDD.n3436 VDD.n3435 8.855
R2623 VDD.n3429 VDD.n3428 8.855
R2624 VDD.n3423 VDD.n3422 8.855
R2625 VDD.n3421 VDD.n3420 8.855
R2626 VDD.n1464 VDD.n1463 8.855
R2627 VDD.n3019 VDD.n3018 8.855
R2628 VDD.n3021 VDD.n3020 8.855
R2629 VDD.n3061 VDD.n3060 8.855
R2630 VDD.n3060 VDD.n3059 8.855
R2631 VDD.n3014 VDD.n3013 8.855
R2632 VDD.n3417 VDD.n3416 8.855
R2633 VDD.n3017 VDD.n3016 8.855
R2634 VDD.n3059 VDD.n3017 8.855
R2635 VDD.n2659 VDD.n2658 8.855
R2636 VDD.n3089 VDD.n3088 8.855
R2637 VDD.n3088 VDD.n3087 8.855
R2638 VDD.n2677 VDD.n2676 8.855
R2639 VDD.n2676 VDD.n2675 8.855
R2640 VDD.n3082 VDD.n3081 8.855
R2641 VDD.n3081 VDD.n3080 8.855
R2642 VDD.n3074 VDD.n3073 8.855
R2643 VDD.n3073 VDD.n3072 8.855
R2644 VDD.n3067 VDD.n2852 8.855
R2645 VDD.n2852 VDD.n2851 8.855
R2646 VDD.n3066 VDD.n3065 8.855
R2647 VDD.n3065 VDD.n3064 8.855
R2648 VDD.n3305 VDD.n3304 8.764
R2649 VDD.n3426 VDD.n3425 8.764
R2650 VDD.n1619 VDD.n1618 8.764
R2651 VDD.n1480 VDD.n1479 8.764
R2652 VDD.n165 VDD.n164 8.764
R2653 VDD.n249 VDD.n248 8.764
R2654 VDD.n1857 VDD.n1856 8.764
R2655 VDD.n750 VDD.n749 8.764
R2656 VDD.n2760 VDD.n2759 8.764
R2657 VDD.n3070 VDD.n3069 8.764
R2658 VDD.n335 VDD.n325 8.762
R2659 VDD.n742 VDD.n732 8.762
R2660 VDD.n425 VDD.n384 8.762
R2661 VDD.n425 VDD.n374 8.762
R2662 VDD.n1166 VDD.n1156 8.762
R2663 VDD.n3059 VDD.n3049 8.762
R2664 VDD.n298 VDD.n295 8.663
R2665 VDD.n705 VDD.n702 8.663
R2666 VDD.n415 VDD.n412 8.662
R2667 VDD.n335 VDD.n269 8.581
R2668 VDD.n742 VDD.n675 8.581
R2669 VDD.n1166 VDD.n1096 8.581
R2670 VDD.n3059 VDD.n2992 8.581
R2671 VDD.n426 VDD.n346 8.448
R2672 VDD.n335 VDD.n334 8.408
R2673 VDD.n742 VDD.n741 8.408
R2674 VDD.n425 VDD.n403 8.408
R2675 VDD.n425 VDD.n355 8.408
R2676 VDD.n1166 VDD.n1165 8.408
R2677 VDD.n3059 VDD.n3058 8.408
R2678 VDD.n3022 VDD.n3019 8.381
R2679 VDD.n1129 VDD.n1128 8.361
R2680 VDD.n1129 VDD.n1126 8.361
R2681 VDD.n3613 VDD.n3609 8.282
R2682 VDD.n2392 VDD.n2389 8.282
R2683 VDD.n415 VDD.n414 8.247
R2684 VDD.n298 VDD.n297 8.247
R2685 VDD.n705 VDD.n704 8.247
R2686 VDD.n335 VDD.n260 8.241
R2687 VDD.n742 VDD.n666 8.241
R2688 VDD.n1166 VDD.n1087 8.241
R2689 VDD.n3059 VDD.n2983 8.241
R2690 VDD.n427 VDD.n426 8.044
R2691 VDD.n423 VDD.n422 8.044
R2692 VDD.n1121 VDD.n1120 8.044
R2693 VDD.n1833 VDD.n1832 8.044
R2694 VDD.n3015 VDD.n3014 8.044
R2695 VDD.n286 VDD.n283 8
R2696 VDD.n693 VDD.n690 8
R2697 VDD.n420 VDD.n417 8
R2698 VDD.n420 VDD.n419 8
R2699 VDD.n286 VDD.n285 7.999
R2700 VDD.n693 VDD.n692 7.999
R2701 VDD.n3022 VDD.n3021 7.98
R2702 VDD.n3600 VDD.t48 7.653
R2703 VDD.n2665 VDD.t55 7.653
R2704 VDD.n3753 VDD.n3752 7.474
R2705 VDD.n3795 VDD.n3794 7.474
R2706 VDD.n3906 VDD.n3905 7.474
R2707 VDD.n3854 VDD.n3853 7.474
R2708 VDD.n4017 VDD.n4016 7.474
R2709 VDD.n3965 VDD.n3964 7.474
R2710 VDD.n4128 VDD.n4127 7.474
R2711 VDD.n4076 VDD.n4075 7.474
R2712 VDD.n4239 VDD.n4238 7.474
R2713 VDD.n4187 VDD.n4186 7.474
R2714 VDD.n4355 VDD.n4354 7.474
R2715 VDD.n4397 VDD.n4396 7.474
R2716 VDD.n4515 VDD.n4514 7.474
R2717 VDD.n4463 VDD.n4462 7.474
R2718 VDD.n4633 VDD.n4632 7.474
R2719 VDD.n4581 VDD.n4580 7.474
R2720 VDD.n4686 VDD.n4685 7.474
R2721 VDD.n23 VDD.n22 7.474
R2722 VDD.n3156 VDD.n3155 6.206
R2723 VDD.n3229 VDD.n3228 6.206
R2724 VDD.n684 VDD.n678 6.206
R2725 VDD.n2325 VDD.n2324 6.206
R2726 VDD.n2088 VDD.n2087 6.206
R2727 VDD.n1948 VDD.n1947 6.206
R2728 VDD.n278 VDD.n272 6.206
R2729 VDD.n3491 VDD.n3490 6.206
R2730 VDD.n364 VDD.n358 6.206
R2731 VDD.n393 VDD.n387 6.206
R2732 VDD.n587 VDD.n585 6.206
R2733 VDD.n621 VDD.n619 6.206
R2734 VDD.n1105 VDD.n1099 6.206
R2735 VDD.n1577 VDD.n1576 6.206
R2736 VDD.n1544 VDD.n1543 6.206
R2737 VDD.n3001 VDD.n2995 6.206
R2738 VDD.n3351 VDD.n3349 6.206
R2739 VDD.n3385 VDD.n3383 6.206
R2740 VDD.n1766 VDD.n1765 6.206
R2741 VDD.n1429 VDD.n1428 6.206
R2742 VDD.n725 VDD.n724 6.023
R2743 VDD.n727 VDD.n726 6.023
R2744 VDD.n719 VDD.n718 6.023
R2745 VDD.n721 VDD.n720 6.023
R2746 VDD.n2301 VDD.n2300 6.023
R2747 VDD.n2309 VDD.n2308 6.023
R2748 VDD.n2064 VDD.n2063 6.023
R2749 VDD.n2072 VDD.n2071 6.023
R2750 VDD.n1964 VDD.n1963 6.023
R2751 VDD.n1956 VDD.n1955 6.023
R2752 VDD.n318 VDD.n317 6.023
R2753 VDD.n320 VDD.n319 6.023
R2754 VDD.n312 VDD.n311 6.023
R2755 VDD.n314 VDD.n313 6.023
R2756 VDD.n3507 VDD.n3506 6.023
R2757 VDD.n3499 VDD.n3498 6.023
R2758 VDD.n367 VDD.n366 6.023
R2759 VDD.n369 VDD.n368 6.023
R2760 VDD.n379 VDD.n378 6.023
R2761 VDD.n381 VDD.n380 6.023
R2762 VDD.n595 VDD.n594 6.023
R2763 VDD.n603 VDD.n602 6.023
R2764 VDD.n1149 VDD.n1148 6.023
R2765 VDD.n1151 VDD.n1150 6.023
R2766 VDD.n1143 VDD.n1142 6.023
R2767 VDD.n1145 VDD.n1144 6.023
R2768 VDD.n1561 VDD.n1560 6.023
R2769 VDD.n1552 VDD.n1551 6.023
R2770 VDD.n1782 VDD.n1781 6.023
R2771 VDD.n1774 VDD.n1773 6.023
R2772 VDD.n1405 VDD.n1404 6.023
R2773 VDD.n1413 VDD.n1412 6.023
R2774 VDD.n3590 VDD.n3589 6.023
R2775 VDD.n3132 VDD.n3131 6.023
R2776 VDD.n3140 VDD.n3139 6.023
R2777 VDD.n3245 VDD.n3244 6.023
R2778 VDD.n3237 VDD.n3236 6.023
R2779 VDD.n2410 VDD.n2407 6.023
R2780 VDD.n3042 VDD.n3041 6.023
R2781 VDD.n3044 VDD.n3043 6.023
R2782 VDD.n3036 VDD.n3035 6.023
R2783 VDD.n3038 VDD.n3037 6.023
R2784 VDD.n3359 VDD.n3358 6.023
R2785 VDD.n3367 VDD.n3366 6.023
R2786 VDD.n3123 VDD.n3122 5.727
R2787 VDD.n3260 VDD.n3259 5.727
R2788 VDD.n675 VDD.n674 5.727
R2789 VDD.n2292 VDD.n2291 5.727
R2790 VDD.n2055 VDD.n2054 5.727
R2791 VDD.n1979 VDD.n1978 5.727
R2792 VDD.n269 VDD.n268 5.727
R2793 VDD.n3522 VDD.n3521 5.727
R2794 VDD.n1096 VDD.n1095 5.727
R2795 VDD.n2992 VDD.n2991 5.727
R2796 VDD.n1797 VDD.n1796 5.727
R2797 VDD.n1396 VDD.n1395 5.727
R2798 VDD.n1903 VDD.n1900 5.661
R2799 VDD.n742 VDD.n685 5.661
R2800 VDD.n425 VDD.n394 5.661
R2801 VDD.n425 VDD.n365 5.661
R2802 VDD.n1166 VDD.n1116 5.661
R2803 VDD.n1166 VDD.n1117 5.661
R2804 VDD.n668 VDD.n667 5.27
R2805 VDD.n670 VDD.n669 5.27
R2806 VDD.n680 VDD.n679 5.27
R2807 VDD.n682 VDD.n681 5.27
R2808 VDD.n2289 VDD.n2288 5.27
R2809 VDD.n2321 VDD.n2320 5.27
R2810 VDD.n2052 VDD.n2051 5.27
R2811 VDD.n2084 VDD.n2083 5.27
R2812 VDD.n1976 VDD.n1975 5.27
R2813 VDD.n1944 VDD.n1943 5.27
R2814 VDD.n262 VDD.n261 5.27
R2815 VDD.n264 VDD.n263 5.27
R2816 VDD.n274 VDD.n273 5.27
R2817 VDD.n276 VDD.n275 5.27
R2818 VDD.n3519 VDD.n3518 5.27
R2819 VDD.n3487 VDD.n3486 5.27
R2820 VDD.n360 VDD.n359 5.27
R2821 VDD.n362 VDD.n361 5.27
R2822 VDD.n389 VDD.n388 5.27
R2823 VDD.n391 VDD.n390 5.27
R2824 VDD.n582 VDD.n581 5.27
R2825 VDD.n616 VDD.n615 5.27
R2826 VDD.n1089 VDD.n1088 5.27
R2827 VDD.n1091 VDD.n1090 5.27
R2828 VDD.n1101 VDD.n1100 5.27
R2829 VDD.n1103 VDD.n1102 5.27
R2830 VDD.n1573 VDD.n1572 5.27
R2831 VDD.n1540 VDD.n1539 5.27
R2832 VDD.n1794 VDD.n1793 5.27
R2833 VDD.n1762 VDD.n1761 5.27
R2834 VDD.n1393 VDD.n1392 5.27
R2835 VDD.n1425 VDD.n1424 5.27
R2836 VDD.n3120 VDD.n3119 5.27
R2837 VDD.n3152 VDD.n3151 5.27
R2838 VDD.n3257 VDD.n3256 5.27
R2839 VDD.n3225 VDD.n3224 5.27
R2840 VDD.n2985 VDD.n2984 5.27
R2841 VDD.n2987 VDD.n2986 5.27
R2842 VDD.n2997 VDD.n2996 5.27
R2843 VDD.n2999 VDD.n2998 5.27
R2844 VDD.n3346 VDD.n3345 5.27
R2845 VDD.n3380 VDD.n3379 5.27
R2846 VDD.n1115 VDD.n1114 5.198
R2847 VDD.n3011 VDD.n3010 5.198
R2848 VDD.n2661 VDD.t46 4.783
R2849 VDD.n2851 VDD.t6 4.783
R2850 VDD.n3306 VDD.n3305 4.65
R2851 VDD.n3427 VDD.n3426 4.65
R2852 VDD.n1620 VDD.n1619 4.65
R2853 VDD.n1481 VDD.n1480 4.65
R2854 VDD.n657 VDD.n656 4.65
R2855 VDD.n2020 VDD.n2019 4.65
R2856 VDD.n2016 VDD.n2015 4.65
R2857 VDD.n2013 VDD.n2012 4.65
R2858 VDD.n428 VDD.n252 4.65
R2859 VDD.n654 VDD.n653 4.65
R2860 VDD.n166 VDD.n165 4.65
R2861 VDD.n2119 VDD.n2022 4.65
R2862 VDD.n1906 VDD.n1905 4.65
R2863 VDD.n250 VDD.n249 4.65
R2864 VDD.n3584 VDD.n3583 4.65
R2865 VDD.n3457 VDD.n342 4.65
R2866 VDD.n2226 VDD.n2225 4.65
R2867 VDD.n2357 VDD.n2356 4.65
R2868 VDD.n1858 VDD.n1857 4.65
R2869 VDD.n751 VDD.n750 4.65
R2870 VDD.n1510 VDD.n1279 4.65
R2871 VDD.n1168 VDD.n744 4.65
R2872 VDD.n1462 VDD.n1461 4.65
R2873 VDD.n929 VDD.n928 4.65
R2874 VDD.n1633 VDD.n1632 4.65
R2875 VDD.n1637 VDD.n1636 4.65
R2876 VDD.n1732 VDD.n1731 4.65
R2877 VDD.n1835 VDD.n1834 4.65
R2878 VDD.n1839 VDD.n1838 4.65
R2879 VDD.n1844 VDD.n1843 4.65
R2880 VDD.n1855 VDD.n1854 4.65
R2881 VDD.n1868 VDD.n1867 4.65
R2882 VDD.n1873 VDD.n1872 4.65
R2883 VDD.n1880 VDD.n1879 4.65
R2884 VDD.n1884 VDD.n1883 4.65
R2885 VDD.n1888 VDD.n1887 4.65
R2886 VDD.n1892 VDD.n1891 4.65
R2887 VDD.n1898 VDD.n1897 4.65
R2888 VDD.n2223 VDD.n2222 4.65
R2889 VDD.n2219 VDD.n2218 4.65
R2890 VDD.n2215 VDD.n2214 4.65
R2891 VDD.n2211 VDD.n2210 4.65
R2892 VDD.n2207 VDD.n2206 4.65
R2893 VDD.n2200 VDD.n2199 4.65
R2894 VDD.n1912 VDD.n1911 4.65
R2895 VDD.n3626 VDD.n3625 4.65
R2896 VDD.n3618 VDD.n3617 4.65
R2897 VDD.n3614 VDD.n3613 4.65
R2898 VDD.n3607 VDD.n3606 4.65
R2899 VDD.n3603 VDD.n3602 4.65
R2900 VDD.n3599 VDD.n3598 4.65
R2901 VDD.n3595 VDD.n3594 4.65
R2902 VDD.n3591 VDD.n3590 4.65
R2903 VDD.n256 VDD.n255 4.65
R2904 VDD.n2664 VDD.n2663 4.65
R2905 VDD.n2668 VDD.n2667 4.65
R2906 VDD.n2672 VDD.n2671 4.65
R2907 VDD.n3191 VDD.n3190 4.65
R2908 VDD.n3294 VDD.n3293 4.65
R2909 VDD.n3194 VDD.n3193 4.65
R2910 VDD.n2414 VDD.n2413 4.65
R2911 VDD.n1469 VDD.n1468 4.65
R2912 VDD.n1478 VDD.n1477 4.65
R2913 VDD.n1490 VDD.n1489 4.65
R2914 VDD.n1494 VDD.n1493 4.65
R2915 VDD.n1508 VDD.n1507 4.65
R2916 VDD.n1503 VDD.n1502 4.65
R2917 VDD.n1500 VDD.n1499 4.65
R2918 VDD.n1497 VDD.n1496 4.65
R2919 VDD.n662 VDD.n661 4.65
R2920 VDD.n2361 VDD.n2360 4.65
R2921 VDD.n2364 VDD.n2363 4.65
R2922 VDD.n2367 VDD.n2366 4.65
R2923 VDD.n2370 VDD.n2369 4.65
R2924 VDD.n2375 VDD.n2374 4.65
R2925 VDD.n2379 VDD.n2378 4.65
R2926 VDD.n2382 VDD.n2381 4.65
R2927 VDD.n2385 VDD.n2384 4.65
R2928 VDD.n2388 VDD.n2387 4.65
R2929 VDD.n2393 VDD.n2392 4.65
R2930 VDD.n2397 VDD.n2396 4.65
R2931 VDD.n2400 VDD.n2399 4.65
R2932 VDD.n2403 VDD.n2402 4.65
R2933 VDD.n2406 VDD.n2405 4.65
R2934 VDD.n2411 VDD.n2410 4.65
R2935 VDD.n3455 VDD.n3454 4.65
R2936 VDD.n3452 VDD.n3451 4.65
R2937 VDD.n3449 VDD.n3448 4.65
R2938 VDD.n3446 VDD.n3445 4.65
R2939 VDD.n3443 VDD.n3442 4.65
R2940 VDD.n3437 VDD.n3436 4.65
R2941 VDD.n3430 VDD.n3429 4.65
R2942 VDD.n3424 VDD.n3423 4.65
R2943 VDD.n3421 VDD.n3419 4.65
R2944 VDD.n1465 VDD.n1464 4.65
R2945 VDD.n3062 VDD.n3061 4.65
R2946 VDD.n3418 VDD.n3417 4.65
R2947 VDD.n2761 VDD.n2760 4.65
R2948 VDD.n3187 VDD.n2659 4.65
R2949 VDD.n3090 VDD.n3089 4.65
R2950 VDD.n3071 VDD.n3070 4.65
R2951 VDD.n2678 VDD.n2677 4.65
R2952 VDD.n3083 VDD.n3082 4.65
R2953 VDD.n3075 VDD.n3074 4.65
R2954 VDD.n3068 VDD.n3067 4.65
R2955 VDD.n3066 VDD.n3063 4.65
R2956 VDD.n3078 VDD.n3077 4.589
R2957 VDD.n2860 VDD.n2859 4.589
R2958 VDD.n3433 VDD.n3432 4.589
R2959 VDD.n2419 VDD.n2418 4.589
R2960 VDD.n1913 VDD.n1908 4.589
R2961 VDD.n3622 VDD.n3621 4.589
R2962 VDD.n1166 VDD.n1124 4.559
R2963 VDD.n734 VDD.n733 4.517
R2964 VDD.n736 VDD.n735 4.517
R2965 VDD.n710 VDD.n709 4.517
R2966 VDD.n712 VDD.n711 4.517
R2967 VDD.n2277 VDD.n2276 4.517
R2968 VDD.n2333 VDD.n2332 4.517
R2969 VDD.n2040 VDD.n2039 4.517
R2970 VDD.n2096 VDD.n2095 4.517
R2971 VDD.n1988 VDD.n1987 4.517
R2972 VDD.n1932 VDD.n1931 4.517
R2973 VDD.n327 VDD.n326 4.517
R2974 VDD.n329 VDD.n328 4.517
R2975 VDD.n303 VDD.n302 4.517
R2976 VDD.n305 VDD.n304 4.517
R2977 VDD.n3531 VDD.n3530 4.517
R2978 VDD.n3474 VDD.n3473 4.517
R2979 VDD.n348 VDD.n347 4.517
R2980 VDD.n350 VDD.n349 4.517
R2981 VDD.n398 VDD.n397 4.517
R2982 VDD.n400 VDD.n399 4.517
R2983 VDD.n570 VDD.n569 4.517
R2984 VDD.n629 VDD.n628 4.517
R2985 VDD.n1158 VDD.n1157 4.517
R2986 VDD.n1160 VDD.n1159 4.517
R2987 VDD.n1134 VDD.n1133 4.517
R2988 VDD.n1136 VDD.n1135 4.517
R2989 VDD.n1585 VDD.n1584 4.517
R2990 VDD.n1528 VDD.n1527 4.517
R2991 VDD.n1806 VDD.n1805 4.517
R2992 VDD.n1750 VDD.n1749 4.517
R2993 VDD.n1381 VDD.n1380 4.517
R2994 VDD.n1437 VDD.n1436 4.517
R2995 VDD.n3108 VDD.n3107 4.517
R2996 VDD.n3164 VDD.n3163 4.517
R2997 VDD.n3269 VDD.n3268 4.517
R2998 VDD.n3212 VDD.n3211 4.517
R2999 VDD.n3051 VDD.n3050 4.517
R3000 VDD.n3053 VDD.n3052 4.517
R3001 VDD.n3027 VDD.n3026 4.517
R3002 VDD.n3029 VDD.n3028 4.517
R3003 VDD.n3334 VDD.n3333 4.517
R3004 VDD.n3393 VDD.n3392 4.517
R3005 VDD.n1635 VDD.n1634 4.279
R3006 VDD.n1631 VDD.n1630 4.279
R3007 VDD.n3189 VDD.n3188 4.079
R3008 VDD.n2018 VDD.n2017 4.079
R3009 VDD.n1124 VDD.n1123 4.079
R3010 VDD.n927 VDD.n926 4.079
R3011 VDD.n1166 VDD.n1115 3.906
R3012 VDD.n3059 VDD.n3011 3.906
R3013 VDD.n2231 VDD.n2230 3.764
R3014 VDD.n2228 VDD.n2227 3.764
R3015 VDD.n698 VDD.n697 3.764
R3016 VDD.n700 VDD.n699 3.764
R3017 VDD.n2265 VDD.n2264 3.764
R3018 VDD.n2345 VDD.n2344 3.764
R3019 VDD.n2028 VDD.n2027 3.764
R3020 VDD.n2108 VDD.n2107 3.764
R3021 VDD.n2000 VDD.n1999 3.764
R3022 VDD.n1921 VDD.n1920 3.764
R3023 VDD.n3582 VDD.n340 3.764
R3024 VDD.n338 VDD.n337 3.764
R3025 VDD.n291 VDD.n290 3.764
R3026 VDD.n293 VDD.n292 3.764
R3027 VDD.n3543 VDD.n3542 3.764
R3028 VDD.n3463 VDD.n3462 3.764
R3029 VDD.n433 VDD.n432 3.764
R3030 VDD.n430 VDD.n429 3.764
R3031 VDD.n408 VDD.n407 3.764
R3032 VDD.n410 VDD.n409 3.764
R3033 VDD.n558 VDD.n557 3.764
R3034 VDD.n641 VDD.n640 3.764
R3035 VDD.n1173 VDD.n1172 3.764
R3036 VDD.n1170 VDD.n1169 3.764
R3037 VDD.n1110 VDD.n1109 3.764
R3038 VDD.n1112 VDD.n1111 3.764
R3039 VDD.n1597 VDD.n1596 3.764
R3040 VDD.n1516 VDD.n1515 3.764
R3041 VDD.n1818 VDD.n1817 3.764
R3042 VDD.n1738 VDD.n1737 3.764
R3043 VDD.n1369 VDD.n1368 3.764
R3044 VDD.n1449 VDD.n1448 3.764
R3045 VDD.n2677 VDD.n2673 3.764
R3046 VDD.n3096 VDD.n3095 3.764
R3047 VDD.n3176 VDD.n3175 3.764
R3048 VDD.n3281 VDD.n3280 3.764
R3049 VDD.n3200 VDD.n3199 3.764
R3050 VDD.n3442 VDD.n3439 3.764
R3051 VDD.n2979 VDD.n2856 3.764
R3052 VDD.n2854 VDD.n2853 3.764
R3053 VDD.n3006 VDD.n3005 3.764
R3054 VDD.n3008 VDD.n3007 3.764
R3055 VDD.n3322 VDD.n3321 3.764
R3056 VDD.n3405 VDD.n3404 3.764
R3057 VDD.n3753 VDD.n3751 3.575
R3058 VDD.n3795 VDD.n3793 3.575
R3059 VDD.n3906 VDD.n3904 3.575
R3060 VDD.n3854 VDD.n3852 3.575
R3061 VDD.n4017 VDD.n4015 3.575
R3062 VDD.n3965 VDD.n3963 3.575
R3063 VDD.n4128 VDD.n4126 3.575
R3064 VDD.n4076 VDD.n4074 3.575
R3065 VDD.n4239 VDD.n4237 3.575
R3066 VDD.n4187 VDD.n4185 3.575
R3067 VDD.n4355 VDD.n4353 3.575
R3068 VDD.n4397 VDD.n4395 3.575
R3069 VDD.n4515 VDD.n4513 3.575
R3070 VDD.n4463 VDD.n4461 3.575
R3071 VDD.n4633 VDD.n4631 3.575
R3072 VDD.n4581 VDD.n4579 3.575
R3073 VDD.n4686 VDD.n4684 3.575
R3074 VDD.n23 VDD.n21 3.575
R3075 VDD.n394 VDD.n393 3.356
R3076 VDD.n621 VDD.n620 3.356
R3077 VDD.n365 VDD.n364 3.356
R3078 VDD.n587 VDD.n586 3.356
R3079 VDD.n3479 VDD.n3478 3.356
R3080 VDD.n3385 VDD.n3384 3.356
R3081 VDD.n3217 VDD.n3216 3.356
R3082 VDD.n3351 VDD.n3350 3.356
R3083 VDD.n2808 VDD.n2807 3.008
R3084 VDD.n798 VDD.n797 3.008
R3085 VDD.n2541 VDD.n2539 3.008
R3086 VDD.n980 VDD.n979 3.008
R3087 VDD.n213 VDD.n212 3.008
R3088 VDD.n2652 VDD.n2651 3
R3089 VDD.n1299 VDD.n1297 3
R3090 VDD.n476 VDD.n474 3
R3091 VDD.n1657 VDD.n1655 3
R3092 VDD.n2881 VDD.n2879 3
R3093 VDD.n2230 VDD.n2229 2.635
R3094 VDD.n2229 VDD.n2228 2.635
R3095 VDD.n701 VDD.n698 2.635
R3096 VDD.n701 VDD.n700 2.635
R3097 VDD.n2270 VDD.n2265 2.635
R3098 VDD.n2349 VDD.n2345 2.635
R3099 VDD.n2033 VDD.n2028 2.635
R3100 VDD.n2113 VDD.n2108 2.635
R3101 VDD.n2005 VDD.n2000 2.635
R3102 VDD.n1925 VDD.n1921 2.635
R3103 VDD.n340 VDD.n339 2.635
R3104 VDD.n339 VDD.n338 2.635
R3105 VDD.n294 VDD.n291 2.635
R3106 VDD.n294 VDD.n293 2.635
R3107 VDD.n3548 VDD.n3543 2.635
R3108 VDD.n3467 VDD.n3463 2.635
R3109 VDD.n432 VDD.n431 2.635
R3110 VDD.n431 VDD.n430 2.635
R3111 VDD.n411 VDD.n408 2.635
R3112 VDD.n411 VDD.n410 2.635
R3113 VDD.n563 VDD.n558 2.635
R3114 VDD.n646 VDD.n641 2.635
R3115 VDD.n1172 VDD.n1171 2.635
R3116 VDD.n1171 VDD.n1170 2.635
R3117 VDD.n1113 VDD.n1110 2.635
R3118 VDD.n1113 VDD.n1112 2.635
R3119 VDD.n1602 VDD.n1597 2.635
R3120 VDD.n1521 VDD.n1516 2.635
R3121 VDD.n1823 VDD.n1818 2.635
R3122 VDD.n1743 VDD.n1738 2.635
R3123 VDD.n1374 VDD.n1369 2.635
R3124 VDD.n1454 VDD.n1449 2.635
R3125 VDD.n3101 VDD.n3096 2.635
R3126 VDD.n3181 VDD.n3176 2.635
R3127 VDD.n3286 VDD.n3281 2.635
R3128 VDD.n3205 VDD.n3200 2.635
R3129 VDD.n2856 VDD.n2855 2.635
R3130 VDD.n2855 VDD.n2854 2.635
R3131 VDD.n3009 VDD.n3006 2.635
R3132 VDD.n3009 VDD.n3008 2.635
R3133 VDD.n3327 VDD.n3322 2.635
R3134 VDD.n3410 VDD.n3405 2.635
R3135 VDD.n3144 VDD.n3143 2.068
R3136 VDD.n3241 VDD.n3240 2.068
R3137 VDD.n723 VDD.n717 2.068
R3138 VDD.n2313 VDD.n2312 2.068
R3139 VDD.n2076 VDD.n2075 2.068
R3140 VDD.n1960 VDD.n1959 2.068
R3141 VDD.n316 VDD.n310 2.068
R3142 VDD.n3503 VDD.n3502 2.068
R3143 VDD.n1147 VDD.n1141 2.068
R3144 VDD.n3040 VDD.n3034 2.068
R3145 VDD.n1778 VDD.n1777 2.068
R3146 VDD.n1417 VDD.n1416 2.068
R3147 VDD.n3135 VDD.n3134 1.949
R3148 VDD.n3248 VDD.n3247 1.949
R3149 VDD.n732 VDD.n731 1.949
R3150 VDD.n2304 VDD.n2303 1.949
R3151 VDD.n2067 VDD.n2066 1.949
R3152 VDD.n1967 VDD.n1966 1.949
R3153 VDD.n325 VDD.n324 1.949
R3154 VDD.n3510 VDD.n3509 1.949
R3155 VDD.n384 VDD.n377 1.949
R3156 VDD.n607 VDD.n606 1.949
R3157 VDD.n598 VDD.n597 1.949
R3158 VDD.n374 VDD.n373 1.949
R3159 VDD.n1156 VDD.n1155 1.949
R3160 VDD.n1556 VDD.n1555 1.949
R3161 VDD.n1564 VDD.n1563 1.949
R3162 VDD.n3049 VDD.n3048 1.949
R3163 VDD.n3371 VDD.n3370 1.949
R3164 VDD.n1785 VDD.n1784 1.949
R3165 VDD.n1408 VDD.n1407 1.949
R3166 VDD.n3362 VDD.n3361 1.949
R3167 VDD.n4258 VDD.n4257 1.94
R3168 VDD.n4147 VDD.n4146 1.94
R3169 VDD.n4036 VDD.n4035 1.94
R3170 VDD.n3925 VDD.n3924 1.94
R3171 VDD.n3814 VDD.n3771 1.94
R3172 VDD.n3814 VDD.n3813 1.94
R3173 VDD.n4705 VDD.n4704 1.94
R3174 VDD.n4652 VDD.n4651 1.94
R3175 VDD.n4534 VDD.n4533 1.94
R3176 VDD.n4416 VDD.n4373 1.94
R3177 VDD.n4416 VDD.n4415 1.94
R3178 VDD.n3925 VDD.n3872 1.94
R3179 VDD.n4036 VDD.n3983 1.94
R3180 VDD.n4147 VDD.n4094 1.94
R3181 VDD.n4258 VDD.n4205 1.94
R3182 VDD.n4534 VDD.n4481 1.94
R3183 VDD.n4652 VDD.n4599 1.94
R3184 VDD.n4705 VDD.n41 1.94
R3185 VDD.n3072 VDD.t1 1.913
R3186 VDD.n737 VDD.n734 1.882
R3187 VDD.n737 VDD.n736 1.882
R3188 VDD.n713 VDD.n710 1.882
R3189 VDD.n713 VDD.n712 1.882
R3190 VDD.n2282 VDD.n2277 1.882
R3191 VDD.n2338 VDD.n2333 1.882
R3192 VDD.n2045 VDD.n2040 1.882
R3193 VDD.n2101 VDD.n2096 1.882
R3194 VDD.n1993 VDD.n1988 1.882
R3195 VDD.n1937 VDD.n1932 1.882
R3196 VDD.n330 VDD.n327 1.882
R3197 VDD.n330 VDD.n329 1.882
R3198 VDD.n306 VDD.n303 1.882
R3199 VDD.n306 VDD.n305 1.882
R3200 VDD.n3536 VDD.n3531 1.882
R3201 VDD.n3480 VDD.n3474 1.882
R3202 VDD.n351 VDD.n348 1.882
R3203 VDD.n351 VDD.n350 1.882
R3204 VDD.n401 VDD.n398 1.882
R3205 VDD.n401 VDD.n400 1.882
R3206 VDD.n575 VDD.n570 1.882
R3207 VDD.n634 VDD.n629 1.882
R3208 VDD.n1161 VDD.n1158 1.882
R3209 VDD.n1161 VDD.n1160 1.882
R3210 VDD.n1137 VDD.n1134 1.882
R3211 VDD.n1137 VDD.n1136 1.882
R3212 VDD.n1590 VDD.n1585 1.882
R3213 VDD.n1533 VDD.n1528 1.882
R3214 VDD.n1811 VDD.n1806 1.882
R3215 VDD.n1755 VDD.n1750 1.882
R3216 VDD.n1386 VDD.n1381 1.882
R3217 VDD.n1442 VDD.n1437 1.882
R3218 VDD.n3113 VDD.n3108 1.882
R3219 VDD.n3169 VDD.n3164 1.882
R3220 VDD.n3274 VDD.n3269 1.882
R3221 VDD.n3218 VDD.n3212 1.882
R3222 VDD.n3054 VDD.n3051 1.882
R3223 VDD.n3054 VDD.n3053 1.882
R3224 VDD.n3030 VDD.n3027 1.882
R3225 VDD.n3030 VDD.n3029 1.882
R3226 VDD.n3339 VDD.n3334 1.882
R3227 VDD.n3398 VDD.n3393 1.882
R3228 VDD.n4260 VDD.n4259 1.135
R3229 VDD.n4267 VDD.n4148 1.135
R3230 VDD.n4274 VDD.n4037 1.135
R3231 VDD.n4281 VDD.n3926 1.135
R3232 VDD.n4288 VDD.n3815 1.135
R3233 VDD.n4662 VDD.n4661 1.135
R3234 VDD.n4654 VDD.n4653 1.135
R3235 VDD.n4536 VDD.n4535 1.135
R3236 VDD.n4418 VDD.n4417 1.135
R3237 VDD.n671 VDD.n668 1.129
R3238 VDD.n671 VDD.n670 1.129
R3239 VDD.n683 VDD.n680 1.129
R3240 VDD.n683 VDD.n682 1.129
R3241 VDD.n2294 VDD.n2289 1.129
R3242 VDD.n2326 VDD.n2321 1.129
R3243 VDD.n2057 VDD.n2052 1.129
R3244 VDD.n2089 VDD.n2084 1.129
R3245 VDD.n1981 VDD.n1976 1.129
R3246 VDD.n1949 VDD.n1944 1.129
R3247 VDD.n265 VDD.n262 1.129
R3248 VDD.n265 VDD.n264 1.129
R3249 VDD.n277 VDD.n274 1.129
R3250 VDD.n277 VDD.n276 1.129
R3251 VDD.n3524 VDD.n3519 1.129
R3252 VDD.n3492 VDD.n3487 1.129
R3253 VDD.n363 VDD.n360 1.129
R3254 VDD.n363 VDD.n362 1.129
R3255 VDD.n392 VDD.n389 1.129
R3256 VDD.n392 VDD.n391 1.129
R3257 VDD.n588 VDD.n582 1.129
R3258 VDD.n622 VDD.n616 1.129
R3259 VDD.n1092 VDD.n1089 1.129
R3260 VDD.n1092 VDD.n1091 1.129
R3261 VDD.n1104 VDD.n1101 1.129
R3262 VDD.n1104 VDD.n1103 1.129
R3263 VDD.n1578 VDD.n1573 1.129
R3264 VDD.n1545 VDD.n1540 1.129
R3265 VDD.n1799 VDD.n1794 1.129
R3266 VDD.n1767 VDD.n1762 1.129
R3267 VDD.n1398 VDD.n1393 1.129
R3268 VDD.n1430 VDD.n1425 1.129
R3269 VDD.n3125 VDD.n3120 1.129
R3270 VDD.n3157 VDD.n3152 1.129
R3271 VDD.n3262 VDD.n3257 1.129
R3272 VDD.n3230 VDD.n3225 1.129
R3273 VDD.n2988 VDD.n2985 1.129
R3274 VDD.n2988 VDD.n2987 1.129
R3275 VDD.n3000 VDD.n2997 1.129
R3276 VDD.n3000 VDD.n2999 1.129
R3277 VDD.n3352 VDD.n3346 1.129
R3278 VDD.n3386 VDD.n3380 1.129
R3279 VDD.n3703 VDD.n3702 0.858
R3280 VDD.n4300 VDD.n4299 0.849
R3281 VDD.n3698 VDD.n3697 0.849
R3282 VDD.n4297 VDD.n4296 0.849
R3283 VDD.n2683 VDD.n2682 0.77
R3284 VDD.n2948 VDD.n2947 0.77
R3285 VDD.n1724 VDD.n1723 0.77
R3286 VDD.n1269 VDD.n1268 0.77
R3287 VDD.n1849 VDD.n1848 0.77
R3288 VDD.n1861 VDD.n1860 0.77
R3289 VDD.n3302 VDD.n3301 0.77
R3290 VDD.n3309 VDD.n3308 0.77
R3291 VDD.n1474 VDD.n1473 0.77
R3292 VDD.n1484 VDD.n1483 0.77
R3293 VDD.n1623 VDD.n1622 0.77
R3294 VDD.n1616 VDD.n1615 0.77
R3295 VDD.n2123 VDD.n2122 0.77
R3296 VDD.n543 VDD.n542 0.77
R3297 VDD.n2004 VDD.n2003 0.646
R3298 VDD.n2032 VDD.n2031 0.646
R3299 VDD.n260 VDD.n257 0.646
R3300 VDD.n3547 VDD.n3546 0.646
R3301 VDD.n666 VDD.n663 0.646
R3302 VDD.n2269 VDD.n2268 0.646
R3303 VDD.n1087 VDD.n1084 0.646
R3304 VDD.n1373 VDD.n1372 0.646
R3305 VDD.n3285 VDD.n3284 0.646
R3306 VDD.n3204 VDD.n3203 0.646
R3307 VDD.n2983 VDD.n2980 0.646
R3308 VDD.n3100 VDD.n3099 0.646
R3309 VDD.n1992 VDD.n1991 0.471
R3310 VDD.n355 VDD.n352 0.471
R3311 VDD.n574 VDD.n573 0.471
R3312 VDD.n403 VDD.n402 0.471
R3313 VDD.n633 VDD.n632 0.471
R3314 VDD.n2044 VDD.n2043 0.471
R3315 VDD.n334 VDD.n331 0.471
R3316 VDD.n3535 VDD.n3534 0.471
R3317 VDD.n741 VDD.n738 0.471
R3318 VDD.n2281 VDD.n2280 0.471
R3319 VDD.n1589 VDD.n1588 0.471
R3320 VDD.n1165 VDD.n1162 0.471
R3321 VDD.n1532 VDD.n1531 0.471
R3322 VDD.n3338 VDD.n3337 0.471
R3323 VDD.n1385 VDD.n1384 0.471
R3324 VDD.n1810 VDD.n1809 0.471
R3325 VDD.n3273 VDD.n3272 0.471
R3326 VDD.n3058 VDD.n3055 0.471
R3327 VDD.n3397 VDD.n3396 0.471
R3328 VDD.n3112 VDD.n3111 0.471
R3329 VDD.n1166 VDD.n1129 0.47
R3330 VDD.n3059 VDD.n3022 0.449
R3331 VDD.n1903 VDD.n1901 0.428
R3332 VDD.n335 VDD.n286 0.428
R3333 VDD.n742 VDD.n693 0.428
R3334 VDD.n3087 VDD.n3085 0.428
R3335 VDD.n425 VDD.n420 0.428
R3336 VDD.n335 VDD.n279 0.416
R3337 VDD.n1903 VDD.n1899 0.416
R3338 VDD.n742 VDD.n686 0.416
R3339 VDD.n425 VDD.n423 0.416
R3340 VDD.n425 VDD.n424 0.416
R3341 VDD.n426 VDD.n425 0.416
R3342 VDD.n1166 VDD.n1121 0.416
R3343 VDD.n1166 VDD.n1118 0.416
R3344 VDD.n1832 VDD.n1831 0.416
R3345 VDD.n1831 VDD.n1829 0.416
R3346 VDD.n3059 VDD.n3015 0.416
R3347 VDD.n3059 VDD.n3012 0.416
R3348 VDD.n728 VDD.n725 0.376
R3349 VDD.n728 VDD.n727 0.376
R3350 VDD.n722 VDD.n719 0.376
R3351 VDD.n722 VDD.n721 0.376
R3352 VDD.n2306 VDD.n2301 0.376
R3353 VDD.n2314 VDD.n2309 0.376
R3354 VDD.n2069 VDD.n2064 0.376
R3355 VDD.n2077 VDD.n2072 0.376
R3356 VDD.n1969 VDD.n1964 0.376
R3357 VDD.n1961 VDD.n1956 0.376
R3358 VDD.n321 VDD.n318 0.376
R3359 VDD.n321 VDD.n320 0.376
R3360 VDD.n315 VDD.n312 0.376
R3361 VDD.n315 VDD.n314 0.376
R3362 VDD.n3512 VDD.n3507 0.376
R3363 VDD.n3504 VDD.n3499 0.376
R3364 VDD.n370 VDD.n367 0.376
R3365 VDD.n370 VDD.n369 0.376
R3366 VDD.n382 VDD.n379 0.376
R3367 VDD.n382 VDD.n381 0.376
R3368 VDD.n600 VDD.n595 0.376
R3369 VDD.n609 VDD.n603 0.376
R3370 VDD.n1152 VDD.n1149 0.376
R3371 VDD.n1152 VDD.n1151 0.376
R3372 VDD.n1146 VDD.n1143 0.376
R3373 VDD.n1146 VDD.n1145 0.376
R3374 VDD.n1566 VDD.n1561 0.376
R3375 VDD.n1558 VDD.n1552 0.376
R3376 VDD.n1787 VDD.n1782 0.376
R3377 VDD.n1779 VDD.n1774 0.376
R3378 VDD.n1410 VDD.n1405 0.376
R3379 VDD.n1418 VDD.n1413 0.376
R3380 VDD.n3137 VDD.n3132 0.376
R3381 VDD.n3145 VDD.n3140 0.376
R3382 VDD.n3250 VDD.n3245 0.376
R3383 VDD.n3242 VDD.n3237 0.376
R3384 VDD.n3045 VDD.n3042 0.376
R3385 VDD.n3045 VDD.n3044 0.376
R3386 VDD.n3039 VDD.n3036 0.376
R3387 VDD.n3039 VDD.n3038 0.376
R3388 VDD.n3364 VDD.n3359 0.376
R3389 VDD.n3373 VDD.n3367 0.376
R3390 VDD.n1903 VDD.n1902 0.327
R3391 VDD.n1831 VDD.n1830 0.327
R3392 VDD.n3087 VDD.n3086 0.327
R3393 VDD.n335 VDD.n298 0.312
R3394 VDD.n742 VDD.n705 0.312
R3395 VDD.n425 VDD.n415 0.312
R3396 VDD.n1980 VDD.n1979 0.288
R3397 VDD.n2056 VDD.n2055 0.288
R3398 VDD.n269 VDD.n266 0.288
R3399 VDD.n3523 VDD.n3522 0.288
R3400 VDD.n675 VDD.n672 0.288
R3401 VDD.n2293 VDD.n2292 0.288
R3402 VDD.n1096 VDD.n1093 0.288
R3403 VDD.n1397 VDD.n1396 0.288
R3404 VDD.n1798 VDD.n1797 0.288
R3405 VDD.n3261 VDD.n3260 0.288
R3406 VDD.n2992 VDD.n2989 0.288
R3407 VDD.n3124 VDD.n3123 0.288
R3408 VDD.n3558 VDD.n3557 0.219
R3409 VDD.n2256 VDD.n2255 0.219
R3410 VDD.n2376 VDD.n657 0.213
R3411 VDD.n2394 VDD.n654 0.213
R3412 VDD.n3585 VDD.n3584 0.213
R3413 VDD.n3457 VDD.n3456 0.213
R3414 VDD.n2225 VDD.n2224 0.213
R3415 VDD.n2358 VDD.n2357 0.213
R3416 VDD.n3296 VDD.n3295 0.208
R3417 VDD.n1629 VDD.n1628 0.208
R3418 VDD.n2120 VDD.n2119 0.208
R3419 VDD.n1732 VDD.n1729 0.208
R3420 VDD.n3187 VDD.n2660 0.208
R3421 VDD.n2819 VDD.n2818 0.189
R3422 VDD.n2793 VDD.n2792 0.189
R3423 VDD.n1245 VDD.n1244 0.189
R3424 VDD.n809 VDD.n808 0.189
R3425 VDD.n783 VDD.n782 0.189
R3426 VDD.n2552 VDD.n2551 0.189
R3427 VDD.n2525 VDD.n2524 0.189
R3428 VDD.n991 VDD.n990 0.189
R3429 VDD.n965 VDD.n964 0.189
R3430 VDD.n1038 VDD.n1037 0.189
R3431 VDD.n1051 VDD.n1050 0.189
R3432 VDD.n224 VDD.n223 0.189
R3433 VDD.n198 VDD.n197 0.189
R3434 VDD.n519 VDD.n518 0.189
R3435 VDD.n505 VDD.n504 0.189
R3436 VDD.n1231 VDD.n1230 0.189
R3437 VDD.n2924 VDD.n2923 0.189
R3438 VDD.n2910 VDD.n2909 0.189
R3439 VDD.n2459 VDD.n2458 0.188
R3440 VDD.n2446 VDD.n2445 0.188
R3441 VDD.n2611 VDD.n2610 0.188
R3442 VDD.n2598 VDD.n2597 0.188
R3443 VDD.n1328 VDD.n1327 0.188
R3444 VDD.n1342 VDD.n1341 0.188
R3445 VDD.n2162 VDD.n2161 0.188
R3446 VDD.n2149 VDD.n2148 0.188
R3447 VDD.n1686 VDD.n1685 0.188
R3448 VDD.n1700 VDD.n1699 0.188
R3449 VDD.n2722 VDD.n2721 0.188
R3450 VDD.n2709 VDD.n2708 0.188
R3451 VDD.n3757 VDD.n3756 0.188
R3452 VDD.n3799 VDD.n3798 0.188
R3453 VDD.n3910 VDD.n3909 0.188
R3454 VDD.n3858 VDD.n3857 0.188
R3455 VDD.n4021 VDD.n4020 0.188
R3456 VDD.n3969 VDD.n3968 0.188
R3457 VDD.n4132 VDD.n4131 0.188
R3458 VDD.n4080 VDD.n4079 0.188
R3459 VDD.n4243 VDD.n4242 0.188
R3460 VDD.n4191 VDD.n4190 0.188
R3461 VDD.n4359 VDD.n4358 0.188
R3462 VDD.n4401 VDD.n4400 0.188
R3463 VDD.n4519 VDD.n4518 0.188
R3464 VDD.n4467 VDD.n4466 0.188
R3465 VDD.n4637 VDD.n4636 0.188
R3466 VDD.n4585 VDD.n4584 0.188
R3467 VDD.n4690 VDD.n4689 0.188
R3468 VDD.n27 VDD.n26 0.188
R3469 VDD.n3315 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/GATE 0.181
R3470 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/GATE VDD.n1609 0.181
R3471 VDD.n549 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/GATE 0.181
R3472 VDD.n1275 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/GATE 0.181
R3473 VDD.n2954 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/GATE 0.181
R3474 VDD.n3071 VDD.n2842 0.18
R3475 VDD.n1858 VDD.n831 0.18
R3476 VDD.n3306 VDD.n2574 0.18
R3477 VDD.n3434 VDD.n2416 0.18
R3478 VDD.n1620 VDD.n1013 0.18
R3479 VDD.n1466 VDD.n1363 0.18
R3480 VDD.n250 VDD.n247 0.18
R3481 VDD.n2129 VDD.n2127 0.18
R3482 VDD.n547 VDD.n540 0.18
R3483 VDD.n1728 VDD.n1721 0.18
R3484 VDD.n1273 VDD.n1266 0.18
R3485 VDD.n2689 VDD.n2687 0.18
R3486 VDD.n2952 VDD.n2945 0.18
R3487 VDD.n2826 VDD.n2825 0.178
R3488 VDD.n2781 VDD.n2780 0.178
R3489 VDD.n816 VDD.n815 0.178
R3490 VDD.n771 VDD.n770 0.178
R3491 VDD.n2559 VDD.n2558 0.178
R3492 VDD.n2514 VDD.n2513 0.178
R3493 VDD.n2591 VDD.n2590 0.178
R3494 VDD.n2439 VDD.n2438 0.178
R3495 VDD.n998 VDD.n997 0.178
R3496 VDD.n953 VDD.n952 0.178
R3497 VDD.n1349 VDD.n1348 0.178
R3498 VDD.n231 VDD.n230 0.178
R3499 VDD.n186 VDD.n185 0.178
R3500 VDD.n2142 VDD.n2141 0.178
R3501 VDD.n1707 VDD.n1706 0.178
R3502 VDD.n2702 VDD.n2701 0.178
R3503 VDD.n2470 VDD.n2469 0.177
R3504 VDD.n2622 VDD.n2621 0.177
R3505 VDD.n1062 VDD.n1061 0.177
R3506 VDD.n1031 VDD.n1030 0.177
R3507 VDD.n1316 VDD.n1315 0.177
R3508 VDD.n2173 VDD.n2172 0.177
R3509 VDD.n493 VDD.n492 0.177
R3510 VDD.n526 VDD.n525 0.177
R3511 VDD.n1674 VDD.n1673 0.177
R3512 VDD.n1219 VDD.n1218 0.177
R3513 VDD.n1252 VDD.n1251 0.177
R3514 VDD.n2733 VDD.n2732 0.177
R3515 VDD.n2898 VDD.n2897 0.177
R3516 VDD.n2931 VDD.n2930 0.177
R3517 VDD.n3769 VDD.n3768 0.177
R3518 VDD.n3811 VDD.n3810 0.177
R3519 VDD.n3922 VDD.n3921 0.177
R3520 VDD.n3870 VDD.n3869 0.177
R3521 VDD.n4033 VDD.n4032 0.177
R3522 VDD.n3981 VDD.n3980 0.177
R3523 VDD.n4144 VDD.n4143 0.177
R3524 VDD.n4092 VDD.n4091 0.177
R3525 VDD.n4255 VDD.n4254 0.177
R3526 VDD.n4203 VDD.n4202 0.177
R3527 VDD.n4371 VDD.n4370 0.177
R3528 VDD.n4413 VDD.n4412 0.177
R3529 VDD.n4531 VDD.n4530 0.177
R3530 VDD.n4479 VDD.n4478 0.177
R3531 VDD.n4649 VDD.n4648 0.177
R3532 VDD.n4597 VDD.n4596 0.177
R3533 VDD.n4702 VDD.n4701 0.177
R3534 VDD.n39 VDD.n38 0.177
R3535 VDD.n2857 VDD.n2421 0.172
R3536 VDD.n3194 VDD.n3191 0.172
R3537 VDD.n1277 VDD.n1276 0.172
R3538 VDD.n1637 VDD.n1633 0.172
R3539 VDD.n2020 VDD.n2016 0.172
R3540 VDD.n2016 VDD.n2013 0.172
R3541 VDD.n551 VDD.n550 0.172
R3542 VDD.n552 VDD.n551 0.172
R3543 VDD.n3607 VDD.n3603 0.172
R3544 VDD.n3603 VDD.n3599 0.172
R3545 VDD.n3599 VDD.n3595 0.172
R3546 VDD.n3595 VDD.n3591 0.172
R3547 VDD.n2664 VDD.n256 0.172
R3548 VDD.n2668 VDD.n2664 0.172
R3549 VDD.n2672 VDD.n2668 0.172
R3550 VDD.n3557 VDD.n3556 0.172
R3551 VDD.n3556 VDD.n3555 0.172
R3552 VDD.n3555 VDD.n3554 0.172
R3553 VDD.n1508 VDD.n1503 0.172
R3554 VDD.n1503 VDD.n1500 0.172
R3555 VDD.n1500 VDD.n1497 0.172
R3556 VDD.n1497 VDD.n662 0.172
R3557 VDD.n2364 VDD.n2361 0.172
R3558 VDD.n2367 VDD.n2364 0.172
R3559 VDD.n2370 VDD.n2367 0.172
R3560 VDD.n2375 VDD.n2370 0.172
R3561 VDD.n2382 VDD.n2379 0.172
R3562 VDD.n2385 VDD.n2382 0.172
R3563 VDD.n2388 VDD.n2385 0.172
R3564 VDD.n2393 VDD.n2388 0.172
R3565 VDD.n2400 VDD.n2397 0.172
R3566 VDD.n2403 VDD.n2400 0.172
R3567 VDD.n2406 VDD.n2403 0.172
R3568 VDD.n2411 VDD.n2406 0.172
R3569 VDD.n3455 VDD.n3452 0.172
R3570 VDD.n3452 VDD.n3449 0.172
R3571 VDD.n3449 VDD.n3446 0.172
R3572 VDD.n2257 VDD.n2256 0.172
R3573 VDD.n2258 VDD.n2257 0.172
R3574 VDD.n2259 VDD.n2258 0.172
R3575 VDD.n1884 VDD.n1880 0.172
R3576 VDD.n1888 VDD.n1884 0.172
R3577 VDD.n1892 VDD.n1888 0.172
R3578 VDD.n1898 VDD.n1892 0.172
R3579 VDD.n2223 VDD.n2219 0.172
R3580 VDD.n2219 VDD.n2215 0.172
R3581 VDD.n2215 VDD.n2211 0.172
R3582 VDD.n2211 VDD.n2207 0.17
R3583 VDD.n2833 VDD.n2832 0.166
R3584 VDD.n2772 VDD.n2771 0.166
R3585 VDD.n1259 VDD.n1258 0.166
R3586 VDD.n823 VDD.n822 0.166
R3587 VDD.n762 VDD.n761 0.166
R3588 VDD.n2566 VDD.n2565 0.166
R3589 VDD.n2505 VDD.n2504 0.166
R3590 VDD.n1005 VDD.n1004 0.166
R3591 VDD.n944 VDD.n943 0.166
R3592 VDD.n1024 VDD.n1023 0.166
R3593 VDD.n238 VDD.n237 0.166
R3594 VDD.n177 VDD.n176 0.166
R3595 VDD.n533 VDD.n532 0.166
R3596 VDD.n2938 VDD.n2937 0.166
R3597 VDD.n2479 VDD.n2478 0.166
R3598 VDD.n2432 VDD.n2431 0.166
R3599 VDD.n2631 VDD.n2630 0.166
R3600 VDD.n2584 VDD.n2583 0.166
R3601 VDD.n1071 VDD.n1070 0.166
R3602 VDD.n1306 VDD.n1305 0.166
R3603 VDD.n1356 VDD.n1355 0.166
R3604 VDD.n2183 VDD.n2182 0.166
R3605 VDD.n2135 VDD.n2134 0.166
R3606 VDD.n483 VDD.n482 0.166
R3607 VDD.n1664 VDD.n1663 0.166
R3608 VDD.n1714 VDD.n1713 0.166
R3609 VDD.n1209 VDD.n1208 0.166
R3610 VDD.n2743 VDD.n2742 0.166
R3611 VDD.n2695 VDD.n2694 0.166
R3612 VDD.n2888 VDD.n2887 0.166
R3613 VDD.n3742 VDD.n3741 0.166
R3614 VDD.n3784 VDD.n3783 0.166
R3615 VDD.n3895 VDD.n3894 0.166
R3616 VDD.n3843 VDD.n3842 0.166
R3617 VDD.n4006 VDD.n4005 0.166
R3618 VDD.n3954 VDD.n3953 0.166
R3619 VDD.n4117 VDD.n4116 0.166
R3620 VDD.n4065 VDD.n4064 0.166
R3621 VDD.n4228 VDD.n4227 0.166
R3622 VDD.n4176 VDD.n4175 0.166
R3623 VDD.n4344 VDD.n4343 0.166
R3624 VDD.n4386 VDD.n4385 0.166
R3625 VDD.n4504 VDD.n4503 0.166
R3626 VDD.n4452 VDD.n4451 0.166
R3627 VDD.n4622 VDD.n4621 0.166
R3628 VDD.n4570 VDD.n4569 0.166
R3629 VDD.n4675 VDD.n4674 0.166
R3630 VDD.n12 VDD.n11 0.166
R3631 VDD.n2955 VDD.n2954 0.161
R3632 VDD.n549 VDD.n457 0.161
R3633 VDD.n2119 VDD.n2118 0.161
R3634 VDD.n1275 VDD.n1197 0.161
R3635 VDD.n1734 VDD.n1732 0.161
R3636 VDD.n3187 VDD.n3186 0.161
R3637 VDD.n2762 VDD.n2761 0.156
R3638 VDD.n752 VDD.n751 0.156
R3639 VDD.n3313 VDD.n2491 0.156
R3640 VDD.n3297 VDD.n2657 0.156
R3641 VDD.n1611 VDD.n1083 0.156
R3642 VDD.n1627 VDD.n930 0.156
R3643 VDD.n167 VDD.n166 0.156
R3644 VDD.n2196 VDD.n2195 0.156
R3645 VDD.n3619 VDD.n251 0.156
R3646 VDD.n1840 VDD.n925 0.156
R3647 VDD.n1869 VDD.n745 0.156
R3648 VDD.n3079 VDD.n2755 0.156
R3649 VDD.n2862 VDD.n2861 0.156
R3650 VDD.n2967 VDD.n2966 0.15
R3651 VDD.n3251 VDD.n3243 0.15
R3652 VDD.n3196 VDD.n2414 0.15
R3653 VDD.n3374 VDD.n3365 0.15
R3654 VDD.n3418 VDD.n3415 0.15
R3655 VDD.n1419 VDD.n1411 0.15
R3656 VDD.n1462 VDD.n1459 0.15
R3657 VDD.n1567 VDD.n1559 0.15
R3658 VDD.n1512 VDD.n1510 0.15
R3659 VDD.n446 VDD.n445 0.15
R3660 VDD.n1970 VDD.n1962 0.15
R3661 VDD.n1917 VDD.n657 0.15
R3662 VDD.n610 VDD.n601 0.15
R3663 VDD.n654 VDD.n651 0.15
R3664 VDD.n2078 VDD.n2070 0.15
R3665 VDD.n3570 VDD.n3569 0.15
R3666 VDD.n3513 VDD.n3505 0.15
R3667 VDD.n3459 VDD.n3457 0.15
R3668 VDD.n2244 VDD.n2243 0.15
R3669 VDD.n2315 VDD.n2307 0.15
R3670 VDD.n2357 VDD.n2354 0.15
R3671 VDD.n1186 VDD.n1185 0.15
R3672 VDD.n1788 VDD.n1780 0.15
R3673 VDD.n3146 VDD.n3138 0.15
R3674 VDD.n4298 VDD.n4297 0.149
R3675 VDD.n3446 VDD.n3443 0.146
R3676 VDD.n2678 VDD.n2672 0.146
R3677 VDD.n2815 VDD.n2813 0.144
R3678 VDD.n3062 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/BULK 0.144
R3679 VDD.n805 VDD.n803 0.144
R3680 VDD.n2548 VDD.n2546 0.144
R3681 VDD.n3294 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/BULK 0.144
R3682 VDD.n2454 VDD.n2451 0.144
R3683 VDD.n2606 VDD.n2603 0.144
R3684 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/BULK VDD.n3316 0.144
R3685 VDD.n987 VDD.n985 0.144
R3686 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/BULK VDD.n929 0.144
R3687 VDD.n1046 VDD.n1043 0.144
R3688 VDD.n1338 VDD.n1336 0.144
R3689 VDD.n1608 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/BULK 0.144
R3690 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/BULK VDD.n252 0.144
R3691 VDD.n2013 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/BULK 0.144
R3692 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/BULK VDD.n552 0.144
R3693 VDD.n220 VDD.n218 0.144
R3694 VDD.n2157 VDD.n2154 0.144
R3695 VDD.n515 VDD.n513 0.144
R3696 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/BULK VDD.n1906 0.144
R3697 VDD.n3584 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/BULK 0.144
R3698 VDD.n3554 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/BULK 0.144
R3699 VDD.n2225 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/BULK 0.144
R3700 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/BULK VDD.n2259 0.144
R3701 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/BULK VDD.n744 0.144
R3702 VDD.n1696 VDD.n1694 0.144
R3703 VDD.n1835 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/BULK 0.144
R3704 VDD.n1241 VDD.n1239 0.144
R3705 VDD.n2717 VDD.n2714 0.144
R3706 VDD.n2920 VDD.n2918 0.144
R3707 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/BULK VDD.n3090 0.144
R3708 VDD.n3585 VDD.n256 0.137
R3709 VDD.n3456 VDD.n3455 0.137
R3710 VDD.n3306 VDD.n3303 0.132
R3711 VDD.n3310 VDD.n3306 0.132
R3712 VDD.n1624 VDD.n1620 0.132
R3713 VDD.n1620 VDD.n1617 0.132
R3714 VDD.n2836 VDD.n2834 0.127
R3715 VDD.n2829 VDD.n2827 0.127
R3716 VDD.n2822 VDD.n2820 0.127
R3717 VDD.n826 VDD.n824 0.127
R3718 VDD.n819 VDD.n817 0.127
R3719 VDD.n812 VDD.n810 0.127
R3720 VDD.n2569 VDD.n2567 0.127
R3721 VDD.n2562 VDD.n2560 0.127
R3722 VDD.n2555 VDD.n2553 0.127
R3723 VDD.n2447 VDD.n2444 0.127
R3724 VDD.n2440 VDD.n2437 0.127
R3725 VDD.n2433 VDD.n2430 0.127
R3726 VDD.n2599 VDD.n2596 0.127
R3727 VDD.n2592 VDD.n2589 0.127
R3728 VDD.n2585 VDD.n2582 0.127
R3729 VDD.n1008 VDD.n1006 0.127
R3730 VDD.n1001 VDD.n999 0.127
R3731 VDD.n994 VDD.n992 0.127
R3732 VDD.n1039 VDD.n1036 0.127
R3733 VDD.n1032 VDD.n1029 0.127
R3734 VDD.n1025 VDD.n1022 0.127
R3735 VDD.n1345 VDD.n1343 0.127
R3736 VDD.n1352 VDD.n1350 0.127
R3737 VDD.n1359 VDD.n1357 0.127
R3738 VDD.n241 VDD.n239 0.127
R3739 VDD.n234 VDD.n232 0.127
R3740 VDD.n227 VDD.n225 0.127
R3741 VDD.n2150 VDD.n2147 0.127
R3742 VDD.n2143 VDD.n2140 0.127
R3743 VDD.n2136 VDD.n2133 0.127
R3744 VDD.n522 VDD.n520 0.127
R3745 VDD.n529 VDD.n527 0.127
R3746 VDD.n536 VDD.n534 0.127
R3747 VDD.n1703 VDD.n1701 0.127
R3748 VDD.n1710 VDD.n1708 0.127
R3749 VDD.n1717 VDD.n1715 0.127
R3750 VDD.n1248 VDD.n1246 0.127
R3751 VDD.n1255 VDD.n1253 0.127
R3752 VDD.n1262 VDD.n1260 0.127
R3753 VDD.n2710 VDD.n2707 0.127
R3754 VDD.n2703 VDD.n2700 0.127
R3755 VDD.n2696 VDD.n2693 0.127
R3756 VDD.n2927 VDD.n2925 0.127
R3757 VDD.n2934 VDD.n2932 0.127
R3758 VDD.n2941 VDD.n2939 0.127
R3759 VDD.n2397 VDD.n2394 0.125
R3760 VDD.n3754 VDD.n3753 0.121
R3761 VDD.n3796 VDD.n3795 0.121
R3762 VDD.n3907 VDD.n3906 0.121
R3763 VDD.n3855 VDD.n3854 0.121
R3764 VDD.n4018 VDD.n4017 0.121
R3765 VDD.n3966 VDD.n3965 0.121
R3766 VDD.n4129 VDD.n4128 0.121
R3767 VDD.n4077 VDD.n4076 0.121
R3768 VDD.n4240 VDD.n4239 0.121
R3769 VDD.n4188 VDD.n4187 0.121
R3770 VDD.n4356 VDD.n4355 0.121
R3771 VDD.n4398 VDD.n4397 0.121
R3772 VDD.n4516 VDD.n4515 0.121
R3773 VDD.n4464 VDD.n4463 0.121
R3774 VDD.n4634 VDD.n4633 0.121
R3775 VDD.n4582 VDD.n4581 0.121
R3776 VDD.n4687 VDD.n4686 0.121
R3777 VDD.n24 VDD.n23 0.121
R3778 VDD.n4537 VDD.n4536 0.119
R3779 VDD.n2976 VDD.n2975 0.114
R3780 VDD.n2973 VDD.n2972 0.114
R3781 VDD.n2970 VDD.n2969 0.114
R3782 VDD.n2964 VDD.n2963 0.114
R3783 VDD.n2961 VDD.n2960 0.114
R3784 VDD.n2958 VDD.n2957 0.114
R3785 VDD.n3287 VDD.n3279 0.114
R3786 VDD.n3275 VDD.n3267 0.114
R3787 VDD.n3263 VDD.n3255 0.114
R3788 VDD.n3233 VDD.n3231 0.114
R3789 VDD.n3221 VDD.n3219 0.114
R3790 VDD.n3208 VDD.n3206 0.114
R3791 VDD.n3330 VDD.n3328 0.114
R3792 VDD.n3342 VDD.n3340 0.114
R3793 VDD.n3355 VDD.n3353 0.114
R3794 VDD.n3387 VDD.n3378 0.114
R3795 VDD.n3399 VDD.n3391 0.114
R3796 VDD.n3411 VDD.n3403 0.114
R3797 VDD.n1377 VDD.n1375 0.114
R3798 VDD.n1389 VDD.n1387 0.114
R3799 VDD.n1401 VDD.n1399 0.114
R3800 VDD.n1431 VDD.n1423 0.114
R3801 VDD.n1443 VDD.n1435 0.114
R3802 VDD.n1455 VDD.n1447 0.114
R3803 VDD.n1603 VDD.n1595 0.114
R3804 VDD.n1591 VDD.n1583 0.114
R3805 VDD.n1579 VDD.n1571 0.114
R3806 VDD.n1548 VDD.n1546 0.114
R3807 VDD.n1536 VDD.n1534 0.114
R3808 VDD.n1524 VDD.n1522 0.114
R3809 VDD.n437 VDD.n436 0.114
R3810 VDD.n440 VDD.n439 0.114
R3811 VDD.n443 VDD.n442 0.114
R3812 VDD.n449 VDD.n448 0.114
R3813 VDD.n452 VDD.n451 0.114
R3814 VDD.n455 VDD.n454 0.114
R3815 VDD.n2006 VDD.n1998 0.114
R3816 VDD.n1994 VDD.n1986 0.114
R3817 VDD.n1982 VDD.n1974 0.114
R3818 VDD.n1952 VDD.n1950 0.114
R3819 VDD.n1940 VDD.n1938 0.114
R3820 VDD.n1928 VDD.n1926 0.114
R3821 VDD.n566 VDD.n564 0.114
R3822 VDD.n578 VDD.n576 0.114
R3823 VDD.n591 VDD.n589 0.114
R3824 VDD.n623 VDD.n614 0.114
R3825 VDD.n635 VDD.n627 0.114
R3826 VDD.n647 VDD.n639 0.114
R3827 VDD.n2036 VDD.n2034 0.114
R3828 VDD.n2048 VDD.n2046 0.114
R3829 VDD.n2060 VDD.n2058 0.114
R3830 VDD.n2090 VDD.n2082 0.114
R3831 VDD.n2102 VDD.n2094 0.114
R3832 VDD.n2114 VDD.n2106 0.114
R3833 VDD.n3579 VDD.n3578 0.114
R3834 VDD.n3576 VDD.n3575 0.114
R3835 VDD.n3573 VDD.n3572 0.114
R3836 VDD.n3567 VDD.n3566 0.114
R3837 VDD.n3564 VDD.n3563 0.114
R3838 VDD.n3561 VDD.n3560 0.114
R3839 VDD.n3549 VDD.n3541 0.114
R3840 VDD.n3537 VDD.n3529 0.114
R3841 VDD.n3525 VDD.n3517 0.114
R3842 VDD.n3495 VDD.n3493 0.114
R3843 VDD.n3483 VDD.n3481 0.114
R3844 VDD.n3470 VDD.n3468 0.114
R3845 VDD.n2235 VDD.n2234 0.114
R3846 VDD.n2238 VDD.n2237 0.114
R3847 VDD.n2241 VDD.n2240 0.114
R3848 VDD.n2247 VDD.n2246 0.114
R3849 VDD.n2250 VDD.n2249 0.114
R3850 VDD.n2253 VDD.n2252 0.114
R3851 VDD.n2273 VDD.n2271 0.114
R3852 VDD.n2285 VDD.n2283 0.114
R3853 VDD.n2297 VDD.n2295 0.114
R3854 VDD.n2327 VDD.n2319 0.114
R3855 VDD.n2339 VDD.n2331 0.114
R3856 VDD.n2350 VDD.n2343 0.114
R3857 VDD.n1177 VDD.n1176 0.114
R3858 VDD.n1180 VDD.n1179 0.114
R3859 VDD.n1183 VDD.n1182 0.114
R3860 VDD.n1189 VDD.n1188 0.114
R3861 VDD.n1192 VDD.n1191 0.114
R3862 VDD.n1195 VDD.n1194 0.114
R3863 VDD.n1824 VDD.n1816 0.114
R3864 VDD.n1812 VDD.n1804 0.114
R3865 VDD.n1800 VDD.n1792 0.114
R3866 VDD.n1770 VDD.n1768 0.114
R3867 VDD.n1758 VDD.n1756 0.114
R3868 VDD.n1746 VDD.n1744 0.114
R3869 VDD.n3104 VDD.n3102 0.114
R3870 VDD.n3116 VDD.n3114 0.114
R3871 VDD.n3128 VDD.n3126 0.114
R3872 VDD.n3158 VDD.n3150 0.114
R3873 VDD.n3170 VDD.n3162 0.114
R3874 VDD.n3182 VDD.n3174 0.114
R3875 VDD.n2379 VDD.n2376 0.112
R3876 VDD.n2361 VDD.n2358 0.099
R3877 VDD.n2224 VDD.n2223 0.099
R3878 VDD.n1968 VDD.n1967 0.098
R3879 VDD.n374 VDD.n371 0.098
R3880 VDD.n599 VDD.n598 0.098
R3881 VDD.n384 VDD.n383 0.098
R3882 VDD.n608 VDD.n607 0.098
R3883 VDD.n2068 VDD.n2067 0.098
R3884 VDD.n325 VDD.n322 0.098
R3885 VDD.n3511 VDD.n3510 0.098
R3886 VDD.n732 VDD.n729 0.098
R3887 VDD.n2305 VDD.n2304 0.098
R3888 VDD.n1565 VDD.n1564 0.098
R3889 VDD.n1156 VDD.n1153 0.098
R3890 VDD.n1557 VDD.n1556 0.098
R3891 VDD.n3363 VDD.n3362 0.098
R3892 VDD.n1409 VDD.n1408 0.098
R3893 VDD.n1786 VDD.n1785 0.098
R3894 VDD.n3249 VDD.n3248 0.098
R3895 VDD.n3049 VDD.n3046 0.098
R3896 VDD.n3372 VDD.n3371 0.098
R3897 VDD.n3136 VDD.n3135 0.098
R3898 VDD.n3628 VDD.n3627 0.092
R3899 VDD.n1851 VDD.n924 0.092
R3900 VDD.n2850 VDD.n2849 0.092
R3901 VDD.n2954 VDD.n2857 0.088
R3902 VDD.n3191 VDD.n3187 0.088
R3903 VDD.n1276 VDD.n1275 0.088
R3904 VDD.n1732 VDD.n1637 0.088
R3905 VDD.n2119 VDD.n2020 0.088
R3906 VDD.n550 VDD.n549 0.088
R3907 VDD.n3608 VDD.n3607 0.085
R3908 VDD.n3063 VDD.n3062 0.079
R3909 VDD.n3419 VDD.n3418 0.079
R3910 VDD.n2358 VDD.n662 0.073
R3911 VDD.n2224 VDD.n1898 0.073
R3912 VDD.n1466 VDD.n1465 0.062
R3913 VDD.n1840 VDD.n1839 0.062
R3914 VDD.n2790 VDD.n2789 0.06
R3915 VDD.n2779 VDD.n2778 0.06
R3916 VDD.n2770 VDD.n2769 0.06
R3917 VDD.n780 VDD.n779 0.06
R3918 VDD.n769 VDD.n768 0.06
R3919 VDD.n760 VDD.n759 0.06
R3920 VDD.n2522 VDD.n2521 0.06
R3921 VDD.n2512 VDD.n2511 0.06
R3922 VDD.n2503 VDD.n2502 0.06
R3923 VDD.n2482 VDD.n2481 0.06
R3924 VDD.n2473 VDD.n2472 0.06
R3925 VDD.n2464 VDD.n2462 0.06
R3926 VDD.n2634 VDD.n2633 0.06
R3927 VDD.n2625 VDD.n2624 0.06
R3928 VDD.n2616 VDD.n2614 0.06
R3929 VDD.n962 VDD.n961 0.06
R3930 VDD.n951 VDD.n950 0.06
R3931 VDD.n942 VDD.n941 0.06
R3932 VDD.n1074 VDD.n1073 0.06
R3933 VDD.n1065 VDD.n1064 0.06
R3934 VDD.n1056 VDD.n1054 0.06
R3935 VDD.n1304 VDD.n1303 0.06
R3936 VDD.n1314 VDD.n1313 0.06
R3937 VDD.n1325 VDD.n1324 0.06
R3938 VDD.n195 VDD.n194 0.06
R3939 VDD.n184 VDD.n183 0.06
R3940 VDD.n175 VDD.n174 0.06
R3941 VDD.n2186 VDD.n2185 0.06
R3942 VDD.n2176 VDD.n2175 0.06
R3943 VDD.n2167 VDD.n2165 0.06
R3944 VDD.n481 VDD.n480 0.06
R3945 VDD.n491 VDD.n490 0.06
R3946 VDD.n502 VDD.n501 0.06
R3947 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/GATE VDD.n3614 0.06
R3948 VDD.n2376 VDD.n2375 0.06
R3949 VDD.n1662 VDD.n1661 0.06
R3950 VDD.n1672 VDD.n1671 0.06
R3951 VDD.n1683 VDD.n1682 0.06
R3952 VDD.n1207 VDD.n1206 0.06
R3953 VDD.n1217 VDD.n1216 0.06
R3954 VDD.n1228 VDD.n1227 0.06
R3955 VDD.n2746 VDD.n2745 0.06
R3956 VDD.n2736 VDD.n2735 0.06
R3957 VDD.n2727 VDD.n2725 0.06
R3958 VDD.n2886 VDD.n2885 0.06
R3959 VDD.n2896 VDD.n2895 0.06
R3960 VDD.n2907 VDD.n2906 0.06
R3961 VDD.n3771 VDD.n3749 0.06
R3962 VDD.n3762 VDD.n3760 0.06
R3963 VDD.n3813 VDD.n3791 0.06
R3964 VDD.n3804 VDD.n3802 0.06
R3965 VDD.n3924 VDD.n3902 0.06
R3966 VDD.n3915 VDD.n3913 0.06
R3967 VDD.n3872 VDD.n3850 0.06
R3968 VDD.n3863 VDD.n3861 0.06
R3969 VDD.n4035 VDD.n4013 0.06
R3970 VDD.n4026 VDD.n4024 0.06
R3971 VDD.n3983 VDD.n3961 0.06
R3972 VDD.n3974 VDD.n3972 0.06
R3973 VDD.n4146 VDD.n4124 0.06
R3974 VDD.n4137 VDD.n4135 0.06
R3975 VDD.n4094 VDD.n4072 0.06
R3976 VDD.n4085 VDD.n4083 0.06
R3977 VDD.n4257 VDD.n4235 0.06
R3978 VDD.n4248 VDD.n4246 0.06
R3979 VDD.n4205 VDD.n4183 0.06
R3980 VDD.n4196 VDD.n4194 0.06
R3981 VDD.n4373 VDD.n4351 0.06
R3982 VDD.n4364 VDD.n4362 0.06
R3983 VDD.n4415 VDD.n4393 0.06
R3984 VDD.n4406 VDD.n4404 0.06
R3985 VDD.n4533 VDD.n4511 0.06
R3986 VDD.n4524 VDD.n4522 0.06
R3987 VDD.n4481 VDD.n4459 0.06
R3988 VDD.n4472 VDD.n4470 0.06
R3989 VDD.n4651 VDD.n4629 0.06
R3990 VDD.n4642 VDD.n4640 0.06
R3991 VDD.n4599 VDD.n4577 0.06
R3992 VDD.n4590 VDD.n4588 0.06
R3993 VDD.n4704 VDD.n4682 0.06
R3994 VDD.n4695 VDD.n4693 0.06
R3995 VDD.n41 VDD.n19 0.06
R3996 VDD.n32 VDD.n30 0.06
R3997 VDD.n3438 VDD.n3437 0.057
R3998 VDD.n1485 VDD.n1481 0.057
R3999 VDD.n1862 VDD.n1858 0.057
R4000 VDD.n3084 VDD.n3083 0.057
R4001 VDD.n1478 VDD.n1475 0.055
R4002 VDD.n1912 VDD.n250 0.053
R4003 VDD.n894 VDD.n893 0.052
R4004 VDD.n3666 VDD.n3665 0.052
R4005 VDD.n3697 VDD.n3695 0.051
R4006 VDD.n120 VDD.n119 0.05
R4007 VDD.n3659 VDD.n3657 0.05
R4008 VDD.n3641 VDD.n3640 0.05
R4009 VDD.n133 VDD.n132 0.05
R4010 VDD.n135 VDD.n134 0.05
R4011 VDD.n3629 VDD.n3628 0.05
R4012 VDD.n912 VDD.n911 0.05
R4013 VDD.n879 VDD.n878 0.05
R4014 VDD.n881 VDD.n880 0.05
R4015 VDD.n865 VDD.n864 0.05
R4016 VDD.n924 VDD.n923 0.05
R4017 VDD.n848 VDD.n847 0.05
R4018 VDD.n2849 VDD.n2848 0.05
R4019 VDD.n109 VDD.n108 0.05
R4020 VDD.n3684 VDD.n3683 0.05
R4021 VDD.n61 VDD.n60 0.05
R4022 VDD.n71 VDD.n70 0.05
R4023 VDD.n89 VDD.n88 0.05
R4024 VDD.n3738 VDD.n3737 0.05
R4025 VDD.n3780 VDD.n3779 0.05
R4026 VDD.n3891 VDD.n3890 0.05
R4027 VDD.n3839 VDD.n3838 0.05
R4028 VDD.n4002 VDD.n4001 0.05
R4029 VDD.n3950 VDD.n3949 0.05
R4030 VDD.n4113 VDD.n4112 0.05
R4031 VDD.n4061 VDD.n4060 0.05
R4032 VDD.n4224 VDD.n4223 0.05
R4033 VDD.n4172 VDD.n4171 0.05
R4034 VDD.n4340 VDD.n4339 0.05
R4035 VDD.n4382 VDD.n4381 0.05
R4036 VDD.n4500 VDD.n4499 0.05
R4037 VDD.n4448 VDD.n4447 0.05
R4038 VDD.n4618 VDD.n4617 0.05
R4039 VDD.n4566 VDD.n4565 0.05
R4040 VDD.n4671 VDD.n4670 0.05
R4041 VDD.n8 VDD.n7 0.05
R4042 VDD.n3626 VDD.n3622 0.049
R4043 VDD.n2200 VDD.n2196 0.047
R4044 VDD.n2394 VDD.n2393 0.047
R4045 VDD.n1494 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/GATE 0.046
R4046 VDD.n1509 VDD.n1508 0.046
R4047 VDD.n1880 VDD.n1874 0.046
R4048 VDD.n1873 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/GATE 0.046
R4049 VDD.n152 VDD.n151 0.043
R4050 VDD.n120 VDD.n117 0.043
R4051 VDD.n120 VDD.n118 0.043
R4052 VDD.n133 VDD.n129 0.043
R4053 VDD.n133 VDD.n131 0.043
R4054 VDD.n3659 VDD.n3656 0.043
R4055 VDD.n3659 VDD.n3658 0.043
R4056 VDD.n3641 VDD.n3638 0.043
R4057 VDD.n3641 VDD.n3639 0.043
R4058 VDD.n3629 VDD.n160 0.043
R4059 VDD.n898 VDD.n897 0.043
R4060 VDD.n912 VDD.n909 0.043
R4061 VDD.n912 VDD.n910 0.043
R4062 VDD.n879 VDD.n875 0.043
R4063 VDD.n879 VDD.n877 0.043
R4064 VDD.n865 VDD.n862 0.043
R4065 VDD.n865 VDD.n863 0.043
R4066 VDD.n848 VDD.n845 0.043
R4067 VDD.n848 VDD.n846 0.043
R4068 VDD.n923 VDD.n832 0.043
R4069 VDD.n3670 VDD.n3669 0.043
R4070 VDD.n109 VDD.n106 0.043
R4071 VDD.n109 VDD.n107 0.043
R4072 VDD.n3684 VDD.n3681 0.043
R4073 VDD.n3684 VDD.n3682 0.043
R4074 VDD.n61 VDD.n59 0.043
R4075 VDD.n71 VDD.n68 0.043
R4076 VDD.n71 VDD.n69 0.043
R4077 VDD.n89 VDD.n86 0.043
R4078 VDD.n89 VDD.n87 0.043
R4079 VDD.n2848 VDD.n2843 0.043
R4080 VDD.n4267 VDD.n4266 0.043
R4081 VDD.n4274 VDD.n4273 0.043
R4082 VDD.n4281 VDD.n4280 0.043
R4083 VDD.n4288 VDD.n4287 0.043
R4084 VDD.n4655 VDD.n4654 0.043
R4085 VDD.n4419 VDD.n4418 0.043
R4086 VDD.n2201 VDD.n2200 0.042
R4087 VDD.n4295 VDD.n4294 0.042
R4088 VDD.n4301 VDD.n4300 0.042
R4089 VDD.n131 VDD.n130 0.041
R4090 VDD.n3656 VDD.n3655 0.041
R4091 VDD.n877 VDD.n876 0.041
R4092 VDD.n862 VDD.n861 0.041
R4093 VDD.n68 VDD.n67 0.041
R4094 VDD.n3630 VDD.n3629 0.041
R4095 VDD.n2848 VDD.n2847 0.041
R4096 VDD.n121 VDD.n120 0.041
R4097 VDD.n3644 VDD.n3641 0.041
R4098 VDD.n3662 VDD.n3659 0.041
R4099 VDD.n141 VDD.n133 0.041
R4100 VDD.n136 VDD.n135 0.041
R4101 VDD.n915 VDD.n912 0.041
R4102 VDD.n887 VDD.n879 0.041
R4103 VDD.n882 VDD.n881 0.041
R4104 VDD.n868 VDD.n865 0.041
R4105 VDD.n851 VDD.n848 0.041
R4106 VDD.n110 VDD.n109 0.041
R4107 VDD.n3689 VDD.n3684 0.041
R4108 VDD.n62 VDD.n61 0.041
R4109 VDD.n74 VDD.n71 0.041
R4110 VDD.n92 VDD.n89 0.041
R4111 VDD.n153 VDD.n152 0.041
R4112 VDD.n923 VDD.n922 0.041
R4113 VDD.n899 VDD.n898 0.041
R4114 VDD.n3671 VDD.n3670 0.041
R4115 VDD.n2820 VDD.n2817 0.038
R4116 VDD.n2769 VDD.n2768 0.038
R4117 VDD.n810 VDD.n807 0.038
R4118 VDD.n759 VDD.n758 0.038
R4119 VDD.n2553 VDD.n2550 0.038
R4120 VDD.n2502 VDD.n2501 0.038
R4121 VDD.n2484 VDD.n2482 0.038
R4122 VDD.n2449 VDD.n2447 0.038
R4123 VDD.n2636 VDD.n2634 0.038
R4124 VDD.n2601 VDD.n2599 0.038
R4125 VDD.n3430 VDD.n3427 0.038
R4126 VDD.n992 VDD.n989 0.038
R4127 VDD.n941 VDD.n940 0.038
R4128 VDD.n1076 VDD.n1074 0.038
R4129 VDD.n1041 VDD.n1039 0.038
R4130 VDD.n1303 VDD.n1302 0.038
R4131 VDD.n1343 VDD.n1340 0.038
R4132 VDD.n225 VDD.n222 0.038
R4133 VDD.n174 VDD.n173 0.038
R4134 VDD.n2188 VDD.n2186 0.038
R4135 VDD.n2152 VDD.n2150 0.038
R4136 VDD.n480 VDD.n479 0.038
R4137 VDD.n520 VDD.n517 0.038
R4138 VDD.n1661 VDD.n1660 0.038
R4139 VDD.n1701 VDD.n1698 0.038
R4140 VDD.n1206 VDD.n1205 0.038
R4141 VDD.n1246 VDD.n1243 0.038
R4142 VDD.n2748 VDD.n2746 0.038
R4143 VDD.n2712 VDD.n2710 0.038
R4144 VDD.n2885 VDD.n2884 0.038
R4145 VDD.n2925 VDD.n2922 0.038
R4146 VDD.n3075 VDD.n3071 0.038
R4147 VDD.n1465 VDD.n1462 0.037
R4148 VDD.n1839 VDD.n1835 0.037
R4149 VDD.n2969 VDD.n2968 0.034
R4150 VDD.n2965 VDD.n2964 0.034
R4151 VDD.n3255 VDD.n3253 0.034
R4152 VDD.n3235 VDD.n3233 0.034
R4153 VDD.n3357 VDD.n3355 0.034
R4154 VDD.n3378 VDD.n3376 0.034
R4155 VDD.n1403 VDD.n1401 0.034
R4156 VDD.n1423 VDD.n1421 0.034
R4157 VDD.n1571 VDD.n1569 0.034
R4158 VDD.n1550 VDD.n1548 0.034
R4159 VDD.n444 VDD.n443 0.034
R4160 VDD.n448 VDD.n447 0.034
R4161 VDD.n1974 VDD.n1972 0.034
R4162 VDD.n1954 VDD.n1952 0.034
R4163 VDD.n593 VDD.n591 0.034
R4164 VDD.n614 VDD.n612 0.034
R4165 VDD.n2062 VDD.n2060 0.034
R4166 VDD.n2082 VDD.n2080 0.034
R4167 VDD.n3591 VDD.n3585 0.034
R4168 VDD.n3572 VDD.n3571 0.034
R4169 VDD.n3568 VDD.n3567 0.034
R4170 VDD.n3517 VDD.n3515 0.034
R4171 VDD.n3497 VDD.n3495 0.034
R4172 VDD.n3456 VDD.n2411 0.034
R4173 VDD.n2242 VDD.n2241 0.034
R4174 VDD.n2246 VDD.n2245 0.034
R4175 VDD.n2299 VDD.n2297 0.034
R4176 VDD.n2319 VDD.n2317 0.034
R4177 VDD.n1184 VDD.n1183 0.034
R4178 VDD.n1188 VDD.n1187 0.034
R4179 VDD.n1792 VDD.n1790 0.034
R4180 VDD.n1772 VDD.n1770 0.034
R4181 VDD.n1855 VDD.n1851 0.034
R4182 VDD.n3130 VDD.n3128 0.034
R4183 VDD.n3150 VDD.n3148 0.034
R4184 VDD.n3424 VDD.n2419 0.034
R4185 VDD.n2827 VDD.n2824 0.033
R4186 VDD.n2782 VDD.n2779 0.033
R4187 VDD.n2778 VDD.n2777 0.033
R4188 VDD.n817 VDD.n814 0.033
R4189 VDD.n772 VDD.n769 0.033
R4190 VDD.n768 VDD.n767 0.033
R4191 VDD.n2560 VDD.n2557 0.033
R4192 VDD.n2515 VDD.n2512 0.033
R4193 VDD.n2511 VDD.n2510 0.033
R4194 VDD.n2475 VDD.n2473 0.033
R4195 VDD.n2472 VDD.n2471 0.033
R4196 VDD.n2442 VDD.n2440 0.033
R4197 VDD.n2627 VDD.n2625 0.033
R4198 VDD.n2624 VDD.n2623 0.033
R4199 VDD.n2594 VDD.n2592 0.033
R4200 VDD.n999 VDD.n996 0.033
R4201 VDD.n954 VDD.n951 0.033
R4202 VDD.n950 VDD.n949 0.033
R4203 VDD.n1067 VDD.n1065 0.033
R4204 VDD.n1064 VDD.n1063 0.033
R4205 VDD.n1034 VDD.n1032 0.033
R4206 VDD.n1313 VDD.n1312 0.033
R4207 VDD.n1317 VDD.n1314 0.033
R4208 VDD.n1350 VDD.n1347 0.033
R4209 VDD.n232 VDD.n229 0.033
R4210 VDD.n187 VDD.n184 0.033
R4211 VDD.n183 VDD.n182 0.033
R4212 VDD.n2178 VDD.n2176 0.033
R4213 VDD.n2175 VDD.n2174 0.033
R4214 VDD.n2145 VDD.n2143 0.033
R4215 VDD.n490 VDD.n489 0.033
R4216 VDD.n494 VDD.n491 0.033
R4217 VDD.n527 VDD.n524 0.033
R4218 VDD.n1671 VDD.n1670 0.033
R4219 VDD.n1675 VDD.n1672 0.033
R4220 VDD.n1708 VDD.n1705 0.033
R4221 VDD.n1216 VDD.n1215 0.033
R4222 VDD.n1220 VDD.n1217 0.033
R4223 VDD.n1253 VDD.n1250 0.033
R4224 VDD.n2738 VDD.n2736 0.033
R4225 VDD.n2735 VDD.n2734 0.033
R4226 VDD.n2705 VDD.n2703 0.033
R4227 VDD.n2895 VDD.n2894 0.033
R4228 VDD.n2899 VDD.n2896 0.033
R4229 VDD.n2932 VDD.n2929 0.033
R4230 VDD.n3771 VDD.n3770 0.033
R4231 VDD.n3813 VDD.n3812 0.033
R4232 VDD.n3924 VDD.n3923 0.033
R4233 VDD.n3872 VDD.n3871 0.033
R4234 VDD.n4035 VDD.n4034 0.033
R4235 VDD.n3983 VDD.n3982 0.033
R4236 VDD.n4146 VDD.n4145 0.033
R4237 VDD.n4094 VDD.n4093 0.033
R4238 VDD.n4257 VDD.n4256 0.033
R4239 VDD.n4205 VDD.n4204 0.033
R4240 VDD.n4373 VDD.n4372 0.033
R4241 VDD.n4415 VDD.n4414 0.033
R4242 VDD.n4533 VDD.n4532 0.033
R4243 VDD.n4481 VDD.n4480 0.033
R4244 VDD.n4651 VDD.n4650 0.033
R4245 VDD.n4599 VDD.n4598 0.033
R4246 VDD.n4704 VDD.n4703 0.033
R4247 VDD.n41 VDD.n40 0.033
R4248 VDD.n3437 VDD.n3434 0.032
R4249 VDD.n1509 VDD.n1494 0.032
R4250 VDD.n1874 VDD.n1873 0.032
R4251 VDD.n3083 VDD.n3079 0.032
R4252 VDD.n3737 VDD.n3736 0.031
R4253 VDD.n3779 VDD.n3778 0.031
R4254 VDD.n3890 VDD.n3889 0.031
R4255 VDD.n3838 VDD.n3837 0.031
R4256 VDD.n4001 VDD.n4000 0.031
R4257 VDD.n3949 VDD.n3948 0.031
R4258 VDD.n4112 VDD.n4111 0.031
R4259 VDD.n4060 VDD.n4059 0.031
R4260 VDD.n4223 VDD.n4222 0.031
R4261 VDD.n4171 VDD.n4170 0.031
R4262 VDD.n4339 VDD.n4338 0.031
R4263 VDD.n4381 VDD.n4380 0.031
R4264 VDD.n4499 VDD.n4498 0.031
R4265 VDD.n4447 VDD.n4446 0.031
R4266 VDD.n4617 VDD.n4616 0.031
R4267 VDD.n4565 VDD.n4564 0.031
R4268 VDD.n4670 VDD.n4669 0.031
R4269 VDD.n7 VDD.n6 0.031
R4270 VDD.n2972 VDD.n2971 0.03
R4271 VDD.n2962 VDD.n2961 0.03
R4272 VDD.n3267 VDD.n3265 0.03
R4273 VDD.n3223 VDD.n3221 0.03
R4274 VDD.n3344 VDD.n3342 0.03
R4275 VDD.n3391 VDD.n3389 0.03
R4276 VDD.n1391 VDD.n1389 0.03
R4277 VDD.n1435 VDD.n1433 0.03
R4278 VDD.n1583 VDD.n1581 0.03
R4279 VDD.n1538 VDD.n1536 0.03
R4280 VDD.n441 VDD.n440 0.03
R4281 VDD.n451 VDD.n450 0.03
R4282 VDD.n1986 VDD.n1984 0.03
R4283 VDD.n1942 VDD.n1940 0.03
R4284 VDD.n580 VDD.n578 0.03
R4285 VDD.n627 VDD.n625 0.03
R4286 VDD.n2050 VDD.n2048 0.03
R4287 VDD.n2094 VDD.n2092 0.03
R4288 VDD.n3575 VDD.n3574 0.03
R4289 VDD.n3565 VDD.n3564 0.03
R4290 VDD.n3529 VDD.n3527 0.03
R4291 VDD.n3485 VDD.n3483 0.03
R4292 VDD.n2239 VDD.n2238 0.03
R4293 VDD.n2249 VDD.n2248 0.03
R4294 VDD.n2287 VDD.n2285 0.03
R4295 VDD.n2331 VDD.n2329 0.03
R4296 VDD.n1181 VDD.n1180 0.03
R4297 VDD.n1191 VDD.n1190 0.03
R4298 VDD.n1804 VDD.n1802 0.03
R4299 VDD.n1760 VDD.n1758 0.03
R4300 VDD.n3118 VDD.n3116 0.03
R4301 VDD.n3162 VDD.n3160 0.03
R4302 VDD.n2834 VDD.n2831 0.028
R4303 VDD.n2789 VDD.n2787 0.028
R4304 VDD.n2773 VDD.n2770 0.028
R4305 VDD.n824 VDD.n821 0.028
R4306 VDD.n779 VDD.n777 0.028
R4307 VDD.n763 VDD.n760 0.028
R4308 VDD.n2567 VDD.n2564 0.028
R4309 VDD.n2521 VDD.n2519 0.028
R4310 VDD.n2506 VDD.n2503 0.028
R4311 VDD.n2481 VDD.n2480 0.028
R4312 VDD.n2466 VDD.n2464 0.028
R4313 VDD.n2435 VDD.n2433 0.028
R4314 VDD.n2633 VDD.n2632 0.028
R4315 VDD.n2618 VDD.n2616 0.028
R4316 VDD.n2587 VDD.n2585 0.028
R4317 VDD.n1006 VDD.n1003 0.028
R4318 VDD.n961 VDD.n959 0.028
R4319 VDD.n945 VDD.n942 0.028
R4320 VDD.n1073 VDD.n1072 0.028
R4321 VDD.n1058 VDD.n1056 0.028
R4322 VDD.n1027 VDD.n1025 0.028
R4323 VDD.n1307 VDD.n1304 0.028
R4324 VDD.n1324 VDD.n1322 0.028
R4325 VDD.n1357 VDD.n1354 0.028
R4326 VDD.n239 VDD.n236 0.028
R4327 VDD.n194 VDD.n192 0.028
R4328 VDD.n178 VDD.n175 0.028
R4329 VDD.n2185 VDD.n2184 0.028
R4330 VDD.n2169 VDD.n2167 0.028
R4331 VDD.n2138 VDD.n2136 0.028
R4332 VDD.n484 VDD.n481 0.028
R4333 VDD.n501 VDD.n499 0.028
R4334 VDD.n534 VDD.n531 0.028
R4335 VDD.n1665 VDD.n1662 0.028
R4336 VDD.n1682 VDD.n1680 0.028
R4337 VDD.n1715 VDD.n1712 0.028
R4338 VDD.n1210 VDD.n1207 0.028
R4339 VDD.n1227 VDD.n1225 0.028
R4340 VDD.n1260 VDD.n1257 0.028
R4341 VDD.n2745 VDD.n2744 0.028
R4342 VDD.n2729 VDD.n2727 0.028
R4343 VDD.n2698 VDD.n2696 0.028
R4344 VDD.n2889 VDD.n2886 0.028
R4345 VDD.n2906 VDD.n2904 0.028
R4346 VDD.n2939 VDD.n2936 0.028
R4347 VDD.n3745 VDD.n3743 0.028
R4348 VDD.n3759 VDD.n3758 0.028
R4349 VDD.n3787 VDD.n3785 0.028
R4350 VDD.n3801 VDD.n3800 0.028
R4351 VDD.n3898 VDD.n3896 0.028
R4352 VDD.n3912 VDD.n3911 0.028
R4353 VDD.n3846 VDD.n3844 0.028
R4354 VDD.n3860 VDD.n3859 0.028
R4355 VDD.n4009 VDD.n4007 0.028
R4356 VDD.n4023 VDD.n4022 0.028
R4357 VDD.n3957 VDD.n3955 0.028
R4358 VDD.n3971 VDD.n3970 0.028
R4359 VDD.n4120 VDD.n4118 0.028
R4360 VDD.n4134 VDD.n4133 0.028
R4361 VDD.n4068 VDD.n4066 0.028
R4362 VDD.n4082 VDD.n4081 0.028
R4363 VDD.n4231 VDD.n4229 0.028
R4364 VDD.n4245 VDD.n4244 0.028
R4365 VDD.n4179 VDD.n4177 0.028
R4366 VDD.n4193 VDD.n4192 0.028
R4367 VDD.n4347 VDD.n4345 0.028
R4368 VDD.n4361 VDD.n4360 0.028
R4369 VDD.n4389 VDD.n4387 0.028
R4370 VDD.n4403 VDD.n4402 0.028
R4371 VDD.n4507 VDD.n4505 0.028
R4372 VDD.n4521 VDD.n4520 0.028
R4373 VDD.n4455 VDD.n4453 0.028
R4374 VDD.n4469 VDD.n4468 0.028
R4375 VDD.n4625 VDD.n4623 0.028
R4376 VDD.n4639 VDD.n4638 0.028
R4377 VDD.n4573 VDD.n4571 0.028
R4378 VDD.n4587 VDD.n4586 0.028
R4379 VDD.n4678 VDD.n4676 0.028
R4380 VDD.n4692 VDD.n4691 0.028
R4381 VDD.n15 VDD.n13 0.028
R4382 VDD.n29 VDD.n28 0.028
R4383 VDD.n3427 VDD.n3424 0.027
R4384 VDD.n3071 VDD.n3068 0.027
R4385 VDD.n2791 VDD.n2790 0.026
R4386 VDD.n2785 VDD.n2783 0.026
R4387 VDD.n781 VDD.n780 0.026
R4388 VDD.n775 VDD.n773 0.026
R4389 VDD.n2523 VDD.n2522 0.026
R4390 VDD.n2517 VDD.n2516 0.026
R4391 VDD.n2468 VDD.n2467 0.026
R4392 VDD.n2462 VDD.n2461 0.026
R4393 VDD.n2620 VDD.n2619 0.026
R4394 VDD.n2614 VDD.n2613 0.026
R4395 VDD.n3299 VDD.n3297 0.026
R4396 VDD.n3313 VDD.n3312 0.026
R4397 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/GATE VDD.n3314 0.026
R4398 VDD.n963 VDD.n962 0.026
R4399 VDD.n957 VDD.n955 0.026
R4400 VDD.n1060 VDD.n1059 0.026
R4401 VDD.n1054 VDD.n1053 0.026
R4402 VDD.n1320 VDD.n1318 0.026
R4403 VDD.n1326 VDD.n1325 0.026
R4404 VDD.n1627 VDD.n1626 0.026
R4405 VDD.n1613 VDD.n1611 0.026
R4406 VDD.n1610 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/GATE 0.026
R4407 VDD.n196 VDD.n195 0.026
R4408 VDD.n190 VDD.n188 0.026
R4409 VDD.n2171 VDD.n2170 0.026
R4410 VDD.n2165 VDD.n2164 0.026
R4411 VDD.n497 VDD.n495 0.026
R4412 VDD.n503 VDD.n502 0.026
R4413 VDD.n2127 VDD.n2126 0.026
R4414 VDD.n547 VDD.n546 0.026
R4415 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/GATE VDD.n548 0.026
R4416 VDD.n1678 VDD.n1676 0.026
R4417 VDD.n1684 VDD.n1683 0.026
R4418 VDD.n1223 VDD.n1221 0.026
R4419 VDD.n1229 VDD.n1228 0.026
R4420 VDD.n1728 VDD.n1727 0.026
R4421 VDD.n1273 VDD.n1272 0.026
R4422 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/GATE VDD.n1274 0.026
R4423 VDD.n2731 VDD.n2730 0.026
R4424 VDD.n2725 VDD.n2724 0.026
R4425 VDD.n2902 VDD.n2900 0.026
R4426 VDD.n2908 VDD.n2907 0.026
R4427 VDD.n2687 VDD.n2686 0.026
R4428 VDD.n2952 VDD.n2951 0.026
R4429 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/GATE VDD.n2953 0.026
R4430 VDD.n3740 VDD.n3739 0.026
R4431 VDD.n3782 VDD.n3781 0.026
R4432 VDD.n3893 VDD.n3892 0.026
R4433 VDD.n3841 VDD.n3840 0.026
R4434 VDD.n4004 VDD.n4003 0.026
R4435 VDD.n3952 VDD.n3951 0.026
R4436 VDD.n4115 VDD.n4114 0.026
R4437 VDD.n4063 VDD.n4062 0.026
R4438 VDD.n4226 VDD.n4225 0.026
R4439 VDD.n4174 VDD.n4173 0.026
R4440 VDD.n4342 VDD.n4341 0.026
R4441 VDD.n4384 VDD.n4383 0.026
R4442 VDD.n4502 VDD.n4501 0.026
R4443 VDD.n4450 VDD.n4449 0.026
R4444 VDD.n4620 VDD.n4619 0.026
R4445 VDD.n4568 VDD.n4567 0.026
R4446 VDD.n4673 VDD.n4672 0.026
R4447 VDD.n10 VDD.n9 0.026
R4448 VDD.n2975 VDD.n2974 0.025
R4449 VDD.n2959 VDD.n2958 0.025
R4450 VDD.n3279 VDD.n3277 0.025
R4451 VDD.n3210 VDD.n3208 0.025
R4452 VDD.n3332 VDD.n3330 0.025
R4453 VDD.n3403 VDD.n3401 0.025
R4454 VDD.n1379 VDD.n1377 0.025
R4455 VDD.n1447 VDD.n1445 0.025
R4456 VDD.n1595 VDD.n1593 0.025
R4457 VDD.n1526 VDD.n1524 0.025
R4458 VDD.n438 VDD.n437 0.025
R4459 VDD.n454 VDD.n453 0.025
R4460 VDD.n1998 VDD.n1996 0.025
R4461 VDD.n1930 VDD.n1928 0.025
R4462 VDD.n568 VDD.n566 0.025
R4463 VDD.n639 VDD.n637 0.025
R4464 VDD.n2038 VDD.n2036 0.025
R4465 VDD.n2106 VDD.n2104 0.025
R4466 VDD.n3578 VDD.n3577 0.025
R4467 VDD.n3562 VDD.n3561 0.025
R4468 VDD.n3541 VDD.n3539 0.025
R4469 VDD.n3472 VDD.n3470 0.025
R4470 VDD.n2236 VDD.n2235 0.025
R4471 VDD.n2252 VDD.n2251 0.025
R4472 VDD.n2275 VDD.n2273 0.025
R4473 VDD.n2343 VDD.n2341 0.025
R4474 VDD.n1178 VDD.n1177 0.025
R4475 VDD.n1194 VDD.n1193 0.025
R4476 VDD.n1816 VDD.n1814 0.025
R4477 VDD.n1748 VDD.n1746 0.025
R4478 VDD.n3106 VDD.n3104 0.025
R4479 VDD.n3174 VDD.n3172 0.025
R4480 VDD.n2842 VDD.n2838 0.024
R4481 VDD.n2813 VDD.n2810 0.024
R4482 VDD.n2808 VDD.n2794 0.024
R4483 VDD.n2765 VDD.n2764 0.024
R4484 VDD.n2764 VDD.n2762 0.024
R4485 VDD.n831 VDD.n828 0.024
R4486 VDD.n803 VDD.n800 0.024
R4487 VDD.n798 VDD.n784 0.024
R4488 VDD.n755 VDD.n754 0.024
R4489 VDD.n754 VDD.n752 0.024
R4490 VDD.n2574 VDD.n2571 0.024
R4491 VDD.n2546 VDD.n2543 0.024
R4492 VDD.n2541 VDD.n2526 0.024
R4493 VDD.n2498 VDD.n2497 0.024
R4494 VDD.n2497 VDD.n2495 0.024
R4495 VDD.n2491 VDD.n2490 0.024
R4496 VDD.n2490 VDD.n2487 0.024
R4497 VDD.n2460 VDD.n2457 0.024
R4498 VDD.n2456 VDD.n2454 0.024
R4499 VDD.n2428 VDD.n2426 0.024
R4500 VDD.n2657 VDD.n2656 0.024
R4501 VDD.n2656 VDD.n2652 0.024
R4502 VDD.n2612 VDD.n2609 0.024
R4503 VDD.n2608 VDD.n2606 0.024
R4504 VDD.n2580 VDD.n2416 0.024
R4505 VDD.n1013 VDD.n1010 0.024
R4506 VDD.n985 VDD.n982 0.024
R4507 VDD.n980 VDD.n966 0.024
R4508 VDD.n937 VDD.n936 0.024
R4509 VDD.n936 VDD.n934 0.024
R4510 VDD.n1083 VDD.n1082 0.024
R4511 VDD.n1082 VDD.n1079 0.024
R4512 VDD.n1052 VDD.n1049 0.024
R4513 VDD.n1048 VDD.n1046 0.024
R4514 VDD.n1020 VDD.n1018 0.024
R4515 VDD.n1283 VDD.n930 0.024
R4516 VDD.n1299 VDD.n1283 0.024
R4517 VDD.n1331 VDD.n1329 0.024
R4518 VDD.n1336 VDD.n1333 0.024
R4519 VDD.n1363 VDD.n1361 0.024
R4520 VDD.n247 VDD.n243 0.024
R4521 VDD.n218 VDD.n215 0.024
R4522 VDD.n213 VDD.n199 0.024
R4523 VDD.n170 VDD.n169 0.024
R4524 VDD.n169 VDD.n167 0.024
R4525 VDD.n2195 VDD.n2194 0.024
R4526 VDD.n2194 VDD.n2191 0.024
R4527 VDD.n2163 VDD.n2160 0.024
R4528 VDD.n2159 VDD.n2157 0.024
R4529 VDD.n2131 VDD.n2129 0.024
R4530 VDD.n460 VDD.n251 0.024
R4531 VDD.n476 VDD.n460 0.024
R4532 VDD.n508 VDD.n506 0.024
R4533 VDD.n513 VDD.n510 0.024
R4534 VDD.n540 VDD.n538 0.024
R4535 VDD.n1641 VDD.n925 0.024
R4536 VDD.n1657 VDD.n1641 0.024
R4537 VDD.n1689 VDD.n1687 0.024
R4538 VDD.n1694 VDD.n1691 0.024
R4539 VDD.n1721 VDD.n1719 0.024
R4540 VDD.n1200 VDD.n745 0.024
R4541 VDD.n1202 VDD.n1200 0.024
R4542 VDD.n1234 VDD.n1232 0.024
R4543 VDD.n1239 VDD.n1236 0.024
R4544 VDD.n1266 VDD.n1264 0.024
R4545 VDD.n2755 VDD.n2754 0.024
R4546 VDD.n2754 VDD.n2751 0.024
R4547 VDD.n2723 VDD.n2720 0.024
R4548 VDD.n2719 VDD.n2717 0.024
R4549 VDD.n2691 VDD.n2689 0.024
R4550 VDD.n2865 VDD.n2862 0.024
R4551 VDD.n2881 VDD.n2865 0.024
R4552 VDD.n2913 VDD.n2911 0.024
R4553 VDD.n2918 VDD.n2915 0.024
R4554 VDD.n2945 VDD.n2943 0.024
R4555 VDD.n3733 VDD.n3731 0.024
R4556 VDD.n3758 VDD.n3755 0.024
R4557 VDD.n3775 VDD.n3773 0.024
R4558 VDD.n3800 VDD.n3797 0.024
R4559 VDD.n3886 VDD.n3884 0.024
R4560 VDD.n3911 VDD.n3908 0.024
R4561 VDD.n3834 VDD.n3832 0.024
R4562 VDD.n3859 VDD.n3856 0.024
R4563 VDD.n3997 VDD.n3995 0.024
R4564 VDD.n4022 VDD.n4019 0.024
R4565 VDD.n3945 VDD.n3943 0.024
R4566 VDD.n3970 VDD.n3967 0.024
R4567 VDD.n4108 VDD.n4106 0.024
R4568 VDD.n4133 VDD.n4130 0.024
R4569 VDD.n4056 VDD.n4054 0.024
R4570 VDD.n4081 VDD.n4078 0.024
R4571 VDD.n4219 VDD.n4217 0.024
R4572 VDD.n4244 VDD.n4241 0.024
R4573 VDD.n4167 VDD.n4165 0.024
R4574 VDD.n4192 VDD.n4189 0.024
R4575 VDD.n4335 VDD.n4333 0.024
R4576 VDD.n4360 VDD.n4357 0.024
R4577 VDD.n4377 VDD.n4375 0.024
R4578 VDD.n4402 VDD.n4399 0.024
R4579 VDD.n4495 VDD.n4493 0.024
R4580 VDD.n4520 VDD.n4517 0.024
R4581 VDD.n4443 VDD.n4441 0.024
R4582 VDD.n4468 VDD.n4465 0.024
R4583 VDD.n4613 VDD.n4611 0.024
R4584 VDD.n4638 VDD.n4635 0.024
R4585 VDD.n4561 VDD.n4559 0.024
R4586 VDD.n4586 VDD.n4583 0.024
R4587 VDD.n4666 VDD.n4664 0.024
R4588 VDD.n4691 VDD.n4688 0.024
R4589 VDD.n3 VDD.n1 0.024
R4590 VDD.n28 VDD.n25 0.024
R4591 VDD.n2806 VDD.n2805 0.023
R4592 VDD.n796 VDD.n795 0.023
R4593 VDD.n2538 VDD.n2537 0.023
R4594 VDD.n2642 VDD.n2641 0.023
R4595 VDD.n978 VDD.n977 0.023
R4596 VDD.n1288 VDD.n1287 0.023
R4597 VDD.n211 VDD.n210 0.023
R4598 VDD.n465 VDD.n464 0.023
R4599 VDD.n2207 VDD.n2201 0.023
R4600 VDD.n1646 VDD.n1645 0.023
R4601 VDD.n2870 VDD.n2869 0.023
R4602 VDD.n3433 VDD.n3430 0.022
R4603 VDD.n3078 VDD.n3075 0.022
R4604 VDD.n2978 VDD.n2977 0.021
R4605 VDD.n2956 VDD.n2955 0.021
R4606 VDD.n3291 VDD.n3289 0.021
R4607 VDD.n3198 VDD.n3196 0.021
R4608 VDD.n3320 VDD.n3318 0.021
R4609 VDD.n3415 VDD.n3413 0.021
R4610 VDD.n1367 VDD.n1365 0.021
R4611 VDD.n1459 VDD.n1457 0.021
R4612 VDD.n1607 VDD.n1605 0.021
R4613 VDD.n1514 VDD.n1512 0.021
R4614 VDD.n435 VDD.n434 0.021
R4615 VDD.n457 VDD.n456 0.021
R4616 VDD.n2010 VDD.n2008 0.021
R4617 VDD.n1919 VDD.n1917 0.021
R4618 VDD.n556 VDD.n554 0.021
R4619 VDD.n651 VDD.n649 0.021
R4620 VDD.n2026 VDD.n2024 0.021
R4621 VDD.n2118 VDD.n2116 0.021
R4622 VDD.n3581 VDD.n3580 0.021
R4623 VDD.n3559 VDD.n3558 0.021
R4624 VDD.n3553 VDD.n3551 0.021
R4625 VDD.n3461 VDD.n3459 0.021
R4626 VDD.n2233 VDD.n2232 0.021
R4627 VDD.n2255 VDD.n2254 0.021
R4628 VDD.n2263 VDD.n2261 0.021
R4629 VDD.n2354 VDD.n2352 0.021
R4630 VDD.n1175 VDD.n1174 0.021
R4631 VDD.n1197 VDD.n1196 0.021
R4632 VDD.n1828 VDD.n1826 0.021
R4633 VDD.n1736 VDD.n1734 0.021
R4634 VDD.n3094 VDD.n3092 0.021
R4635 VDD.n3186 VDD.n3184 0.021
R4636 VDD.n3749 VDD.n3748 0.021
R4637 VDD.n3770 VDD.n3767 0.021
R4638 VDD.n3791 VDD.n3790 0.021
R4639 VDD.n3812 VDD.n3809 0.021
R4640 VDD.n3902 VDD.n3901 0.021
R4641 VDD.n3923 VDD.n3920 0.021
R4642 VDD.n3850 VDD.n3849 0.021
R4643 VDD.n3871 VDD.n3868 0.021
R4644 VDD.n4013 VDD.n4012 0.021
R4645 VDD.n4034 VDD.n4031 0.021
R4646 VDD.n3961 VDD.n3960 0.021
R4647 VDD.n3982 VDD.n3979 0.021
R4648 VDD.n4124 VDD.n4123 0.021
R4649 VDD.n4145 VDD.n4142 0.021
R4650 VDD.n4072 VDD.n4071 0.021
R4651 VDD.n4093 VDD.n4090 0.021
R4652 VDD.n4235 VDD.n4234 0.021
R4653 VDD.n4256 VDD.n4253 0.021
R4654 VDD.n4183 VDD.n4182 0.021
R4655 VDD.n4204 VDD.n4201 0.021
R4656 VDD.n4351 VDD.n4350 0.021
R4657 VDD.n4372 VDD.n4369 0.021
R4658 VDD.n4393 VDD.n4392 0.021
R4659 VDD.n4414 VDD.n4411 0.021
R4660 VDD.n4511 VDD.n4510 0.021
R4661 VDD.n4532 VDD.n4529 0.021
R4662 VDD.n4459 VDD.n4458 0.021
R4663 VDD.n4480 VDD.n4477 0.021
R4664 VDD.n4629 VDD.n4628 0.021
R4665 VDD.n4650 VDD.n4647 0.021
R4666 VDD.n4577 VDD.n4576 0.021
R4667 VDD.n4598 VDD.n4595 0.021
R4668 VDD.n4682 VDD.n4681 0.021
R4669 VDD.n4703 VDD.n4700 0.021
R4670 VDD.n19 VDD.n18 0.021
R4671 VDD.n40 VDD.n37 0.021
R4672 VDD.n1851 VDD.n1850 0.02
R4673 VDD.n3315 VDD.n2421 0.019
R4674 VDD.n3295 VDD.n3194 0.019
R4675 VDD.n1609 VDD.n1277 0.019
R4676 VDD.n1633 VDD.n1629 0.019
R4677 VDD.n2860 VDD.n2850 0.019
R4678 VDD.n3614 VDD.n3608 0.018
R4679 VDD.n2838 VDD.n2836 0.016
R4680 VDD.n2810 VDD.n2808 0.016
R4681 VDD.n2774 VDD.n2773 0.016
R4682 VDD.n828 VDD.n826 0.016
R4683 VDD.n800 VDD.n798 0.016
R4684 VDD.n764 VDD.n763 0.016
R4685 VDD.n2571 VDD.n2569 0.016
R4686 VDD.n2543 VDD.n2541 0.016
R4687 VDD.n2507 VDD.n2506 0.016
R4688 VDD.n2480 VDD.n2477 0.016
R4689 VDD.n2457 VDD.n2456 0.016
R4690 VDD.n2430 VDD.n2428 0.016
R4691 VDD.n2632 VDD.n2629 0.016
R4692 VDD.n2609 VDD.n2608 0.016
R4693 VDD.n2582 VDD.n2580 0.016
R4694 VDD.n1010 VDD.n1008 0.016
R4695 VDD.n982 VDD.n980 0.016
R4696 VDD.n946 VDD.n945 0.016
R4697 VDD.n1072 VDD.n1069 0.016
R4698 VDD.n1049 VDD.n1048 0.016
R4699 VDD.n1022 VDD.n1020 0.016
R4700 VDD.n1308 VDD.n1307 0.016
R4701 VDD.n1333 VDD.n1331 0.016
R4702 VDD.n1361 VDD.n1359 0.016
R4703 VDD.n154 VDD.n150 0.016
R4704 VDD.n121 VDD.n114 0.016
R4705 VDD.n121 VDD.n116 0.016
R4706 VDD.n141 VDD.n128 0.016
R4707 VDD.n141 VDD.n140 0.016
R4708 VDD.n137 VDD.n136 0.016
R4709 VDD.n3662 VDD.n3654 0.016
R4710 VDD.n3662 VDD.n3661 0.016
R4711 VDD.n3644 VDD.n3637 0.016
R4712 VDD.n3644 VDD.n3643 0.016
R4713 VDD.n3631 VDD.n159 0.016
R4714 VDD.n243 VDD.n241 0.016
R4715 VDD.n215 VDD.n213 0.016
R4716 VDD.n179 VDD.n178 0.016
R4717 VDD.n2184 VDD.n2181 0.016
R4718 VDD.n2160 VDD.n2159 0.016
R4719 VDD.n2133 VDD.n2131 0.016
R4720 VDD.n485 VDD.n484 0.016
R4721 VDD.n510 VDD.n508 0.016
R4722 VDD.n538 VDD.n536 0.016
R4723 VDD.n902 VDD.n901 0.016
R4724 VDD.n915 VDD.n908 0.016
R4725 VDD.n915 VDD.n914 0.016
R4726 VDD.n887 VDD.n874 0.016
R4727 VDD.n887 VDD.n886 0.016
R4728 VDD.n883 VDD.n882 0.016
R4729 VDD.n868 VDD.n860 0.016
R4730 VDD.n868 VDD.n867 0.016
R4731 VDD.n851 VDD.n844 0.016
R4732 VDD.n851 VDD.n850 0.016
R4733 VDD.n921 VDD.n834 0.016
R4734 VDD.n1666 VDD.n1665 0.016
R4735 VDD.n1691 VDD.n1689 0.016
R4736 VDD.n1719 VDD.n1717 0.016
R4737 VDD.n1211 VDD.n1210 0.016
R4738 VDD.n1236 VDD.n1234 0.016
R4739 VDD.n1264 VDD.n1262 0.016
R4740 VDD.n2744 VDD.n2741 0.016
R4741 VDD.n2720 VDD.n2719 0.016
R4742 VDD.n2693 VDD.n2691 0.016
R4743 VDD.n2890 VDD.n2889 0.016
R4744 VDD.n2915 VDD.n2913 0.016
R4745 VDD.n2943 VDD.n2941 0.016
R4746 VDD.n3674 VDD.n3673 0.016
R4747 VDD.n110 VDD.n103 0.016
R4748 VDD.n110 VDD.n105 0.016
R4749 VDD.n3689 VDD.n3680 0.016
R4750 VDD.n3689 VDD.n3688 0.016
R4751 VDD.n63 VDD.n62 0.016
R4752 VDD.n74 VDD.n66 0.016
R4753 VDD.n74 VDD.n73 0.016
R4754 VDD.n92 VDD.n85 0.016
R4755 VDD.n92 VDD.n91 0.016
R4756 VDD.n2846 VDD.n2845 0.016
R4757 VDD.n3735 VDD.n3733 0.016
R4758 VDD.n3765 VDD.n3763 0.016
R4759 VDD.n3777 VDD.n3775 0.016
R4760 VDD.n3807 VDD.n3805 0.016
R4761 VDD.n3888 VDD.n3886 0.016
R4762 VDD.n3918 VDD.n3916 0.016
R4763 VDD.n3836 VDD.n3834 0.016
R4764 VDD.n3866 VDD.n3864 0.016
R4765 VDD.n3999 VDD.n3997 0.016
R4766 VDD.n4029 VDD.n4027 0.016
R4767 VDD.n3947 VDD.n3945 0.016
R4768 VDD.n3977 VDD.n3975 0.016
R4769 VDD.n4110 VDD.n4108 0.016
R4770 VDD.n4140 VDD.n4138 0.016
R4771 VDD.n4058 VDD.n4056 0.016
R4772 VDD.n4088 VDD.n4086 0.016
R4773 VDD.n4221 VDD.n4219 0.016
R4774 VDD.n4251 VDD.n4249 0.016
R4775 VDD.n4169 VDD.n4167 0.016
R4776 VDD.n4199 VDD.n4197 0.016
R4777 VDD.n4337 VDD.n4335 0.016
R4778 VDD.n4367 VDD.n4365 0.016
R4779 VDD.n4379 VDD.n4377 0.016
R4780 VDD.n4409 VDD.n4407 0.016
R4781 VDD.n4497 VDD.n4495 0.016
R4782 VDD.n4527 VDD.n4525 0.016
R4783 VDD.n4445 VDD.n4443 0.016
R4784 VDD.n4475 VDD.n4473 0.016
R4785 VDD.n4615 VDD.n4613 0.016
R4786 VDD.n4645 VDD.n4643 0.016
R4787 VDD.n4563 VDD.n4561 0.016
R4788 VDD.n4593 VDD.n4591 0.016
R4789 VDD.n4668 VDD.n4666 0.016
R4790 VDD.n4698 VDD.n4696 0.016
R4791 VDD.n5 VDD.n3 0.016
R4792 VDD.n35 VDD.n33 0.016
R4793 VDD.n2977 VDD.n2976 0.015
R4794 VDD.n2957 VDD.n2956 0.015
R4795 VDD.n3289 VDD.n3287 0.015
R4796 VDD.n3206 VDD.n3198 0.015
R4797 VDD.n3328 VDD.n3320 0.015
R4798 VDD.n3413 VDD.n3411 0.015
R4799 VDD.n1375 VDD.n1367 0.015
R4800 VDD.n1457 VDD.n1455 0.015
R4801 VDD.n1605 VDD.n1603 0.015
R4802 VDD.n1522 VDD.n1514 0.015
R4803 VDD.n436 VDD.n435 0.015
R4804 VDD.n456 VDD.n455 0.015
R4805 VDD.n2008 VDD.n2006 0.015
R4806 VDD.n1926 VDD.n1919 0.015
R4807 VDD.n564 VDD.n556 0.015
R4808 VDD.n649 VDD.n647 0.015
R4809 VDD.n2034 VDD.n2026 0.015
R4810 VDD.n2116 VDD.n2114 0.015
R4811 VDD.n3580 VDD.n3579 0.015
R4812 VDD.n3560 VDD.n3559 0.015
R4813 VDD.n3551 VDD.n3549 0.015
R4814 VDD.n3468 VDD.n3461 0.015
R4815 VDD.n2234 VDD.n2233 0.015
R4816 VDD.n2254 VDD.n2253 0.015
R4817 VDD.n2271 VDD.n2263 0.015
R4818 VDD.n2352 VDD.n2350 0.015
R4819 VDD.n1176 VDD.n1175 0.015
R4820 VDD.n1196 VDD.n1195 0.015
R4821 VDD.n1826 VDD.n1824 0.015
R4822 VDD.n1744 VDD.n1736 0.015
R4823 VDD.n3102 VDD.n3094 0.015
R4824 VDD.n3184 VDD.n3182 0.015
R4825 VDD.n3068 VDD.n2850 0.014
R4826 VDD.n2803 VDD.n2802 0.013
R4827 VDD.n2799 VDD.n2798 0.013
R4828 VDD.n793 VDD.n792 0.013
R4829 VDD.n789 VDD.n788 0.013
R4830 VDD.n2535 VDD.n2534 0.013
R4831 VDD.n2531 VDD.n2530 0.013
R4832 VDD.n2649 VDD.n2648 0.013
R4833 VDD.n2645 VDD.n2644 0.013
R4834 VDD.n975 VDD.n974 0.013
R4835 VDD.n971 VDD.n970 0.013
R4836 VDD.n1295 VDD.n1294 0.013
R4837 VDD.n1291 VDD.n1290 0.013
R4838 VDD.n208 VDD.n207 0.013
R4839 VDD.n204 VDD.n203 0.013
R4840 VDD.n472 VDD.n471 0.013
R4841 VDD.n468 VDD.n467 0.013
R4842 VDD.n1653 VDD.n1652 0.013
R4843 VDD.n1649 VDD.n1648 0.013
R4844 VDD.n2877 VDD.n2876 0.013
R4845 VDD.n2873 VDD.n2872 0.013
R4846 VDD.n2831 VDD.n2829 0.012
R4847 VDD.n2794 VDD.n2791 0.012
R4848 VDD.n2787 VDD.n2785 0.012
R4849 VDD.n2777 VDD.n2775 0.012
R4850 VDD.n2775 VDD.n2774 0.012
R4851 VDD.n821 VDD.n819 0.012
R4852 VDD.n784 VDD.n781 0.012
R4853 VDD.n777 VDD.n775 0.012
R4854 VDD.n767 VDD.n765 0.012
R4855 VDD.n765 VDD.n764 0.012
R4856 VDD.n2564 VDD.n2562 0.012
R4857 VDD.n2526 VDD.n2523 0.012
R4858 VDD.n2519 VDD.n2517 0.012
R4859 VDD.n2510 VDD.n2508 0.012
R4860 VDD.n2508 VDD.n2507 0.012
R4861 VDD.n2477 VDD.n2476 0.012
R4862 VDD.n2476 VDD.n2475 0.012
R4863 VDD.n2467 VDD.n2466 0.012
R4864 VDD.n2461 VDD.n2460 0.012
R4865 VDD.n2437 VDD.n2435 0.012
R4866 VDD.n2629 VDD.n2628 0.012
R4867 VDD.n2628 VDD.n2627 0.012
R4868 VDD.n2619 VDD.n2618 0.012
R4869 VDD.n2613 VDD.n2612 0.012
R4870 VDD.n2589 VDD.n2587 0.012
R4871 VDD.n1003 VDD.n1001 0.012
R4872 VDD.n966 VDD.n963 0.012
R4873 VDD.n959 VDD.n957 0.012
R4874 VDD.n949 VDD.n947 0.012
R4875 VDD.n947 VDD.n946 0.012
R4876 VDD.n1069 VDD.n1068 0.012
R4877 VDD.n1068 VDD.n1067 0.012
R4878 VDD.n1059 VDD.n1058 0.012
R4879 VDD.n1053 VDD.n1052 0.012
R4880 VDD.n1029 VDD.n1027 0.012
R4881 VDD.n1310 VDD.n1308 0.012
R4882 VDD.n1312 VDD.n1310 0.012
R4883 VDD.n1322 VDD.n1320 0.012
R4884 VDD.n1329 VDD.n1326 0.012
R4885 VDD.n1354 VDD.n1352 0.012
R4886 VDD.n139 VDD.n138 0.012
R4887 VDD.n3653 VDD.n3652 0.012
R4888 VDD.n236 VDD.n234 0.012
R4889 VDD.n199 VDD.n196 0.012
R4890 VDD.n192 VDD.n190 0.012
R4891 VDD.n182 VDD.n180 0.012
R4892 VDD.n180 VDD.n179 0.012
R4893 VDD.n2181 VDD.n2180 0.012
R4894 VDD.n2180 VDD.n2178 0.012
R4895 VDD.n2170 VDD.n2169 0.012
R4896 VDD.n2164 VDD.n2163 0.012
R4897 VDD.n2140 VDD.n2138 0.012
R4898 VDD.n487 VDD.n485 0.012
R4899 VDD.n489 VDD.n487 0.012
R4900 VDD.n499 VDD.n497 0.012
R4901 VDD.n506 VDD.n503 0.012
R4902 VDD.n531 VDD.n529 0.012
R4903 VDD.n885 VDD.n884 0.012
R4904 VDD.n859 VDD.n858 0.012
R4905 VDD.n1668 VDD.n1666 0.012
R4906 VDD.n1670 VDD.n1668 0.012
R4907 VDD.n1680 VDD.n1678 0.012
R4908 VDD.n1687 VDD.n1684 0.012
R4909 VDD.n1712 VDD.n1710 0.012
R4910 VDD.n1213 VDD.n1211 0.012
R4911 VDD.n1215 VDD.n1213 0.012
R4912 VDD.n1225 VDD.n1223 0.012
R4913 VDD.n1232 VDD.n1229 0.012
R4914 VDD.n1257 VDD.n1255 0.012
R4915 VDD.n2741 VDD.n2740 0.012
R4916 VDD.n2740 VDD.n2738 0.012
R4917 VDD.n2730 VDD.n2729 0.012
R4918 VDD.n2724 VDD.n2723 0.012
R4919 VDD.n2700 VDD.n2698 0.012
R4920 VDD.n2892 VDD.n2890 0.012
R4921 VDD.n2894 VDD.n2892 0.012
R4922 VDD.n2904 VDD.n2902 0.012
R4923 VDD.n2911 VDD.n2908 0.012
R4924 VDD.n2936 VDD.n2934 0.012
R4925 VDD.n3687 VDD.n3686 0.012
R4926 VDD.n65 VDD.n64 0.012
R4927 VDD.n3747 VDD.n3745 0.012
R4928 VDD.n3748 VDD.n3747 0.012
R4929 VDD.n3766 VDD.n3765 0.012
R4930 VDD.n3763 VDD.n3762 0.012
R4931 VDD.n3789 VDD.n3787 0.012
R4932 VDD.n3790 VDD.n3789 0.012
R4933 VDD.n3808 VDD.n3807 0.012
R4934 VDD.n3805 VDD.n3804 0.012
R4935 VDD.n3814 VDD.n3729 0.012
R4936 VDD.n3722 VDD.n3721 0.012
R4937 VDD.n3900 VDD.n3898 0.012
R4938 VDD.n3901 VDD.n3900 0.012
R4939 VDD.n3919 VDD.n3918 0.012
R4940 VDD.n3916 VDD.n3915 0.012
R4941 VDD.n3848 VDD.n3846 0.012
R4942 VDD.n3849 VDD.n3848 0.012
R4943 VDD.n3867 VDD.n3866 0.012
R4944 VDD.n3864 VDD.n3863 0.012
R4945 VDD.n3925 VDD.n3882 0.012
R4946 VDD.n3875 VDD.n3874 0.012
R4947 VDD.n4011 VDD.n4009 0.012
R4948 VDD.n4012 VDD.n4011 0.012
R4949 VDD.n4030 VDD.n4029 0.012
R4950 VDD.n4027 VDD.n4026 0.012
R4951 VDD.n3959 VDD.n3957 0.012
R4952 VDD.n3960 VDD.n3959 0.012
R4953 VDD.n3978 VDD.n3977 0.012
R4954 VDD.n3975 VDD.n3974 0.012
R4955 VDD.n4036 VDD.n3993 0.012
R4956 VDD.n3986 VDD.n3985 0.012
R4957 VDD.n4122 VDD.n4120 0.012
R4958 VDD.n4123 VDD.n4122 0.012
R4959 VDD.n4141 VDD.n4140 0.012
R4960 VDD.n4138 VDD.n4137 0.012
R4961 VDD.n4070 VDD.n4068 0.012
R4962 VDD.n4071 VDD.n4070 0.012
R4963 VDD.n4089 VDD.n4088 0.012
R4964 VDD.n4086 VDD.n4085 0.012
R4965 VDD.n4147 VDD.n4104 0.012
R4966 VDD.n4097 VDD.n4096 0.012
R4967 VDD.n4233 VDD.n4231 0.012
R4968 VDD.n4234 VDD.n4233 0.012
R4969 VDD.n4252 VDD.n4251 0.012
R4970 VDD.n4249 VDD.n4248 0.012
R4971 VDD.n4181 VDD.n4179 0.012
R4972 VDD.n4182 VDD.n4181 0.012
R4973 VDD.n4200 VDD.n4199 0.012
R4974 VDD.n4197 VDD.n4196 0.012
R4975 VDD.n4258 VDD.n4215 0.012
R4976 VDD.n4208 VDD.n4207 0.012
R4977 VDD.n4349 VDD.n4347 0.012
R4978 VDD.n4350 VDD.n4349 0.012
R4979 VDD.n4368 VDD.n4367 0.012
R4980 VDD.n4365 VDD.n4364 0.012
R4981 VDD.n4391 VDD.n4389 0.012
R4982 VDD.n4392 VDD.n4391 0.012
R4983 VDD.n4410 VDD.n4409 0.012
R4984 VDD.n4407 VDD.n4406 0.012
R4985 VDD.n4416 VDD.n4331 0.012
R4986 VDD.n4324 VDD.n4323 0.012
R4987 VDD.n4509 VDD.n4507 0.012
R4988 VDD.n4510 VDD.n4509 0.012
R4989 VDD.n4528 VDD.n4527 0.012
R4990 VDD.n4525 VDD.n4524 0.012
R4991 VDD.n4457 VDD.n4455 0.012
R4992 VDD.n4458 VDD.n4457 0.012
R4993 VDD.n4476 VDD.n4475 0.012
R4994 VDD.n4473 VDD.n4472 0.012
R4995 VDD.n4534 VDD.n4491 0.012
R4996 VDD.n4484 VDD.n4483 0.012
R4997 VDD.n4627 VDD.n4625 0.012
R4998 VDD.n4628 VDD.n4627 0.012
R4999 VDD.n4646 VDD.n4645 0.012
R5000 VDD.n4643 VDD.n4642 0.012
R5001 VDD.n4575 VDD.n4573 0.012
R5002 VDD.n4576 VDD.n4575 0.012
R5003 VDD.n4594 VDD.n4593 0.012
R5004 VDD.n4591 VDD.n4590 0.012
R5005 VDD.n4652 VDD.n4609 0.012
R5006 VDD.n4602 VDD.n4601 0.012
R5007 VDD.n4680 VDD.n4678 0.012
R5008 VDD.n4681 VDD.n4680 0.012
R5009 VDD.n4699 VDD.n4698 0.012
R5010 VDD.n4696 VDD.n4695 0.012
R5011 VDD.n17 VDD.n15 0.012
R5012 VDD.n18 VDD.n17 0.012
R5013 VDD.n36 VDD.n35 0.012
R5014 VDD.n33 VDD.n32 0.012
R5015 VDD.n4706 VDD.n4705 0.012
R5016 VDD.n4714 VDD.n4713 0.012
R5017 VDD.n125 VDD.n124 0.011
R5018 VDD.n853 VDD.n852 0.011
R5019 VDD.n3693 VDD.n3676 0.011
R5020 VDD.n3692 VDD.n3691 0.011
R5021 VDD.n3694 VDD.n3693 0.011
R5022 VDD.n904 VDD.n903 0.011
R5023 VDD.n3664 VDD.n3663 0.011
R5024 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/GATE VDD.n2420 0.011
R5025 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/GATE VDD.n1491 0.011
R5026 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/GATE VDD.n1869 0.011
R5027 VDD.n2861 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/GATE 0.011
R5028 VDD.n3647 VDD.n3633 0.011
R5029 VDD.n3647 VDD.n3646 0.011
R5030 VDD.n3647 VDD.n155 0.011
R5031 VDD.n3647 VDD.n145 0.011
R5032 VDD.n919 VDD.n890 0.011
R5033 VDD.n919 VDD.n918 0.011
R5034 VDD.n919 VDD.n871 0.011
R5035 VDD.n920 VDD.n919 0.011
R5036 VDD.n3693 VDD.n111 0.011
R5037 VDD.n3079 VDD.n3078 0.01
R5038 VDD.n2861 VDD.n2860 0.01
R5039 VDD.n3434 VDD.n3433 0.01
R5040 VDD.n2420 VDD.n2419 0.01
R5041 VDD.n2196 VDD.n1913 0.01
R5042 VDD.n3622 VDD.n3619 0.01
R5043 VDD.n2802 VDD.n2801 0.01
R5044 VDD.n2800 VDD.n2799 0.01
R5045 VDD.n2798 VDD.n2797 0.01
R5046 VDD.n2796 VDD.n2795 0.01
R5047 VDD.n2974 VDD.n2973 0.01
R5048 VDD.n2960 VDD.n2959 0.01
R5049 VDD.n792 VDD.n791 0.01
R5050 VDD.n790 VDD.n789 0.01
R5051 VDD.n788 VDD.n787 0.01
R5052 VDD.n786 VDD.n785 0.01
R5053 VDD.n2534 VDD.n2533 0.01
R5054 VDD.n2532 VDD.n2531 0.01
R5055 VDD.n2530 VDD.n2529 0.01
R5056 VDD.n2528 VDD.n2527 0.01
R5057 VDD.n3295 VDD.n3294 0.01
R5058 VDD.n3277 VDD.n3275 0.01
R5059 VDD.n3219 VDD.n3210 0.01
R5060 VDD.n3438 VDD.n2414 0.01
R5061 VDD.n2651 VDD.n2638 0.01
R5062 VDD.n2650 VDD.n2649 0.01
R5063 VDD.n2648 VDD.n2647 0.01
R5064 VDD.n2646 VDD.n2645 0.01
R5065 VDD.n3316 VDD.n3315 0.01
R5066 VDD.n3340 VDD.n3332 0.01
R5067 VDD.n3401 VDD.n3399 0.01
R5068 VDD.n974 VDD.n973 0.01
R5069 VDD.n972 VDD.n971 0.01
R5070 VDD.n970 VDD.n969 0.01
R5071 VDD.n968 VDD.n967 0.01
R5072 VDD.n1629 VDD.n929 0.01
R5073 VDD.n1387 VDD.n1379 0.01
R5074 VDD.n1445 VDD.n1443 0.01
R5075 VDD.n1297 VDD.n1284 0.01
R5076 VDD.n1296 VDD.n1295 0.01
R5077 VDD.n1294 VDD.n1293 0.01
R5078 VDD.n1292 VDD.n1291 0.01
R5079 VDD.n1609 VDD.n1608 0.01
R5080 VDD.n1593 VDD.n1591 0.01
R5081 VDD.n1534 VDD.n1526 0.01
R5082 VDD.n1510 VDD.n1509 0.01
R5083 VDD.n3608 VDD.n252 0.01
R5084 VDD.n439 VDD.n438 0.01
R5085 VDD.n453 VDD.n452 0.01
R5086 VDD.n1996 VDD.n1994 0.01
R5087 VDD.n1938 VDD.n1930 0.01
R5088 VDD.n576 VDD.n568 0.01
R5089 VDD.n637 VDD.n635 0.01
R5090 VDD.n207 VDD.n206 0.01
R5091 VDD.n205 VDD.n204 0.01
R5092 VDD.n203 VDD.n202 0.01
R5093 VDD.n201 VDD.n200 0.01
R5094 VDD.n474 VDD.n461 0.01
R5095 VDD.n473 VDD.n472 0.01
R5096 VDD.n471 VDD.n470 0.01
R5097 VDD.n469 VDD.n468 0.01
R5098 VDD.n2201 VDD.n1906 0.01
R5099 VDD.n2046 VDD.n2038 0.01
R5100 VDD.n2104 VDD.n2102 0.01
R5101 VDD.n3577 VDD.n3576 0.01
R5102 VDD.n3563 VDD.n3562 0.01
R5103 VDD.n3539 VDD.n3537 0.01
R5104 VDD.n3481 VDD.n3472 0.01
R5105 VDD.n2237 VDD.n2236 0.01
R5106 VDD.n2251 VDD.n2250 0.01
R5107 VDD.n2283 VDD.n2275 0.01
R5108 VDD.n2341 VDD.n2339 0.01
R5109 VDD.n1874 VDD.n744 0.01
R5110 VDD.n1179 VDD.n1178 0.01
R5111 VDD.n1193 VDD.n1192 0.01
R5112 VDD.n1655 VDD.n1642 0.01
R5113 VDD.n1654 VDD.n1653 0.01
R5114 VDD.n1652 VDD.n1651 0.01
R5115 VDD.n1650 VDD.n1649 0.01
R5116 VDD.n1814 VDD.n1812 0.01
R5117 VDD.n1756 VDD.n1748 0.01
R5118 VDD.n2879 VDD.n2866 0.01
R5119 VDD.n2878 VDD.n2877 0.01
R5120 VDD.n2876 VDD.n2875 0.01
R5121 VDD.n2874 VDD.n2873 0.01
R5122 VDD.n3090 VDD.n3084 0.01
R5123 VDD.n3114 VDD.n3106 0.01
R5124 VDD.n3172 VDD.n3170 0.01
R5125 VDD.n4263 VDD.n4262 0.01
R5126 VDD.n4264 VDD.n4263 0.01
R5127 VDD.n4270 VDD.n4269 0.01
R5128 VDD.n4271 VDD.n4270 0.01
R5129 VDD.n4277 VDD.n4276 0.01
R5130 VDD.n4278 VDD.n4277 0.01
R5131 VDD.n4284 VDD.n4283 0.01
R5132 VDD.n4285 VDD.n4284 0.01
R5133 VDD.n4291 VDD.n4290 0.01
R5134 VDD.n4292 VDD.n4291 0.01
R5135 VDD.n4659 VDD.n4658 0.01
R5136 VDD.n4658 VDD.n4657 0.01
R5137 VDD.n4541 VDD.n4540 0.01
R5138 VDD.n4540 VDD.n4539 0.01
R5139 VDD.n4423 VDD.n4422 0.01
R5140 VDD.n4422 VDD.n4421 0.01
R5141 VDD.n4305 VDD.n4304 0.01
R5142 VDD.n4304 VDD.n4303 0.01
R5143 VDD.n124 VDD.n121 0.01
R5144 VDD.n921 VDD.n920 0.01
R5145 VDD.n3691 VDD.n3689 0.01
R5146 VDD.n80 VDD.n74 0.01
R5147 VDD.n93 VDD.n92 0.01
R5148 VDD.n3646 VDD.n3644 0.01
R5149 VDD.n155 VDD.n154 0.01
R5150 VDD.n145 VDD.n141 0.01
R5151 VDD.n890 VDD.n887 0.01
R5152 VDD.n918 VDD.n915 0.01
R5153 VDD.n871 VDD.n868 0.01
R5154 VDD.n852 VDD.n851 0.01
R5155 VDD.n3675 VDD.n3674 0.01
R5156 VDD.n3663 VDD.n3662 0.01
R5157 VDD.n903 VDD.n902 0.01
R5158 VDD.n3633 VDD.n3631 0.01
R5159 VDD.n2846 VDD.n97 0.01
R5160 VDD.n111 VDD.n110 0.01
R5161 VDD.n3706 VDD.n3705 0.009
R5162 VDD.n3817 VDD.n3816 0.009
R5163 VDD.n3928 VDD.n3927 0.009
R5164 VDD.n4039 VDD.n4038 0.009
R5165 VDD.n4150 VDD.n4149 0.009
R5166 VDD.n4308 VDD.n4307 0.009
R5167 VDD.n4426 VDD.n4425 0.009
R5168 VDD.n4544 VDD.n4543 0.009
R5169 VDD.n43 VDD.n42 0.009
R5170 VDD.n2768 VDD.n2766 0.009
R5171 VDD.n758 VDD.n756 0.009
R5172 VDD.n2501 VDD.n2499 0.009
R5173 VDD.n2485 VDD.n2484 0.009
R5174 VDD.n2639 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/SOURCE 0.009
R5175 VDD.n2637 VDD.n2636 0.009
R5176 VDD.n3419 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/GATE 0.009
R5177 VDD.n940 VDD.n938 0.009
R5178 VDD.n1077 VDD.n1076 0.009
R5179 VDD.n1285 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/SOURCE 0.009
R5180 VDD.n1302 VDD.n1300 0.009
R5181 VDD.n1471 VDD.n1469 0.009
R5182 VDD.n173 VDD.n171 0.009
R5183 VDD.n2189 VDD.n2188 0.009
R5184 VDD.n462 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/SOURCE 0.009
R5185 VDD.n479 VDD.n477 0.009
R5186 VDD.n3627 VDD.n3626 0.009
R5187 VDD.n1643 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/SOURCE 0.009
R5188 VDD.n1660 VDD.n1658 0.009
R5189 VDD.n1846 VDD.n1844 0.009
R5190 VDD.n1205 VDD.n1203 0.009
R5191 VDD.n2749 VDD.n2748 0.009
R5192 VDD.n2867 VDD 0.009
R5193 VDD.n2884 VDD.n2882 0.009
R5194 VDD.n3063 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/GATE 0.009
R5195 VDD.n3739 VDD.n3738 0.009
R5196 VDD.n3760 VDD.n3759 0.009
R5197 VDD.n3755 VDD.n3754 0.009
R5198 VDD.n3781 VDD.n3780 0.009
R5199 VDD.n3802 VDD.n3801 0.009
R5200 VDD.n3797 VDD.n3796 0.009
R5201 VDD.n3892 VDD.n3891 0.009
R5202 VDD.n3913 VDD.n3912 0.009
R5203 VDD.n3908 VDD.n3907 0.009
R5204 VDD.n3840 VDD.n3839 0.009
R5205 VDD.n3861 VDD.n3860 0.009
R5206 VDD.n3856 VDD.n3855 0.009
R5207 VDD.n4003 VDD.n4002 0.009
R5208 VDD.n4024 VDD.n4023 0.009
R5209 VDD.n4019 VDD.n4018 0.009
R5210 VDD.n3951 VDD.n3950 0.009
R5211 VDD.n3972 VDD.n3971 0.009
R5212 VDD.n3967 VDD.n3966 0.009
R5213 VDD.n4114 VDD.n4113 0.009
R5214 VDD.n4135 VDD.n4134 0.009
R5215 VDD.n4130 VDD.n4129 0.009
R5216 VDD.n4062 VDD.n4061 0.009
R5217 VDD.n4083 VDD.n4082 0.009
R5218 VDD.n4078 VDD.n4077 0.009
R5219 VDD.n4225 VDD.n4224 0.009
R5220 VDD.n4246 VDD.n4245 0.009
R5221 VDD.n4241 VDD.n4240 0.009
R5222 VDD.n4173 VDD.n4172 0.009
R5223 VDD.n4194 VDD.n4193 0.009
R5224 VDD.n4189 VDD.n4188 0.009
R5225 VDD.n4341 VDD.n4340 0.009
R5226 VDD.n4362 VDD.n4361 0.009
R5227 VDD.n4357 VDD.n4356 0.009
R5228 VDD.n4383 VDD.n4382 0.009
R5229 VDD.n4404 VDD.n4403 0.009
R5230 VDD.n4399 VDD.n4398 0.009
R5231 VDD.n4501 VDD.n4500 0.009
R5232 VDD.n4522 VDD.n4521 0.009
R5233 VDD.n4517 VDD.n4516 0.009
R5234 VDD.n4449 VDD.n4448 0.009
R5235 VDD.n4470 VDD.n4469 0.009
R5236 VDD.n4465 VDD.n4464 0.009
R5237 VDD.n4619 VDD.n4618 0.009
R5238 VDD.n4640 VDD.n4639 0.009
R5239 VDD.n4635 VDD.n4634 0.009
R5240 VDD.n4567 VDD.n4566 0.009
R5241 VDD.n4588 VDD.n4587 0.009
R5242 VDD.n4583 VDD.n4582 0.009
R5243 VDD.n4672 VDD.n4671 0.009
R5244 VDD.n4693 VDD.n4692 0.009
R5245 VDD.n4688 VDD.n4687 0.009
R5246 VDD.n9 VDD.n8 0.009
R5247 VDD.n30 VDD.n29 0.009
R5248 VDD.n25 VDD.n24 0.009
R5249 VDD.n4299 VDD.n3699 0.009
R5250 VDD.n3701 VDD.n3700 0.009
R5251 VDD.n58 VDD.n57 0.008
R5252 VDD.n4299 VDD.n4298 0.008
R5253 VDD.n2804 VDD.n2803 0.008
R5254 VDD.n794 VDD.n793 0.008
R5255 VDD.n2536 VDD.n2535 0.008
R5256 VDD.n2644 VDD.n2643 0.008
R5257 VDD.n2640 VDD.n2639 0.008
R5258 VDD.n3443 VDD.n3438 0.008
R5259 VDD.n976 VDD.n975 0.008
R5260 VDD.n1290 VDD.n1289 0.008
R5261 VDD.n1286 VDD.n1285 0.008
R5262 VDD.n209 VDD.n208 0.008
R5263 VDD.n467 VDD.n466 0.008
R5264 VDD.n463 VDD.n462 0.008
R5265 VDD.n1648 VDD.n1647 0.008
R5266 VDD.n1644 VDD.n1643 0.008
R5267 VDD.n2872 VDD.n2871 0.008
R5268 VDD.n2868 VDD.n2867 0.008
R5269 VDD.n3084 VDD.n2678 0.008
R5270 VDD.n4296 VDD.n3704 0.008
R5271 VDD.n3698 VDD.n58 0.008
R5272 VDD.n3703 VDD.n3701 0.008
R5273 VDD.n3697 VDD.n3696 0.008
R5274 VDD.n4300 VDD.n3698 0.008
R5275 VDD.n4297 VDD.n3703 0.008
R5276 VDD.n4296 VDD.n4295 0.008
R5277 VDD.n1913 VDD.n1912 0.008
R5278 VDD.n2824 VDD.n2822 0.007
R5279 VDD.n2766 VDD.n2765 0.007
R5280 VDD.n814 VDD.n812 0.007
R5281 VDD.n756 VDD.n755 0.007
R5282 VDD.n2557 VDD.n2555 0.007
R5283 VDD.n2499 VDD.n2498 0.007
R5284 VDD.n2487 VDD.n2485 0.007
R5285 VDD.n2444 VDD.n2442 0.007
R5286 VDD.n2652 VDD.n2637 0.007
R5287 VDD.n2596 VDD.n2594 0.007
R5288 VDD.n996 VDD.n994 0.007
R5289 VDD.n938 VDD.n937 0.007
R5290 VDD.n1079 VDD.n1077 0.007
R5291 VDD.n1036 VDD.n1034 0.007
R5292 VDD.n1300 VDD.n1299 0.007
R5293 VDD.n1347 VDD.n1345 0.007
R5294 VDD.n1491 VDD.n1490 0.007
R5295 VDD.n229 VDD.n227 0.007
R5296 VDD.n171 VDD.n170 0.007
R5297 VDD.n2191 VDD.n2189 0.007
R5298 VDD.n2147 VDD.n2145 0.007
R5299 VDD.n477 VDD.n476 0.007
R5300 VDD.n524 VDD.n522 0.007
R5301 VDD.n1658 VDD.n1657 0.007
R5302 VDD.n1705 VDD.n1703 0.007
R5303 VDD.n1869 VDD.n1868 0.007
R5304 VDD.n1203 VDD.n1202 0.007
R5305 VDD.n1250 VDD.n1248 0.007
R5306 VDD.n2751 VDD.n2749 0.007
R5307 VDD.n2707 VDD.n2705 0.007
R5308 VDD.n2882 VDD.n2881 0.007
R5309 VDD.n2929 VDD.n2927 0.007
R5310 VDD.n3736 VDD.n3735 0.007
R5311 VDD.n3767 VDD.n3766 0.007
R5312 VDD.n3778 VDD.n3777 0.007
R5313 VDD.n3809 VDD.n3808 0.007
R5314 VDD.n3716 VDD.n3715 0.007
R5315 VDD.n3720 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/SOURCE 0.007
R5316 VDD.n3889 VDD.n3888 0.007
R5317 VDD.n3920 VDD.n3919 0.007
R5318 VDD.n3837 VDD.n3836 0.007
R5319 VDD.n3868 VDD.n3867 0.007
R5320 VDD.n3827 VDD.n3826 0.007
R5321 VDD.n3873 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/SOURCE 0.007
R5322 VDD.n4000 VDD.n3999 0.007
R5323 VDD.n4031 VDD.n4030 0.007
R5324 VDD.n3948 VDD.n3947 0.007
R5325 VDD.n3979 VDD.n3978 0.007
R5326 VDD.n3938 VDD.n3937 0.007
R5327 VDD.n3984 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/SOURCE 0.007
R5328 VDD.n4111 VDD.n4110 0.007
R5329 VDD.n4142 VDD.n4141 0.007
R5330 VDD.n4059 VDD.n4058 0.007
R5331 VDD.n4090 VDD.n4089 0.007
R5332 VDD.n4049 VDD.n4048 0.007
R5333 VDD.n4095 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/SOURCE 0.007
R5334 VDD.n4222 VDD.n4221 0.007
R5335 VDD.n4253 VDD.n4252 0.007
R5336 VDD.n4170 VDD.n4169 0.007
R5337 VDD.n4201 VDD.n4200 0.007
R5338 VDD.n4160 VDD.n4159 0.007
R5339 VDD.n4206 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/SOURCE 0.007
R5340 VDD.n4338 VDD.n4337 0.007
R5341 VDD.n4369 VDD.n4368 0.007
R5342 VDD.n4380 VDD.n4379 0.007
R5343 VDD.n4411 VDD.n4410 0.007
R5344 VDD.n4318 VDD.n4317 0.007
R5345 VDD.n4322 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/SOURCE 0.007
R5346 VDD.n4498 VDD.n4497 0.007
R5347 VDD.n4529 VDD.n4528 0.007
R5348 VDD.n4446 VDD.n4445 0.007
R5349 VDD.n4477 VDD.n4476 0.007
R5350 VDD.n4436 VDD.n4435 0.007
R5351 VDD.n4482 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/SOURCE 0.007
R5352 VDD.n4616 VDD.n4615 0.007
R5353 VDD.n4647 VDD.n4646 0.007
R5354 VDD.n4564 VDD.n4563 0.007
R5355 VDD.n4595 VDD.n4594 0.007
R5356 VDD.n4554 VDD.n4553 0.007
R5357 VDD.n4600 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/SOURCE 0.007
R5358 VDD.n4669 VDD.n4668 0.007
R5359 VDD.n4700 VDD.n4699 0.007
R5360 VDD.n6 VDD.n5 0.007
R5361 VDD.n37 VDD.n36 0.007
R5362 VDD.n53 VDD.n52 0.007
R5363 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/SOURCE VDD.n4715 0.007
R5364 VDD.n3726 VDD.n3725 0.007
R5365 VDD.n3879 VDD.n3878 0.007
R5366 VDD.n3990 VDD.n3989 0.007
R5367 VDD.n4101 VDD.n4100 0.007
R5368 VDD.n4212 VDD.n4211 0.007
R5369 VDD.n4328 VDD.n4327 0.007
R5370 VDD.n4488 VDD.n4487 0.007
R5371 VDD.n4606 VDD.n4605 0.007
R5372 VDD.n4710 VDD.n4709 0.007
R5373 VDD.n4259 VDD.n4258 0.006
R5374 VDD.n4148 VDD.n4147 0.006
R5375 VDD.n4037 VDD.n4036 0.006
R5376 VDD.n3926 VDD.n3925 0.006
R5377 VDD.n3815 VDD.n3814 0.006
R5378 VDD.n4705 VDD.n4662 0.006
R5379 VDD.n4653 VDD.n4652 0.006
R5380 VDD.n4535 VDD.n4534 0.006
R5381 VDD.n4417 VDD.n4416 0.006
R5382 VDD.n2807 VDD.n2806 0.006
R5383 VDD.n2805 VDD.n2804 0.006
R5384 VDD.n2978 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/BULK 0.006
R5385 VDD.n2971 VDD.n2970 0.006
R5386 VDD.n2963 VDD.n2962 0.006
R5387 VDD.n797 VDD.n796 0.006
R5388 VDD.n795 VDD.n794 0.006
R5389 VDD.n2539 VDD.n2538 0.006
R5390 VDD.n2537 VDD.n2536 0.006
R5391 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/BULK VDD.n3291 0.006
R5392 VDD.n3265 VDD.n3263 0.006
R5393 VDD.n3231 VDD.n3223 0.006
R5394 VDD.n2643 VDD.n2642 0.006
R5395 VDD.n2641 VDD.n2640 0.006
R5396 VDD.n3318 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/BULK 0.006
R5397 VDD.n3353 VDD.n3344 0.006
R5398 VDD.n3389 VDD.n3387 0.006
R5399 VDD.n979 VDD.n978 0.006
R5400 VDD.n977 VDD.n976 0.006
R5401 VDD.n1365 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/BULK 0.006
R5402 VDD.n1399 VDD.n1391 0.006
R5403 VDD.n1433 VDD.n1431 0.006
R5404 VDD.n1289 VDD.n1288 0.006
R5405 VDD.n1287 VDD.n1286 0.006
R5406 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/BULK VDD.n1607 0.006
R5407 VDD.n1581 VDD.n1579 0.006
R5408 VDD.n1546 VDD.n1538 0.006
R5409 VDD.n434 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/BULK 0.006
R5410 VDD.n442 VDD.n441 0.006
R5411 VDD.n450 VDD.n449 0.006
R5412 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/BULK VDD.n2010 0.006
R5413 VDD.n1984 VDD.n1982 0.006
R5414 VDD.n1950 VDD.n1942 0.006
R5415 VDD.n554 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/BULK 0.006
R5416 VDD.n589 VDD.n580 0.006
R5417 VDD.n625 VDD.n623 0.006
R5418 VDD.n212 VDD.n211 0.006
R5419 VDD.n210 VDD.n209 0.006
R5420 VDD.n466 VDD.n465 0.006
R5421 VDD.n464 VDD.n463 0.006
R5422 VDD.n2024 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/BULK 0.006
R5423 VDD.n2058 VDD.n2050 0.006
R5424 VDD.n2092 VDD.n2090 0.006
R5425 VDD.n3619 VDD.n3618 0.006
R5426 VDD.n3581 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/BULK 0.006
R5427 VDD.n3574 VDD.n3573 0.006
R5428 VDD.n3566 VDD.n3565 0.006
R5429 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/BULK VDD.n3553 0.006
R5430 VDD.n3527 VDD.n3525 0.006
R5431 VDD.n3493 VDD.n3485 0.006
R5432 VDD.n2232 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/BULK 0.006
R5433 VDD.n2240 VDD.n2239 0.006
R5434 VDD.n2248 VDD.n2247 0.006
R5435 VDD.n2261 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/BULK 0.006
R5436 VDD.n2295 VDD.n2287 0.006
R5437 VDD.n2329 VDD.n2327 0.006
R5438 VDD.n1174 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/BULK 0.006
R5439 VDD.n1182 VDD.n1181 0.006
R5440 VDD.n1190 VDD.n1189 0.006
R5441 VDD.n1647 VDD.n1646 0.006
R5442 VDD.n1645 VDD.n1644 0.006
R5443 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/BULK VDD.n1828 0.006
R5444 VDD.n1802 VDD.n1800 0.006
R5445 VDD.n1768 VDD.n1760 0.006
R5446 VDD.n2871 VDD.n2870 0.006
R5447 VDD.n2869 VDD.n2868 0.006
R5448 VDD.n3092 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/BULK 0.006
R5449 VDD.n3126 VDD.n3118 0.006
R5450 VDD.n3160 VDD.n3158 0.006
R5451 VDD.n3711 VDD.n3710 0.006
R5452 VDD.n3715 VDD.n3714 0.006
R5453 VDD.n3728 VDD.n3727 0.006
R5454 VDD.n3822 VDD.n3821 0.006
R5455 VDD.n3826 VDD.n3825 0.006
R5456 VDD.n3881 VDD.n3880 0.006
R5457 VDD.n3933 VDD.n3932 0.006
R5458 VDD.n3937 VDD.n3936 0.006
R5459 VDD.n3992 VDD.n3991 0.006
R5460 VDD.n4044 VDD.n4043 0.006
R5461 VDD.n4048 VDD.n4047 0.006
R5462 VDD.n4103 VDD.n4102 0.006
R5463 VDD.n4155 VDD.n4154 0.006
R5464 VDD.n4159 VDD.n4158 0.006
R5465 VDD.n4214 VDD.n4213 0.006
R5466 VDD.n4313 VDD.n4312 0.006
R5467 VDD.n4317 VDD.n4316 0.006
R5468 VDD.n4330 VDD.n4329 0.006
R5469 VDD.n4431 VDD.n4430 0.006
R5470 VDD.n4435 VDD.n4434 0.006
R5471 VDD.n4490 VDD.n4489 0.006
R5472 VDD.n4549 VDD.n4548 0.006
R5473 VDD.n4553 VDD.n4552 0.006
R5474 VDD.n4608 VDD.n4607 0.006
R5475 VDD.n48 VDD.n47 0.006
R5476 VDD.n52 VDD.n51 0.006
R5477 VDD.n4708 VDD.n4707 0.006
R5478 VDD.n3707 VDD.n3706 0.005
R5479 VDD.n3717 VDD.n3716 0.005
R5480 VDD.n3818 VDD.n3817 0.005
R5481 VDD.n3828 VDD.n3827 0.005
R5482 VDD.n3929 VDD.n3928 0.005
R5483 VDD.n3939 VDD.n3938 0.005
R5484 VDD.n4040 VDD.n4039 0.005
R5485 VDD.n4050 VDD.n4049 0.005
R5486 VDD.n4151 VDD.n4150 0.005
R5487 VDD.n4161 VDD.n4160 0.005
R5488 VDD.n4309 VDD.n4308 0.005
R5489 VDD.n4319 VDD.n4318 0.005
R5490 VDD.n4427 VDD.n4426 0.005
R5491 VDD.n4437 VDD.n4436 0.005
R5492 VDD.n4545 VDD.n4544 0.005
R5493 VDD.n4555 VDD.n4554 0.005
R5494 VDD.n44 VDD.n43 0.005
R5495 VDD.n54 VDD.n53 0.005
R5496 VDD.n3725 VDD.n3724 0.004
R5497 VDD.n3878 VDD.n3877 0.004
R5498 VDD.n3989 VDD.n3988 0.004
R5499 VDD.n4100 VDD.n4099 0.004
R5500 VDD.n4211 VDD.n4210 0.004
R5501 VDD.n4327 VDD.n4326 0.004
R5502 VDD.n4487 VDD.n4486 0.004
R5503 VDD.n4605 VDD.n4604 0.004
R5504 VDD.n4711 VDD.n4710 0.004
R5505 VDD.n3667 VDD.n3666 0.004
R5506 VDD.n2795 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/DRAIN 0.004
R5507 VDD.n785 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/DRAIN 0.004
R5508 VDD.n2527 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/DRAIN 0.004
R5509 VDD.n967 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/DRAIN 0.004
R5510 VDD.n1490 VDD.n1487 0.004
R5511 VDD.n200 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/DRAIN 0.004
R5512 VDD.n3618 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/GATE 0.004
R5513 VDD.n1868 VDD.n1864 0.004
R5514 VDD.n3718 VDD.n3717 0.004
R5515 VDD.n3719 VDD.n3718 0.004
R5516 VDD.n3829 VDD.n3828 0.004
R5517 VDD.n3830 VDD.n3829 0.004
R5518 VDD.n3940 VDD.n3939 0.004
R5519 VDD.n3941 VDD.n3940 0.004
R5520 VDD.n4051 VDD.n4050 0.004
R5521 VDD.n4052 VDD.n4051 0.004
R5522 VDD.n4162 VDD.n4161 0.004
R5523 VDD.n4163 VDD.n4162 0.004
R5524 VDD.n4320 VDD.n4319 0.004
R5525 VDD.n4321 VDD.n4320 0.004
R5526 VDD.n4438 VDD.n4437 0.004
R5527 VDD.n4439 VDD.n4438 0.004
R5528 VDD.n4556 VDD.n4555 0.004
R5529 VDD.n4557 VDD.n4556 0.004
R5530 VDD.n55 VDD.n54 0.004
R5531 VDD.n56 VDD.n55 0.004
R5532 VDD.n3815 VDD.n3719 0.003
R5533 VDD.n3926 VDD.n3830 0.003
R5534 VDD.n4037 VDD.n3941 0.003
R5535 VDD.n4148 VDD.n4052 0.003
R5536 VDD.n4259 VDD.n4163 0.003
R5537 VDD.n4417 VDD.n4321 0.003
R5538 VDD.n4535 VDD.n4439 0.003
R5539 VDD.n4653 VDD.n4557 0.003
R5540 VDD.n4662 VDD.n56 0.003
R5541 VDD.n79 VDD.n78 0.003
R5542 VDD.n3695 VDD.n3694 0.003
R5543 VDD.n3692 VDD.n3677 0.003
R5544 VDD.n3665 VDD.n3664 0.003
R5545 VDD.n904 VDD.n894 0.003
R5546 VDD.n3303 VDD.n3299 0.003
R5547 VDD.n3312 VDD.n3310 0.003
R5548 VDD.n1626 VDD.n1624 0.003
R5549 VDD.n1617 VDD.n1613 0.003
R5550 VDD.n155 VDD.n146 0.003
R5551 VDD.n155 VDD.n148 0.003
R5552 VDD.n124 VDD.n112 0.003
R5553 VDD.n124 VDD.n123 0.003
R5554 VDD.n145 VDD.n126 0.003
R5555 VDD.n145 VDD.n144 0.003
R5556 VDD.n143 VDD.n142 0.003
R5557 VDD.n3663 VDD.n3649 0.003
R5558 VDD.n3663 VDD.n3650 0.003
R5559 VDD.n3646 VDD.n3635 0.003
R5560 VDD.n3646 VDD.n3645 0.003
R5561 VDD.n3633 VDD.n157 0.003
R5562 VDD.n3633 VDD.n3632 0.003
R5563 VDD.n2126 VDD.n2124 0.003
R5564 VDD.n546 VDD.n544 0.003
R5565 VDD.n903 VDD.n895 0.003
R5566 VDD.n903 VDD.n896 0.003
R5567 VDD.n918 VDD.n906 0.003
R5568 VDD.n918 VDD.n917 0.003
R5569 VDD.n890 VDD.n872 0.003
R5570 VDD.n890 VDD.n889 0.003
R5571 VDD.n855 VDD.n854 0.003
R5572 VDD.n871 VDD.n856 0.003
R5573 VDD.n871 VDD.n870 0.003
R5574 VDD.n852 VDD.n840 0.003
R5575 VDD.n852 VDD.n842 0.003
R5576 VDD.n920 VDD.n835 0.003
R5577 VDD.n920 VDD.n836 0.003
R5578 VDD.n1727 VDD.n1725 0.003
R5579 VDD.n1272 VDD.n1270 0.003
R5580 VDD.n2686 VDD.n2684 0.003
R5581 VDD.n2951 VDD.n2949 0.003
R5582 VDD.n3675 VDD.n3668 0.003
R5583 VDD.n111 VDD.n99 0.003
R5584 VDD.n111 VDD.n101 0.003
R5585 VDD.n3691 VDD.n3678 0.003
R5586 VDD.n3691 VDD.n3690 0.003
R5587 VDD.n76 VDD.n75 0.003
R5588 VDD.n77 VDD.n76 0.003
R5589 VDD.n81 VDD.n80 0.003
R5590 VDD.n93 VDD.n83 0.003
R5591 VDD.n94 VDD.n93 0.003
R5592 VDD.n97 VDD.n96 0.003
R5593 VDD.n3677 VDD 0.003
R5594 VDD.n3709 VDD.n3708 0.002
R5595 VDD.n3712 VDD.n3711 0.002
R5596 VDD.n3820 VDD.n3819 0.002
R5597 VDD.n3823 VDD.n3822 0.002
R5598 VDD.n3931 VDD.n3930 0.002
R5599 VDD.n3934 VDD.n3933 0.002
R5600 VDD.n4042 VDD.n4041 0.002
R5601 VDD.n4045 VDD.n4044 0.002
R5602 VDD.n4153 VDD.n4152 0.002
R5603 VDD.n4156 VDD.n4155 0.002
R5604 VDD.n4261 VDD.n4260 0.002
R5605 VDD.n4265 VDD.n4264 0.002
R5606 VDD.n4268 VDD.n4267 0.002
R5607 VDD.n4272 VDD.n4271 0.002
R5608 VDD.n4275 VDD.n4274 0.002
R5609 VDD.n4279 VDD.n4278 0.002
R5610 VDD.n4282 VDD.n4281 0.002
R5611 VDD.n4286 VDD.n4285 0.002
R5612 VDD.n4289 VDD.n4288 0.002
R5613 VDD.n4293 VDD.n4292 0.002
R5614 VDD.n4290 VDD.n4289 0.002
R5615 VDD.n4283 VDD.n4282 0.002
R5616 VDD.n4276 VDD.n4275 0.002
R5617 VDD.n4269 VDD.n4268 0.002
R5618 VDD.n4262 VDD.n4261 0.002
R5619 VDD.n4213 VDD.n4212 0.002
R5620 VDD.n4157 VDD.n4156 0.002
R5621 VDD.n4152 VDD.n4151 0.002
R5622 VDD.n4266 VDD.n4265 0.002
R5623 VDD.n4102 VDD.n4101 0.002
R5624 VDD.n4046 VDD.n4045 0.002
R5625 VDD.n4041 VDD.n4040 0.002
R5626 VDD.n4273 VDD.n4272 0.002
R5627 VDD.n3991 VDD.n3990 0.002
R5628 VDD.n3935 VDD.n3934 0.002
R5629 VDD.n3930 VDD.n3929 0.002
R5630 VDD.n4280 VDD.n4279 0.002
R5631 VDD.n3880 VDD.n3879 0.002
R5632 VDD.n3824 VDD.n3823 0.002
R5633 VDD.n3819 VDD.n3818 0.002
R5634 VDD.n4287 VDD.n4286 0.002
R5635 VDD.n3727 VDD.n3726 0.002
R5636 VDD.n3713 VDD.n3712 0.002
R5637 VDD.n3708 VDD.n3707 0.002
R5638 VDD.n4294 VDD.n4293 0.002
R5639 VDD.n4311 VDD.n4310 0.002
R5640 VDD.n4314 VDD.n4313 0.002
R5641 VDD.n4429 VDD.n4428 0.002
R5642 VDD.n4432 VDD.n4431 0.002
R5643 VDD.n4547 VDD.n4546 0.002
R5644 VDD.n4550 VDD.n4549 0.002
R5645 VDD.n46 VDD.n45 0.002
R5646 VDD.n49 VDD.n48 0.002
R5647 VDD.n4661 VDD.n4660 0.002
R5648 VDD.n4657 VDD.n4656 0.002
R5649 VDD.n4654 VDD.n4542 0.002
R5650 VDD.n4539 VDD.n4538 0.002
R5651 VDD.n4536 VDD.n4424 0.002
R5652 VDD.n4421 VDD.n4420 0.002
R5653 VDD.n4418 VDD.n4306 0.002
R5654 VDD.n4303 VDD.n4302 0.002
R5655 VDD.n4306 VDD.n4305 0.002
R5656 VDD.n4424 VDD.n4423 0.002
R5657 VDD.n4542 VDD.n4541 0.002
R5658 VDD.n4660 VDD.n4659 0.002
R5659 VDD.n4709 VDD.n4708 0.002
R5660 VDD.n50 VDD.n49 0.002
R5661 VDD.n45 VDD.n44 0.002
R5662 VDD.n4656 VDD.n4655 0.002
R5663 VDD.n4607 VDD.n4606 0.002
R5664 VDD.n4551 VDD.n4550 0.002
R5665 VDD.n4546 VDD.n4545 0.002
R5666 VDD.n4538 VDD.n4537 0.002
R5667 VDD.n4489 VDD.n4488 0.002
R5668 VDD.n4433 VDD.n4432 0.002
R5669 VDD.n4428 VDD.n4427 0.002
R5670 VDD.n4420 VDD.n4419 0.002
R5671 VDD.n4329 VDD.n4328 0.002
R5672 VDD.n4315 VDD.n4314 0.002
R5673 VDD.n4310 VDD.n4309 0.002
R5674 VDD.n4302 VDD.n4301 0.002
R5675 VDD.n2801 VDD.n2800 0.002
R5676 VDD.n2817 VDD.n2815 0.002
R5677 VDD.n2783 VDD.n2782 0.002
R5678 VDD.n2968 VDD.n2967 0.002
R5679 VDD.n2966 VDD.n2965 0.002
R5680 VDD.n791 VDD.n790 0.002
R5681 VDD.n807 VDD.n805 0.002
R5682 VDD.n773 VDD.n772 0.002
R5683 VDD.n2533 VDD.n2532 0.002
R5684 VDD.n2550 VDD.n2548 0.002
R5685 VDD.n2516 VDD.n2515 0.002
R5686 VDD.n3253 VDD.n3251 0.002
R5687 VDD.n3243 VDD.n3235 0.002
R5688 VDD.n2471 VDD.n2468 0.002
R5689 VDD.n2451 VDD.n2449 0.002
R5690 VDD.n2647 VDD.n2646 0.002
R5691 VDD.n2623 VDD.n2620 0.002
R5692 VDD.n2603 VDD.n2601 0.002
R5693 VDD.n3365 VDD.n3357 0.002
R5694 VDD.n3376 VDD.n3374 0.002
R5695 VDD.n973 VDD.n972 0.002
R5696 VDD.n989 VDD.n987 0.002
R5697 VDD.n955 VDD.n954 0.002
R5698 VDD.n1411 VDD.n1403 0.002
R5699 VDD.n1421 VDD.n1419 0.002
R5700 VDD.n1063 VDD.n1060 0.002
R5701 VDD.n1043 VDD.n1041 0.002
R5702 VDD.n1293 VDD.n1292 0.002
R5703 VDD.n1318 VDD.n1317 0.002
R5704 VDD.n1340 VDD.n1338 0.002
R5705 VDD.n1569 VDD.n1567 0.002
R5706 VDD.n1559 VDD.n1550 0.002
R5707 VDD.n1469 VDD.n1466 0.002
R5708 VDD.n1481 VDD.n1478 0.002
R5709 VDD.n445 VDD.n444 0.002
R5710 VDD.n447 VDD.n446 0.002
R5711 VDD.n1972 VDD.n1970 0.002
R5712 VDD.n1962 VDD.n1954 0.002
R5713 VDD.n601 VDD.n593 0.002
R5714 VDD.n612 VDD.n610 0.002
R5715 VDD.n206 VDD.n205 0.002
R5716 VDD.n222 VDD.n220 0.002
R5717 VDD.n188 VDD.n187 0.002
R5718 VDD.n2174 VDD.n2171 0.002
R5719 VDD.n2154 VDD.n2152 0.002
R5720 VDD.n470 VDD.n469 0.002
R5721 VDD.n495 VDD.n494 0.002
R5722 VDD.n517 VDD.n515 0.002
R5723 VDD.n2070 VDD.n2062 0.002
R5724 VDD.n2080 VDD.n2078 0.002
R5725 VDD.n3627 VDD.n250 0.002
R5726 VDD.n3571 VDD.n3570 0.002
R5727 VDD.n3569 VDD.n3568 0.002
R5728 VDD.n3515 VDD.n3513 0.002
R5729 VDD.n3505 VDD.n3497 0.002
R5730 VDD.n2243 VDD.n2242 0.002
R5731 VDD.n2245 VDD.n2244 0.002
R5732 VDD.n2307 VDD.n2299 0.002
R5733 VDD.n2317 VDD.n2315 0.002
R5734 VDD.n1185 VDD.n1184 0.002
R5735 VDD.n1187 VDD.n1186 0.002
R5736 VDD.n1651 VDD.n1650 0.002
R5737 VDD.n1676 VDD.n1675 0.002
R5738 VDD.n1698 VDD.n1696 0.002
R5739 VDD.n1790 VDD.n1788 0.002
R5740 VDD.n1780 VDD.n1772 0.002
R5741 VDD.n1844 VDD.n1840 0.002
R5742 VDD.n1858 VDD.n1855 0.002
R5743 VDD.n1221 VDD.n1220 0.002
R5744 VDD.n1243 VDD.n1241 0.002
R5745 VDD.n2734 VDD.n2731 0.002
R5746 VDD.n2714 VDD.n2712 0.002
R5747 VDD.n2875 VDD.n2874 0.002
R5748 VDD.n2900 VDD.n2899 0.002
R5749 VDD.n2922 VDD.n2920 0.002
R5750 VDD.n3138 VDD.n3130 0.002
R5751 VDD.n3148 VDD.n3146 0.002
R5752 VDD.n3743 VDD.n3740 0.002
R5753 VDD.n3785 VDD.n3782 0.002
R5754 VDD.n3710 VDD.n3709 0.002
R5755 VDD.n3714 VDD.n3713 0.002
R5756 VDD.n3724 VDD.n3723 0.002
R5757 VDD.n3723 VDD.n3722 0.002
R5758 VDD.n3721 VDD.n3720 0.002
R5759 VDD.n3896 VDD.n3893 0.002
R5760 VDD.n3844 VDD.n3841 0.002
R5761 VDD.n3821 VDD.n3820 0.002
R5762 VDD.n3825 VDD.n3824 0.002
R5763 VDD.n3877 VDD.n3876 0.002
R5764 VDD.n3876 VDD.n3875 0.002
R5765 VDD.n3874 VDD.n3873 0.002
R5766 VDD.n4007 VDD.n4004 0.002
R5767 VDD.n3955 VDD.n3952 0.002
R5768 VDD.n3932 VDD.n3931 0.002
R5769 VDD.n3936 VDD.n3935 0.002
R5770 VDD.n3988 VDD.n3987 0.002
R5771 VDD.n3987 VDD.n3986 0.002
R5772 VDD.n3985 VDD.n3984 0.002
R5773 VDD.n4118 VDD.n4115 0.002
R5774 VDD.n4066 VDD.n4063 0.002
R5775 VDD.n4043 VDD.n4042 0.002
R5776 VDD.n4047 VDD.n4046 0.002
R5777 VDD.n4099 VDD.n4098 0.002
R5778 VDD.n4098 VDD.n4097 0.002
R5779 VDD.n4096 VDD.n4095 0.002
R5780 VDD.n4229 VDD.n4226 0.002
R5781 VDD.n4177 VDD.n4174 0.002
R5782 VDD.n4154 VDD.n4153 0.002
R5783 VDD.n4158 VDD.n4157 0.002
R5784 VDD.n4210 VDD.n4209 0.002
R5785 VDD.n4209 VDD.n4208 0.002
R5786 VDD.n4207 VDD.n4206 0.002
R5787 VDD.n4345 VDD.n4342 0.002
R5788 VDD.n4387 VDD.n4384 0.002
R5789 VDD.n4312 VDD.n4311 0.002
R5790 VDD.n4316 VDD.n4315 0.002
R5791 VDD.n4326 VDD.n4325 0.002
R5792 VDD.n4325 VDD.n4324 0.002
R5793 VDD.n4323 VDD.n4322 0.002
R5794 VDD.n4505 VDD.n4502 0.002
R5795 VDD.n4453 VDD.n4450 0.002
R5796 VDD.n4430 VDD.n4429 0.002
R5797 VDD.n4434 VDD.n4433 0.002
R5798 VDD.n4486 VDD.n4485 0.002
R5799 VDD.n4485 VDD.n4484 0.002
R5800 VDD.n4483 VDD.n4482 0.002
R5801 VDD.n4623 VDD.n4620 0.002
R5802 VDD.n4571 VDD.n4568 0.002
R5803 VDD.n4548 VDD.n4547 0.002
R5804 VDD.n4552 VDD.n4551 0.002
R5805 VDD.n4604 VDD.n4603 0.002
R5806 VDD.n4603 VDD.n4602 0.002
R5807 VDD.n4601 VDD.n4600 0.002
R5808 VDD.n4676 VDD.n4673 0.002
R5809 VDD.n13 VDD.n10 0.002
R5810 VDD.n47 VDD.n46 0.002
R5811 VDD.n51 VDD.n50 0.002
R5812 VDD.n4712 VDD.n4711 0.002
R5813 VDD.n4713 VDD.n4712 0.002
R5814 VDD.n4715 VDD.n4714 0.002
R5815 VDD.n838 VDD.n837 0.002
R5816 VDD.n893 VDD.n892 0.002
R5817 VDD.n839 VDD.n838 0.002
R5818 VDD.n892 VDD.n891 0.002
R5819 VDD.n3631 VDD.n3630 0.002
R5820 VDD.n2847 VDD.n2846 0.002
R5821 VDD.n2797 VDD.n2796 0.001
R5822 VDD.n787 VDD.n786 0.001
R5823 VDD.n2529 VDD.n2528 0.001
R5824 VDD.n2651 VDD.n2650 0.001
R5825 VDD.n3297 VDD.n3296 0.001
R5826 VDD.n3314 VDD.n3313 0.001
R5827 VDD.n969 VDD.n968 0.001
R5828 VDD.n1297 VDD.n1296 0.001
R5829 VDD.n1628 VDD.n1627 0.001
R5830 VDD.n1611 VDD.n1610 0.001
R5831 VDD.n1475 VDD.n1471 0.001
R5832 VDD.n1487 VDD.n1485 0.001
R5833 VDD.n148 VDD.n147 0.001
R5834 VDD.n123 VDD.n122 0.001
R5835 VDD.n144 VDD.n143 0.001
R5836 VDD.n3649 VDD.n3648 0.001
R5837 VDD.n3635 VDD.n3634 0.001
R5838 VDD.n157 VDD.n156 0.001
R5839 VDD.n150 VDD.n149 0.001
R5840 VDD.n114 VDD.n113 0.001
R5841 VDD.n116 VDD.n115 0.001
R5842 VDD.n128 VDD.n127 0.001
R5843 VDD.n140 VDD.n139 0.001
R5844 VDD.n138 VDD.n137 0.001
R5845 VDD.n3652 VDD.n3651 0.001
R5846 VDD.n3654 VDD.n3653 0.001
R5847 VDD.n3661 VDD.n3660 0.001
R5848 VDD.n3637 VDD.n3636 0.001
R5849 VDD.n3643 VDD.n3642 0.001
R5850 VDD.n159 VDD.n158 0.001
R5851 VDD.n202 VDD.n201 0.001
R5852 VDD.n474 VDD.n473 0.001
R5853 VDD.n2127 VDD.n2120 0.001
R5854 VDD.n548 VDD.n547 0.001
R5855 VDD.n906 VDD.n905 0.001
R5856 VDD.n917 VDD.n916 0.001
R5857 VDD.n889 VDD.n888 0.001
R5858 VDD.n856 VDD.n855 0.001
R5859 VDD.n870 VDD.n869 0.001
R5860 VDD.n842 VDD.n841 0.001
R5861 VDD.n901 VDD.n900 0.001
R5862 VDD.n908 VDD.n907 0.001
R5863 VDD.n914 VDD.n913 0.001
R5864 VDD.n874 VDD.n873 0.001
R5865 VDD.n886 VDD.n885 0.001
R5866 VDD.n884 VDD.n883 0.001
R5867 VDD.n858 VDD.n857 0.001
R5868 VDD.n860 VDD.n859 0.001
R5869 VDD.n867 VDD.n866 0.001
R5870 VDD.n844 VDD.n843 0.001
R5871 VDD.n850 VDD.n849 0.001
R5872 VDD.n834 VDD.n833 0.001
R5873 VDD.n1655 VDD.n1654 0.001
R5874 VDD.n1850 VDD.n1846 0.001
R5875 VDD.n1864 VDD.n1862 0.001
R5876 VDD.n1729 VDD.n1728 0.001
R5877 VDD.n1274 VDD.n1273 0.001
R5878 VDD.n2879 VDD.n2878 0.001
R5879 VDD.n2687 VDD.n2660 0.001
R5880 VDD.n2953 VDD.n2952 0.001
R5881 VDD.n3673 VDD.n3672 0.001
R5882 VDD.n103 VDD.n102 0.001
R5883 VDD.n105 VDD.n104 0.001
R5884 VDD.n3680 VDD.n3679 0.001
R5885 VDD.n3688 VDD.n3687 0.001
R5886 VDD.n3686 VDD.n3685 0.001
R5887 VDD.n64 VDD.n63 0.001
R5888 VDD.n66 VDD.n65 0.001
R5889 VDD.n73 VDD.n72 0.001
R5890 VDD.n85 VDD.n84 0.001
R5891 VDD.n91 VDD.n90 0.001
R5892 VDD.n2845 VDD.n2844 0.001
R5893 VDD.n3729 VDD.n3728 0.001
R5894 VDD.n3882 VDD.n3881 0.001
R5895 VDD.n3993 VDD.n3992 0.001
R5896 VDD.n4104 VDD.n4103 0.001
R5897 VDD.n4215 VDD.n4214 0.001
R5898 VDD.n4331 VDD.n4330 0.001
R5899 VDD.n4491 VDD.n4490 0.001
R5900 VDD.n4609 VDD.n4608 0.001
R5901 VDD.n4707 VDD.n4706 0.001
R5902 VDD.n99 VDD.n98 0.001
R5903 VDD.n101 VDD.n100 0.001
R5904 VDD.n78 VDD.n77 0.001
R5905 VDD.n82 VDD.n81 0.001
R5906 VDD.n83 VDD.n82 0.001
R5907 VDD.n95 VDD.n94 0.001
R5908 VDD.n96 VDD.n95 0.001
R5909 VDD.n154 VDD.n153 0.001
R5910 VDD.n922 VDD.n921 0.001
R5911 VDD.n902 VDD.n899 0.001
R5912 VDD.n3674 VDD.n3671 0.001
R5913 VDD.n3693 VDD.n3667 0.001
R5914 VDD.n919 VDD.n904 0.001
R5915 VDD.n3664 VDD.n3647 0.001
R5916 VDD.n3693 VDD.n3692 0.001
R5917 VDD.n80 VDD.n79 0.001
R5918 VDD.n3694 VDD.n97 0.001
R5919 VDD.n3676 VDD.n3675 0.001
R5920 VDD.n919 VDD.n853 0.001
R5921 VDD.n3647 VDD.n125 0.001
R5922 VDD.n853 VDD.n839 0.001
R5923 VDD.n891 VDD.n125 0.001
R5924 IND_CT.n241 IND_CT.n236 9.3
R5925 IND_CT.n265 IND_CT.n264 9.3
R5926 IND_CT.n269 IND_CT.n268 9.3
R5927 IND_CT.n262 IND_CT.n261 9.3
R5928 IND_CT.n247 IND_CT.n246 9.3
R5929 IND_CT.n251 IND_CT.n250 9.3
R5930 IND_CT.n258 IND_CT.n257 9.3
R5931 IND_CT.n239 IND_CT.n238 9.3
R5932 IND_CT.n204 IND_CT.n203 9.3
R5933 IND_CT.n219 IND_CT.n218 9.3
R5934 IND_CT.n223 IND_CT.n222 9.3
R5935 IND_CT.n216 IND_CT.n215 9.3
R5936 IND_CT.n211 IND_CT.n210 9.3
R5937 IND_CT.n195 IND_CT.n190 9.3
R5938 IND_CT.n192 IND_CT.n191 9.3
R5939 IND_CT.n201 IND_CT.n200 9.3
R5940 IND_CT.n133 IND_CT.n128 9.3
R5941 IND_CT.n157 IND_CT.n156 9.3
R5942 IND_CT.n161 IND_CT.n160 9.3
R5943 IND_CT.n154 IND_CT.n153 9.3
R5944 IND_CT.n139 IND_CT.n138 9.3
R5945 IND_CT.n143 IND_CT.n142 9.3
R5946 IND_CT.n150 IND_CT.n149 9.3
R5947 IND_CT.n131 IND_CT.n130 9.3
R5948 IND_CT.n96 IND_CT.n95 9.3
R5949 IND_CT.n111 IND_CT.n110 9.3
R5950 IND_CT.n115 IND_CT.n114 9.3
R5951 IND_CT.n108 IND_CT.n107 9.3
R5952 IND_CT.n103 IND_CT.n102 9.3
R5953 IND_CT.n87 IND_CT.n82 9.3
R5954 IND_CT.n84 IND_CT.n83 9.3
R5955 IND_CT.n93 IND_CT.n92 9.3
R5956 IND_CT.n352 IND_CT.n351 9.3
R5957 IND_CT.n399 IND_CT.n398 9.3
R5958 IND_CT.n404 IND_CT.n403 9.3
R5959 IND_CT.n396 IND_CT.n395 9.3
R5960 IND_CT.n360 IND_CT.n359 9.3
R5961 IND_CT.n363 IND_CT.n362 9.3
R5962 IND_CT.n391 IND_CT.n390 9.3
R5963 IND_CT.n349 IND_CT.n348 9.3
R5964 IND_CT.n439 IND_CT.n438 9.3
R5965 IND_CT.n463 IND_CT.n462 9.3
R5966 IND_CT.n460 IND_CT.n459 9.3
R5967 IND_CT.n452 IND_CT.n451 9.3
R5968 IND_CT.n449 IND_CT.n448 9.3
R5969 IND_CT.n427 IND_CT.n426 9.3
R5970 IND_CT.n431 IND_CT.n430 9.3
R5971 IND_CT.n434 IND_CT.n433 9.3
R5972 IND_CT.n496 IND_CT.n495 9.3
R5973 IND_CT.n543 IND_CT.n542 9.3
R5974 IND_CT.n548 IND_CT.n547 9.3
R5975 IND_CT.n540 IND_CT.n539 9.3
R5976 IND_CT.n504 IND_CT.n503 9.3
R5977 IND_CT.n507 IND_CT.n506 9.3
R5978 IND_CT.n535 IND_CT.n534 9.3
R5979 IND_CT.n493 IND_CT.n492 9.3
R5980 IND_CT.n10 IND_CT.n9 9.3
R5981 IND_CT.n7 IND_CT.n6 9.3
R5982 IND_CT.n15 IND_CT.n14 9.3
R5983 IND_CT.n34 IND_CT.n33 9.3
R5984 IND_CT.n45 IND_CT.n44 9.3
R5985 IND_CT.n42 IND_CT.n41 9.3
R5986 IND_CT.n30 IND_CT.n29 9.3
R5987 IND_CT.n3 IND_CT.n2 9.3
R5988 IND_CT.n233 IND_CT.t3 9.162
R5989 IND_CT.n233 IND_CT.t8 9.162
R5990 IND_CT.n187 IND_CT.t5 9.162
R5991 IND_CT.n187 IND_CT.t14 9.162
R5992 IND_CT.n125 IND_CT.t15 9.162
R5993 IND_CT.n125 IND_CT.t1 9.162
R5994 IND_CT.n79 IND_CT.t6 9.162
R5995 IND_CT.n79 IND_CT.t12 9.162
R5996 IND_CT.n387 IND_CT.t9 9.162
R5997 IND_CT.n387 IND_CT.t11 9.162
R5998 IND_CT.n422 IND_CT.t7 9.162
R5999 IND_CT.n422 IND_CT.t2 9.162
R6000 IND_CT.n531 IND_CT.t4 9.162
R6001 IND_CT.n531 IND_CT.t0 9.162
R6002 IND_CT.n18 IND_CT.t10 9.162
R6003 IND_CT.n18 IND_CT.t13 9.162
R6004 IND_CT.n249 IND_CT.n248 9
R6005 IND_CT.n260 IND_CT.n235 9
R6006 IND_CT.n240 IND_CT.n237 9
R6007 IND_CT.n214 IND_CT.n213 9
R6008 IND_CT.n194 IND_CT.n193 9
R6009 IND_CT.n202 IND_CT.n189 9
R6010 IND_CT.n141 IND_CT.n140 9
R6011 IND_CT.n152 IND_CT.n127 9
R6012 IND_CT.n132 IND_CT.n129 9
R6013 IND_CT.n106 IND_CT.n105 9
R6014 IND_CT.n86 IND_CT.n85 9
R6015 IND_CT.n94 IND_CT.n81 9
R6016 IND_CT.n361 IND_CT.n346 9
R6017 IND_CT.n394 IND_CT.n393 9
R6018 IND_CT.n350 IND_CT.n347 9
R6019 IND_CT.n450 IND_CT.n447 9
R6020 IND_CT.n461 IND_CT.n446 9
R6021 IND_CT.n429 IND_CT.n424 9
R6022 IND_CT.n505 IND_CT.n490 9
R6023 IND_CT.n538 IND_CT.n537 9
R6024 IND_CT.n494 IND_CT.n491 9
R6025 IND_CT.n43 IND_CT.n28 9
R6026 IND_CT.n32 IND_CT.n31 9
R6027 IND_CT.n5 IND_CT.n0 9
R6028 IND_CT.n19 IND_CT.n17 7.474
R6029 IND_CT.n234 IND_CT.n232 7.474
R6030 IND_CT.n188 IND_CT.n186 7.474
R6031 IND_CT.n126 IND_CT.n124 7.474
R6032 IND_CT.n80 IND_CT.n78 7.474
R6033 IND_CT.n388 IND_CT.n386 7.474
R6034 IND_CT.n423 IND_CT.n421 7.474
R6035 IND_CT.n532 IND_CT.n530 7.474
R6036 IND_CT.n234 IND_CT.n233 3.575
R6037 IND_CT.n188 IND_CT.n187 3.575
R6038 IND_CT.n126 IND_CT.n125 3.575
R6039 IND_CT.n80 IND_CT.n79 3.575
R6040 IND_CT.n388 IND_CT.n387 3.575
R6041 IND_CT.n423 IND_CT.n422 3.575
R6042 IND_CT.n532 IND_CT.n531 3.575
R6043 IND_CT.n19 IND_CT.n18 3.575
R6044 IND_CT.n511 IND_CT.n510 2.473
R6045 IND_CT.n367 IND_CT.n366 2.473
R6046 IND_CT.n467 IND_CT.n466 2.473
R6047 IND_CT.n49 IND_CT.n48 2.473
R6048 IND_CT.n272 IND_CT.n271 2.263
R6049 IND_CT.n226 IND_CT.n225 2.263
R6050 IND_CT.n164 IND_CT.n163 2.263
R6051 IND_CT.n118 IND_CT.n117 2.263
R6052 IND_CT.n407 IND_CT.n406 2.261
R6053 IND_CT.n442 IND_CT.n441 2.261
R6054 IND_CT.n551 IND_CT.n550 2.261
R6055 IND_CT.n21 IND_CT.n20 2.261
R6056 IND_CT.n555 IND_CT.n526 1.135
R6057 IND_CT.n483 IND_CT.n482 1.135
R6058 IND_CT.n411 IND_CT.n382 1.135
R6059 IND_CT.n566 IND_CT.n565 1.135
R6060 IND_CT.n324 IND_CT.n323 1.135
R6061 IND_CT.n294 IND_CT.n293 1.135
R6062 IND_CT.n301 IND_CT.n228 1.135
R6063 IND_CT.n331 IND_CT.n120 1.135
R6064 IND_CT.n324 IND_CT.n166 1.135
R6065 IND_CT.n294 IND_CT.n274 1.135
R6066 IND_CT.n555 IND_CT.n554 1.135
R6067 IND_CT.n411 IND_CT.n410 1.135
R6068 IND_CT.n483 IND_CT.n445 1.135
R6069 IND_CT.n53 IND_CT.n52 0.857
R6070 IND_CT.n342 IND_CT.n341 0.849
R6071 IND_CT.n339 IND_CT.n338 0.849
R6072 IND_CT.n336 IND_CT.n335 0.849
R6073 IND_CT.n268 IND_CT.n267 0.189
R6074 IND_CT.n222 IND_CT.n221 0.189
R6075 IND_CT.n160 IND_CT.n159 0.189
R6076 IND_CT.n114 IND_CT.n113 0.189
R6077 IND_CT.n403 IND_CT.n402 0.189
R6078 IND_CT.n438 IND_CT.n437 0.189
R6079 IND_CT.n547 IND_CT.n546 0.189
R6080 IND_CT.n14 IND_CT.n13 0.189
R6081 IND_CT.n257 IND_CT.n256 0.178
R6082 IND_CT.n210 IND_CT.n209 0.178
R6083 IND_CT.n149 IND_CT.n148 0.178
R6084 IND_CT.n102 IND_CT.n101 0.178
R6085 IND_CT.n390 IND_CT.n389 0.178
R6086 IND_CT.n426 IND_CT.n425 0.178
R6087 IND_CT.n534 IND_CT.n533 0.178
R6088 IND_CT.n2 IND_CT.n1 0.178
R6089 IND_CT.n246 IND_CT.n245 0.166
R6090 IND_CT.n200 IND_CT.n199 0.166
R6091 IND_CT.n138 IND_CT.n137 0.166
R6092 IND_CT.n92 IND_CT.n91 0.166
R6093 IND_CT.n359 IND_CT.n358 0.166
R6094 IND_CT.n459 IND_CT.n458 0.166
R6095 IND_CT.n503 IND_CT.n502 0.166
R6096 IND_CT.n41 IND_CT.n40 0.166
R6097 IND_CT.n340 IND_CT.n339 0.15
R6098 IND_CT.n271 IND_CT.n234 0.131
R6099 IND_CT.n225 IND_CT.n188 0.131
R6100 IND_CT.n163 IND_CT.n126 0.131
R6101 IND_CT.n117 IND_CT.n80 0.131
R6102 IND_CT.n406 IND_CT.n388 0.129
R6103 IND_CT.n441 IND_CT.n423 0.129
R6104 IND_CT.n550 IND_CT.n532 0.129
R6105 IND_CT.n20 IND_CT.n19 0.128
R6106 IND_CT.n305 IND_CT.n304 0.12
R6107 IND_CT.n487 IND_CT.n486 0.12
R6108 IND_CT.n55 IND_CT 0.088
R6109 IND_CT.n266 IND_CT.n265 0.062
R6110 IND_CT.n220 IND_CT.n219 0.062
R6111 IND_CT.n158 IND_CT.n157 0.062
R6112 IND_CT.n112 IND_CT.n111 0.062
R6113 IND_CT.n243 IND_CT.n242 0.06
R6114 IND_CT.n197 IND_CT.n196 0.06
R6115 IND_CT.n135 IND_CT.n134 0.06
R6116 IND_CT.n89 IND_CT.n88 0.06
R6117 IND_CT.n400 IND_CT.n399 0.06
R6118 IND_CT.n366 IND_CT.n365 0.06
R6119 IND_CT.n435 IND_CT.n434 0.06
R6120 IND_CT.n466 IND_CT.n465 0.06
R6121 IND_CT.n544 IND_CT.n543 0.06
R6122 IND_CT.n510 IND_CT.n509 0.06
R6123 IND_CT.n11 IND_CT.n10 0.06
R6124 IND_CT.n48 IND_CT.n47 0.06
R6125 IND_CT.n254 IND_CT.n253 0.052
R6126 IND_CT.n207 IND_CT.n206 0.052
R6127 IND_CT.n146 IND_CT.n145 0.052
R6128 IND_CT.n99 IND_CT.n98 0.052
R6129 IND_CT.n355 IND_CT.n354 0.05
R6130 IND_CT.n455 IND_CT.n454 0.05
R6131 IND_CT.n499 IND_CT.n498 0.05
R6132 IND_CT.n37 IND_CT.n36 0.05
R6133 IND_CT.n328 IND_CT.n327 0.045
R6134 IND_CT.n298 IND_CT.n297 0.045
R6135 IND_CT.n415 IND_CT.n414 0.045
R6136 IND_CT.n559 IND_CT.n558 0.045
R6137 IND_CT.n335 IND_CT.n334 0.043
R6138 IND_CT.n343 IND_CT.n342 0.043
R6139 IND_CT.n242 IND_CT.n241 0.038
R6140 IND_CT.n196 IND_CT.n195 0.038
R6141 IND_CT.n134 IND_CT.n133 0.038
R6142 IND_CT.n88 IND_CT.n87 0.038
R6143 IND_CT.n269 IND_CT.n266 0.037
R6144 IND_CT.n223 IND_CT.n220 0.037
R6145 IND_CT.n161 IND_CT.n158 0.037
R6146 IND_CT.n115 IND_CT.n112 0.037
R6147 IND_CT.n258 IND_CT.n255 0.033
R6148 IND_CT.n211 IND_CT.n208 0.033
R6149 IND_CT.n150 IND_CT.n147 0.033
R6150 IND_CT.n103 IND_CT.n100 0.033
R6151 IND_CT.n354 IND_CT.n353 0.031
R6152 IND_CT.n454 IND_CT.n453 0.031
R6153 IND_CT.n498 IND_CT.n497 0.031
R6154 IND_CT.n36 IND_CT.n35 0.031
R6155 IND_CT.n253 IND_CT.n252 0.028
R6156 IND_CT.n249 IND_CT.n247 0.028
R6157 IND_CT.n206 IND_CT.n205 0.028
R6158 IND_CT.n202 IND_CT.n201 0.028
R6159 IND_CT.n145 IND_CT.n144 0.028
R6160 IND_CT.n141 IND_CT.n139 0.028
R6161 IND_CT.n98 IND_CT.n97 0.028
R6162 IND_CT.n94 IND_CT.n93 0.028
R6163 IND_CT.n404 IND_CT.n401 0.028
R6164 IND_CT.n361 IND_CT.n360 0.028
R6165 IND_CT.n439 IND_CT.n436 0.028
R6166 IND_CT.n461 IND_CT.n460 0.028
R6167 IND_CT.n548 IND_CT.n545 0.028
R6168 IND_CT.n505 IND_CT.n504 0.028
R6169 IND_CT.n15 IND_CT.n12 0.028
R6170 IND_CT.n43 IND_CT.n42 0.028
R6171 IND_CT.n357 IND_CT.n356 0.026
R6172 IND_CT.n457 IND_CT.n456 0.026
R6173 IND_CT.n501 IND_CT.n500 0.026
R6174 IND_CT.n39 IND_CT.n38 0.026
R6175 IND_CT.n270 IND_CT.n269 0.024
R6176 IND_CT.n240 IND_CT.n239 0.024
R6177 IND_CT.n224 IND_CT.n223 0.024
R6178 IND_CT.n194 IND_CT.n192 0.024
R6179 IND_CT.n162 IND_CT.n161 0.024
R6180 IND_CT.n132 IND_CT.n131 0.024
R6181 IND_CT.n116 IND_CT.n115 0.024
R6182 IND_CT.n86 IND_CT.n84 0.024
R6183 IND_CT.n405 IND_CT.n404 0.024
R6184 IND_CT.n350 IND_CT.n349 0.024
R6185 IND_CT.n440 IND_CT.n439 0.024
R6186 IND_CT.n450 IND_CT.n449 0.024
R6187 IND_CT.n549 IND_CT.n548 0.024
R6188 IND_CT.n494 IND_CT.n493 0.024
R6189 IND_CT.n16 IND_CT.n15 0.024
R6190 IND_CT.n32 IND_CT.n30 0.024
R6191 IND_CT.n260 IND_CT.n259 0.021
R6192 IND_CT.n214 IND_CT.n212 0.021
R6193 IND_CT.n152 IND_CT.n151 0.021
R6194 IND_CT.n106 IND_CT.n104 0.021
R6195 IND_CT.n392 IND_CT.n391 0.021
R6196 IND_CT.n365 IND_CT.n364 0.021
R6197 IND_CT.n428 IND_CT.n427 0.021
R6198 IND_CT.n465 IND_CT.n464 0.021
R6199 IND_CT.n536 IND_CT.n535 0.021
R6200 IND_CT.n509 IND_CT.n508 0.021
R6201 IND_CT.n4 IND_CT.n3 0.021
R6202 IND_CT.n47 IND_CT.n46 0.021
R6203 IND_CT.n265 IND_CT.n263 0.019
R6204 IND_CT.n219 IND_CT.n217 0.019
R6205 IND_CT.n157 IND_CT.n155 0.019
R6206 IND_CT.n111 IND_CT.n109 0.019
R6207 IND_CT.n247 IND_CT.n244 0.016
R6208 IND_CT.n241 IND_CT.n240 0.016
R6209 IND_CT.n201 IND_CT.n198 0.016
R6210 IND_CT.n195 IND_CT.n194 0.016
R6211 IND_CT.n139 IND_CT.n136 0.016
R6212 IND_CT.n133 IND_CT.n132 0.016
R6213 IND_CT.n93 IND_CT.n90 0.016
R6214 IND_CT.n87 IND_CT.n86 0.016
R6215 IND_CT.n397 IND_CT.n396 0.016
R6216 IND_CT.n352 IND_CT.n350 0.016
R6217 IND_CT.n432 IND_CT.n431 0.016
R6218 IND_CT.n452 IND_CT.n450 0.016
R6219 IND_CT.n541 IND_CT.n540 0.016
R6220 IND_CT.n496 IND_CT.n494 0.016
R6221 IND_CT.n8 IND_CT.n7 0.016
R6222 IND_CT.n34 IND_CT.n32 0.016
R6223 IND_CT.n262 IND_CT.n260 0.012
R6224 IND_CT.n251 IND_CT.n249 0.012
R6225 IND_CT.n244 IND_CT.n243 0.012
R6226 IND_CT.n216 IND_CT.n214 0.012
R6227 IND_CT.n204 IND_CT.n202 0.012
R6228 IND_CT.n198 IND_CT.n197 0.012
R6229 IND_CT.n154 IND_CT.n152 0.012
R6230 IND_CT.n143 IND_CT.n141 0.012
R6231 IND_CT.n136 IND_CT.n135 0.012
R6232 IND_CT.n108 IND_CT.n106 0.012
R6233 IND_CT.n96 IND_CT.n94 0.012
R6234 IND_CT.n90 IND_CT.n89 0.012
R6235 IND_CT.n399 IND_CT.n397 0.012
R6236 IND_CT.n396 IND_CT.n394 0.012
R6237 IND_CT.n364 IND_CT.n363 0.012
R6238 IND_CT.n363 IND_CT.n361 0.012
R6239 IND_CT.n434 IND_CT.n432 0.012
R6240 IND_CT.n431 IND_CT.n429 0.012
R6241 IND_CT.n464 IND_CT.n463 0.012
R6242 IND_CT.n463 IND_CT.n461 0.012
R6243 IND_CT.n543 IND_CT.n541 0.012
R6244 IND_CT.n540 IND_CT.n538 0.012
R6245 IND_CT.n508 IND_CT.n507 0.012
R6246 IND_CT.n507 IND_CT.n505 0.012
R6247 IND_CT.n10 IND_CT.n8 0.012
R6248 IND_CT.n7 IND_CT.n5 0.012
R6249 IND_CT.n46 IND_CT.n45 0.012
R6250 IND_CT.n45 IND_CT.n43 0.012
R6251 IND_CT.n49 IND_CT.n27 0.012
R6252 IND_CT.n287 IND_CT.n286 0.01
R6253 IND_CT.n279 IND_CT.n278 0.01
R6254 IND_CT.n176 IND_CT.n175 0.01
R6255 IND_CT.n168 IND_CT.n167 0.01
R6256 IND_CT.n317 IND_CT.n316 0.01
R6257 IND_CT.n309 IND_CT.n308 0.01
R6258 IND_CT.n68 IND_CT.n67 0.01
R6259 IND_CT.n60 IND_CT.n59 0.01
R6260 IND_CT.n334 IND_CT.n333 0.01
R6261 IND_CT.n329 IND_CT.n328 0.01
R6262 IND_CT.n327 IND_CT.n326 0.01
R6263 IND_CT.n306 IND_CT.n305 0.01
R6264 IND_CT.n304 IND_CT.n303 0.01
R6265 IND_CT.n299 IND_CT.n298 0.01
R6266 IND_CT.n297 IND_CT.n296 0.01
R6267 IND_CT.n276 IND_CT.n275 0.01
R6268 IND_CT.n344 IND_CT.n343 0.01
R6269 IND_CT.n414 IND_CT.n413 0.01
R6270 IND_CT.n416 IND_CT.n415 0.01
R6271 IND_CT.n486 IND_CT.n485 0.01
R6272 IND_CT.n488 IND_CT.n487 0.01
R6273 IND_CT.n558 IND_CT.n557 0.01
R6274 IND_CT.n560 IND_CT.n559 0.01
R6275 IND_CT.n563 IND_CT.n562 0.01
R6276 IND_CT.n369 IND_CT.n368 0.009
R6277 IND_CT.n469 IND_CT.n468 0.009
R6278 IND_CT.n513 IND_CT.n512 0.009
R6279 IND_CT.n580 IND_CT.n579 0.009
R6280 IND_CT.n263 IND_CT.n262 0.009
R6281 IND_CT.n217 IND_CT.n216 0.009
R6282 IND_CT.n183 IND_CT.n182 0.009
R6283 IND_CT.n155 IND_CT.n154 0.009
R6284 IND_CT.n109 IND_CT.n108 0.009
R6285 IND_CT.n75 IND_CT.n74 0.009
R6286 IND_CT.n401 IND_CT.n400 0.009
R6287 IND_CT.n356 IND_CT.n355 0.009
R6288 IND_CT.n436 IND_CT.n435 0.009
R6289 IND_CT.n456 IND_CT.n455 0.009
R6290 IND_CT.n545 IND_CT.n544 0.009
R6291 IND_CT.n500 IND_CT.n499 0.009
R6292 IND_CT.n12 IND_CT.n11 0.009
R6293 IND_CT.n38 IND_CT.n37 0.009
R6294 IND_CT.n181 IND_CT.n180 0.009
R6295 IND_CT.n73 IND_CT.n72 0.009
R6296 IND_CT.n341 IND_CT.n54 0.009
R6297 IND_CT.n335 IND_CT.n58 0.009
R6298 IND_CT.n57 IND_CT.n56 0.009
R6299 IND_CT.n374 IND_CT.n373 0.008
R6300 IND_CT.n518 IND_CT.n517 0.008
R6301 IND_CT.n575 IND_CT.n574 0.008
R6302 IND_CT.n51 IND_CT.n50 0.008
R6303 IND_CT.n56 IND_CT.n55 0.008
R6304 IND_CT.n341 IND_CT.n340 0.008
R6305 IND_CT.n338 IND_CT.n337 0.008
R6306 IND_CT.n53 IND_CT.n51 0.008
R6307 IND_CT.n336 IND_CT.n57 0.008
R6308 IND_CT.n342 IND_CT.n53 0.008
R6309 IND_CT.n339 IND_CT.n336 0.008
R6310 IND_CT.n410 IND_CT.n409 0.008
R6311 IND_CT.n445 IND_CT.n444 0.008
R6312 IND_CT.n554 IND_CT.n553 0.008
R6313 IND_CT.n24 IND_CT.n23 0.008
R6314 IND_CT.n566 IND_CT.n49 0.007
R6315 IND_CT.n526 IND_CT.n511 0.007
R6316 IND_CT.n382 IND_CT.n367 0.007
R6317 IND_CT.n482 IND_CT.n467 0.007
R6318 IND_CT.n259 IND_CT.n258 0.007
R6319 IND_CT.n255 IND_CT.n254 0.007
R6320 IND_CT.n285 IND_CT.n284 0.007
R6321 IND_CT.n212 IND_CT.n211 0.007
R6322 IND_CT.n208 IND_CT.n207 0.007
R6323 IND_CT.n174 IND_CT.n173 0.007
R6324 IND_CT.n151 IND_CT.n150 0.007
R6325 IND_CT.n147 IND_CT.n146 0.007
R6326 IND_CT.n315 IND_CT.n314 0.007
R6327 IND_CT.n104 IND_CT.n103 0.007
R6328 IND_CT.n100 IND_CT.n99 0.007
R6329 IND_CT.n66 IND_CT.n65 0.007
R6330 IND_CT.n394 IND_CT.n392 0.007
R6331 IND_CT.n353 IND_CT.n352 0.007
R6332 IND_CT.n378 IND_CT.n377 0.007
R6333 IND_CT.n429 IND_CT.n428 0.007
R6334 IND_CT.n453 IND_CT.n452 0.007
R6335 IND_CT.n478 IND_CT.n477 0.007
R6336 IND_CT.n538 IND_CT.n536 0.007
R6337 IND_CT.n497 IND_CT.n496 0.007
R6338 IND_CT.n522 IND_CT.n521 0.007
R6339 IND_CT.n5 IND_CT.n4 0.007
R6340 IND_CT.n35 IND_CT.n34 0.007
R6341 IND_CT.n571 IND_CT.n570 0.007
R6342 IND_CT.n323 IND_CT.n322 0.007
R6343 IND_CT.n293 IND_CT.n292 0.007
R6344 IND_CT.n120 IND_CT.n119 0.006
R6345 IND_CT.n166 IND_CT.n165 0.006
R6346 IND_CT.n228 IND_CT.n227 0.006
R6347 IND_CT.n274 IND_CT.n273 0.006
R6348 IND_CT.n274 IND_CT.n231 0.006
R6349 IND_CT.n228 IND_CT.n185 0.006
R6350 IND_CT.n166 IND_CT.n123 0.006
R6351 IND_CT.n120 IND_CT.n77 0.006
R6352 IND_CT.n410 IND_CT.n385 0.006
R6353 IND_CT.n445 IND_CT.n420 0.006
R6354 IND_CT.n554 IND_CT.n529 0.006
R6355 IND_CT.n25 IND_CT.n24 0.006
R6356 IND_CT.n273 IND_CT.n272 0.006
R6357 IND_CT.n289 IND_CT.n288 0.006
R6358 IND_CT.n284 IND_CT.n283 0.006
R6359 IND_CT.n227 IND_CT.n226 0.006
R6360 IND_CT.n178 IND_CT.n177 0.006
R6361 IND_CT.n173 IND_CT.n172 0.006
R6362 IND_CT.n165 IND_CT.n164 0.006
R6363 IND_CT.n319 IND_CT.n318 0.006
R6364 IND_CT.n314 IND_CT.n313 0.006
R6365 IND_CT.n119 IND_CT.n118 0.006
R6366 IND_CT.n70 IND_CT.n69 0.006
R6367 IND_CT.n65 IND_CT.n64 0.006
R6368 IND_CT.n385 IND_CT.n384 0.006
R6369 IND_CT.n377 IND_CT.n376 0.006
R6370 IND_CT.n420 IND_CT.n419 0.006
R6371 IND_CT.n477 IND_CT.n476 0.006
R6372 IND_CT.n474 IND_CT.n473 0.006
R6373 IND_CT.n529 IND_CT.n528 0.006
R6374 IND_CT.n521 IND_CT.n520 0.006
R6375 IND_CT.n26 IND_CT.n25 0.006
R6376 IND_CT.n572 IND_CT.n571 0.006
R6377 IND_CT.n368 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/DRAIN 0.006
R6378 IND_CT.n468 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/DRAIN 0.006
R6379 IND_CT.n512 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/DRAIN 0.006
R6380 IND_CT IND_CT.n580 0.006
R6381 IND_CT.n293 IND_CT.n290 0.005
R6382 IND_CT.n323 IND_CT.n320 0.005
R6383 IND_CT.n283 IND_CT.n282 0.005
R6384 IND_CT.n172 IND_CT.n171 0.005
R6385 IND_CT.n313 IND_CT.n312 0.005
R6386 IND_CT.n64 IND_CT.n63 0.005
R6387 IND_CT.n379 IND_CT.n378 0.005
R6388 IND_CT.n370 IND_CT.n369 0.005
R6389 IND_CT.n479 IND_CT.n478 0.005
R6390 IND_CT.n470 IND_CT.n469 0.005
R6391 IND_CT.n523 IND_CT.n522 0.005
R6392 IND_CT.n514 IND_CT.n513 0.005
R6393 IND_CT.n570 IND_CT.n569 0.005
R6394 IND_CT.n579 IND_CT.n578 0.005
R6395 IND_CT.n252 IND_CT.n251 0.004
R6396 IND_CT.n231 IND_CT.n230 0.004
R6397 IND_CT.n230 IND_CT.n229 0.004
R6398 IND_CT.n278 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/DRAIN 0.004
R6399 IND_CT.n205 IND_CT.n204 0.004
R6400 IND_CT.n185 IND_CT.n184 0.004
R6401 IND_CT.n184 IND_CT.n183 0.004
R6402 IND_CT.n167 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/DRAIN 0.004
R6403 IND_CT.n144 IND_CT.n143 0.004
R6404 IND_CT.n123 IND_CT.n122 0.004
R6405 IND_CT.n122 IND_CT.n121 0.004
R6406 IND_CT.n308 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/DRAIN 0.004
R6407 IND_CT.n97 IND_CT.n96 0.004
R6408 IND_CT.n77 IND_CT.n76 0.004
R6409 IND_CT.n76 IND_CT.n75 0.004
R6410 IND_CT.n59 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/DRAIN 0.004
R6411 IND_CT.n381 IND_CT.n380 0.004
R6412 IND_CT.n380 IND_CT.n379 0.004
R6413 IND_CT.n481 IND_CT.n480 0.004
R6414 IND_CT.n480 IND_CT.n479 0.004
R6415 IND_CT.n475 IND_CT.n474 0.004
R6416 IND_CT.n525 IND_CT.n524 0.004
R6417 IND_CT.n524 IND_CT.n523 0.004
R6418 IND_CT.n568 IND_CT.n567 0.004
R6419 IND_CT.n569 IND_CT.n568 0.004
R6420 IND_CT.n482 IND_CT.n481 0.004
R6421 IND_CT.n567 IND_CT.n566 0.004
R6422 IND_CT.n526 IND_CT.n525 0.004
R6423 IND_CT.n382 IND_CT.n381 0.004
R6424 IND_CT.n288 IND_CT.n287 0.003
R6425 IND_CT.n280 IND_CT.n279 0.003
R6426 IND_CT.n177 IND_CT.n176 0.003
R6427 IND_CT.n169 IND_CT.n168 0.003
R6428 IND_CT.n318 IND_CT.n317 0.003
R6429 IND_CT.n310 IND_CT.n309 0.003
R6430 IND_CT.n69 IND_CT.n68 0.003
R6431 IND_CT.n61 IND_CT.n60 0.003
R6432 IND_CT.n333 IND_CT.n332 0.003
R6433 IND_CT.n330 IND_CT.n329 0.003
R6434 IND_CT.n326 IND_CT.n325 0.003
R6435 IND_CT.n307 IND_CT.n306 0.003
R6436 IND_CT.n303 IND_CT.n302 0.003
R6437 IND_CT.n300 IND_CT.n299 0.003
R6438 IND_CT.n295 IND_CT.n294 0.003
R6439 IND_CT.n277 IND_CT.n276 0.003
R6440 IND_CT.n296 IND_CT.n295 0.003
R6441 IND_CT.n294 IND_CT.n277 0.003
R6442 IND_CT.n301 IND_CT.n300 0.003
R6443 IND_CT.n302 IND_CT.n301 0.003
R6444 IND_CT.n325 IND_CT.n324 0.003
R6445 IND_CT.n331 IND_CT.n330 0.003
R6446 IND_CT.n332 IND_CT.n331 0.003
R6447 IND_CT.n324 IND_CT.n307 0.003
R6448 IND_CT.n411 IND_CT.n345 0.003
R6449 IND_CT.n413 IND_CT.n412 0.003
R6450 IND_CT.n483 IND_CT.n417 0.003
R6451 IND_CT.n485 IND_CT.n484 0.003
R6452 IND_CT.n555 IND_CT.n489 0.003
R6453 IND_CT.n557 IND_CT.n556 0.003
R6454 IND_CT.n565 IND_CT.n561 0.003
R6455 IND_CT.n564 IND_CT.n563 0.003
R6456 IND_CT.n561 IND_CT.n560 0.003
R6457 IND_CT.n556 IND_CT.n555 0.003
R6458 IND_CT.n489 IND_CT.n488 0.003
R6459 IND_CT.n412 IND_CT.n411 0.003
R6460 IND_CT.n345 IND_CT.n344 0.003
R6461 IND_CT.n484 IND_CT.n483 0.003
R6462 IND_CT.n417 IND_CT.n416 0.003
R6463 IND_CT.n565 IND_CT.n564 0.003
R6464 IND_CT.n406 IND_CT.n405 0.003
R6465 IND_CT.n441 IND_CT.n440 0.003
R6466 IND_CT.n550 IND_CT.n549 0.003
R6467 IND_CT.n20 IND_CT.n16 0.003
R6468 IND_CT.n371 IND_CT.n370 0.002
R6469 IND_CT.n471 IND_CT.n470 0.002
R6470 IND_CT.n515 IND_CT.n514 0.002
R6471 IND_CT.n577 IND_CT.n576 0.002
R6472 IND_CT.n578 IND_CT.n577 0.002
R6473 IND_CT.n519 IND_CT.n518 0.002
R6474 IND_CT.n375 IND_CT.n374 0.002
R6475 IND_CT.n372 IND_CT.n371 0.002
R6476 IND_CT.n472 IND_CT.n471 0.002
R6477 IND_CT.n516 IND_CT.n515 0.002
R6478 IND_CT.n574 IND_CT.n573 0.002
R6479 IND_CT.n286 IND_CT.n285 0.002
R6480 IND_CT.n175 IND_CT.n174 0.002
R6481 IND_CT.n316 IND_CT.n315 0.002
R6482 IND_CT.n67 IND_CT.n66 0.002
R6483 IND_CT.n360 IND_CT.n357 0.002
R6484 IND_CT.n408 IND_CT.n407 0.002
R6485 IND_CT.n409 IND_CT.n408 0.002
R6486 IND_CT.n376 IND_CT.n375 0.002
R6487 IND_CT.n373 IND_CT.n372 0.002
R6488 IND_CT.n460 IND_CT.n457 0.002
R6489 IND_CT.n443 IND_CT.n442 0.002
R6490 IND_CT.n444 IND_CT.n443 0.002
R6491 IND_CT.n476 IND_CT.n475 0.002
R6492 IND_CT.n473 IND_CT.n472 0.002
R6493 IND_CT.n504 IND_CT.n501 0.002
R6494 IND_CT.n552 IND_CT.n551 0.002
R6495 IND_CT.n553 IND_CT.n552 0.002
R6496 IND_CT.n520 IND_CT.n519 0.002
R6497 IND_CT.n517 IND_CT.n516 0.002
R6498 IND_CT.n42 IND_CT.n39 0.002
R6499 IND_CT.n22 IND_CT.n21 0.002
R6500 IND_CT.n23 IND_CT.n22 0.002
R6501 IND_CT.n573 IND_CT.n572 0.002
R6502 IND_CT.n576 IND_CT.n575 0.002
R6503 IND_CT.n281 IND_CT.n280 0.002
R6504 IND_CT.n170 IND_CT.n169 0.002
R6505 IND_CT.n311 IND_CT.n310 0.002
R6506 IND_CT.n62 IND_CT.n61 0.002
R6507 IND_CT.n63 IND_CT.n62 0.002
R6508 IND_CT.n312 IND_CT.n311 0.002
R6509 IND_CT.n171 IND_CT.n170 0.002
R6510 IND_CT.n282 IND_CT.n281 0.002
R6511 IND_CT.n72 IND_CT.n71 0.002
R6512 IND_CT.n180 IND_CT.n179 0.002
R6513 IND_CT.n271 IND_CT.n270 0.001
R6514 IND_CT.n225 IND_CT.n224 0.001
R6515 IND_CT.n163 IND_CT.n162 0.001
R6516 IND_CT.n117 IND_CT.n116 0.001
R6517 IND_CT.n292 IND_CT.n291 0.001
R6518 IND_CT.n290 IND_CT.n289 0.001
R6519 IND_CT.n182 IND_CT.n181 0.001
R6520 IND_CT.n179 IND_CT.n178 0.001
R6521 IND_CT.n322 IND_CT.n321 0.001
R6522 IND_CT.n320 IND_CT.n319 0.001
R6523 IND_CT.n74 IND_CT.n73 0.001
R6524 IND_CT.n71 IND_CT.n70 0.001
R6525 IND_CT.n384 IND_CT.n383 0.001
R6526 IND_CT.n419 IND_CT.n418 0.001
R6527 IND_CT.n528 IND_CT.n527 0.001
R6528 IND_CT.n27 IND_CT.n26 0.001
R6529 VBIAS.n78 VBIAS.t0 4.85
R6530 VBIAS.n79 VBIAS.n78 1.137
R6531 VBIAS.n60 VBIAS.n59 1.136
R6532 VBIAS.n30 VBIAS.n29 1.136
R6533 VBIAS.n10 VBIAS.n3 1.136
R6534 VBIAS.n54 VBIAS.n53 0.019
R6535 VBIAS.n78 VBIAS.n71 0.017
R6536 VBIAS.n78 VBIAS.n77 0.015
R6537 VBIAS VBIAS.n80 0.015
R6538 VBIAS.n54 VBIAS.n52 0.011
R6539 VBIAS.n46 VBIAS.n45 0.01
R6540 VBIAS.n27 VBIAS.n26 0.01
R6541 VBIAS.n55 VBIAS.n54 0.008
R6542 VBIAS.n1 VBIAS.n0 0.008
R6543 VBIAS.n45 VBIAS.n44 0.007
R6544 VBIAS.n26 VBIAS.n25 0.007
R6545 VBIAS.n77 VBIAS.n76 0.007
R6546 VBIAS.n44 VBIAS.n43 0.007
R6547 VBIAS.n25 VBIAS.n24 0.007
R6548 VBIAS.n62 VBIAS.n61 0.006
R6549 VBIAS.n2 VBIAS.n1 0.005
R6550 VBIAS.n56 VBIAS.n55 0.005
R6551 VBIAS.n59 VBIAS.n46 0.004
R6552 VBIAS.n40 VBIAS.n39 0.003
R6553 VBIAS.n29 VBIAS.n27 0.003
R6554 VBIAS.n57 VBIAS.n56 0.003
R6555 VBIAS.n3 VBIAS.n2 0.003
R6556 VBIAS.n78 VBIAS.n62 0.003
R6557 VBIAS.n22 VBIAS.n21 0.003
R6558 VBIAS.n73 VBIAS.n72 0.003
R6559 VBIAS.n21 VBIAS.n20 0.003
R6560 VBIAS.n74 VBIAS.n73 0.003
R6561 VBIAS.n70 VBIAS.n69 0.003
R6562 VBIAS.n67 VBIAS.n66 0.002
R6563 VBIAS.n50 VBIAS.n49 0.002
R6564 VBIAS.n66 VBIAS.n65 0.002
R6565 VBIAS.n49 VBIAS.n48 0.002
R6566 VBIAS.n59 VBIAS.n58 0.002
R6567 VBIAS.n10 VBIAS.n9 0.002
R6568 VBIAS.n16 VBIAS.n15 0.002
R6569 VBIAS.n33 VBIAS.n32 0.002
R6570 VBIAS.n34 VBIAS.n33 0.002
R6571 VBIAS.n9 VBIAS.n8 0.002
R6572 VBIAS.n15 VBIAS.n14 0.002
R6573 VBIAS.n8 VBIAS.n7 0.002
R6574 VBIAS.n80 VBIAS.n79 0.002
R6575 VBIAS.n39 VBIAS.n38 0.002
R6576 VBIAS.n29 VBIAS.n28 0.002
R6577 VBIAS.n58 VBIAS.n57 0.002
R6578 VBIAS.n71 VBIAS.n70 0.002
R6579 VBIAS.n19 VBIAS.n18 0.001
R6580 VBIAS.n23 VBIAS.n22 0.001
R6581 VBIAS.n65 VBIAS.n64 0.001
R6582 VBIAS.n69 VBIAS.n68 0.001
R6583 VBIAS.n75 VBIAS.n74 0.001
R6584 VBIAS.n51 VBIAS.n50 0.001
R6585 VBIAS.n48 VBIAS.n47 0.001
R6586 VBIAS.n6 VBIAS.n5 0.001
R6587 VBIAS.n60 VBIAS.n41 0.001
R6588 VBIAS.n41 VBIAS.n40 0.001
R6589 VBIAS.n20 VBIAS.n19 0.001
R6590 VBIAS.n68 VBIAS.n67 0.001
R6591 VBIAS.n5 VBIAS.n4 0.001
R6592 VBIAS.n43 VBIAS.n42 0.001
R6593 VBIAS.n76 VBIAS.n75 0.001
R6594 VBIAS.n52 VBIAS.n51 0.001
R6595 VBIAS.n64 VBIAS.n63 0.001
R6596 VBIAS.n24 VBIAS.n23 0.001
R6597 VBIAS.n32 VBIAS.n31 0.001
R6598 VBIAS.n7 VBIAS.n6 0.001
R6599 VBIAS.n79 VBIAS.n60 0.001
R6600 VBIAS.n12 VBIAS.n11 0.001
R6601 VBIAS.n30 VBIAS.n17 0.001
R6602 VBIAS.n38 VBIAS.n37 0.001
R6603 VBIAS.n17 VBIAS.n16 0.001
R6604 VBIAS.n37 VBIAS.n36 0.001
R6605 VBIAS.n11 VBIAS.n10 0.001
R6606 VBIAS.n31 VBIAS.n30 0.001
R6607 VBIAS.n14 VBIAS.n13 0.001
R6608 VBIAS.n36 VBIAS.n35 0.001
R6609 VBIAS.n35 VBIAS.n34 0.001
R6610 VBIAS.n13 VBIAS.n12 0.001
R6611 GND.n368 GND.n367 195.121
R6612 GND.n360 GND.n359 195.121
R6613 GND.n353 GND.n352 195.121
R6614 GND.n346 GND.n345 195.121
R6615 GND.n339 GND.n338 195.121
R6616 GND.n332 GND.n331 195.121
R6617 GND.n325 GND.n324 195.121
R6618 GND.n318 GND.n317 195.121
R6619 GND.n311 GND.n310 195.121
R6620 GND.n291 GND.n290 195.121
R6621 GND.n284 GND.n283 195.121
R6622 GND.n277 GND.n276 195.121
R6623 GND.n270 GND.n269 195.121
R6624 GND.n263 GND.n262 195.121
R6625 GND.n256 GND.n255 195.121
R6626 GND.n249 GND.n248 195.121
R6627 GND.n242 GND.n241 195.121
R6628 GND.n235 GND.n234 195.121
R6629 GND.n376 GND.n375 146.341
R6630 GND.n228 GND.n227 126.829
R6631 GND.n100 GND.n99 112.571
R6632 GND.n94 GND.n93 112.571
R6633 GND.n89 GND.n88 112.571
R6634 GND.n84 GND.n83 112.571
R6635 GND.n79 GND.n78 112.571
R6636 GND.n74 GND.n73 112.571
R6637 GND.n69 GND.n68 112.571
R6638 GND.n64 GND.n63 112.571
R6639 GND.n59 GND.n58 112.571
R6640 GND.n51 GND.n50 112.571
R6641 GND.n46 GND.n45 112.571
R6642 GND.n41 GND.n40 112.571
R6643 GND.n36 GND.n35 112.571
R6644 GND.n31 GND.n30 112.571
R6645 GND.n26 GND.n25 112.571
R6646 GND.n21 GND.n20 112.571
R6647 GND.n16 GND.n15 112.571
R6648 GND.n11 GND.n10 112.571
R6649 GND.n369 GND.n366 112.571
R6650 GND.n361 GND.n358 112.571
R6651 GND.n354 GND.n351 112.571
R6652 GND.n347 GND.n344 112.571
R6653 GND.n340 GND.n337 112.571
R6654 GND.n333 GND.n330 112.571
R6655 GND.n326 GND.n323 112.571
R6656 GND.n319 GND.n316 112.571
R6657 GND.n312 GND.n309 112.571
R6658 GND.n292 GND.n289 112.571
R6659 GND.n285 GND.n282 112.571
R6660 GND.n278 GND.n275 112.571
R6661 GND.n271 GND.n268 112.571
R6662 GND.n264 GND.n261 112.571
R6663 GND.n257 GND.n254 112.571
R6664 GND.n250 GND.n247 112.571
R6665 GND.n243 GND.n240 112.571
R6666 GND.n236 GND.n233 112.571
R6667 GND.t0 GND.n297 102.439
R6668 GND.n107 GND.n106 84.428
R6669 GND.n377 GND.n374 84.428
R6670 GND.n6 GND.n5 73.171
R6671 GND.n229 GND.n226 73.171
R6672 GND.n142 GND.n133 68.292
R6673 GND.n198 GND.n182 68.292
R6674 GND.n301 GND.n298 59.1
R6675 GND.n302 GND.n296 59.1
R6676 GND.n370 GND.n364 15.058
R6677 GND.n370 GND.n365 15.058
R6678 GND.n362 GND.n357 15.058
R6679 GND.n355 GND.n350 15.058
R6680 GND.n348 GND.n343 15.058
R6681 GND.n341 GND.n336 15.058
R6682 GND.n334 GND.n329 15.058
R6683 GND.n327 GND.n322 15.058
R6684 GND.n320 GND.n315 15.058
R6685 GND.n313 GND.n308 15.058
R6686 GND.n293 GND.n288 15.058
R6687 GND.n286 GND.n281 15.058
R6688 GND.n279 GND.n274 15.058
R6689 GND.n272 GND.n267 15.058
R6690 GND.n265 GND.n260 15.058
R6691 GND.n258 GND.n253 15.058
R6692 GND.n251 GND.n246 15.058
R6693 GND.n244 GND.n239 15.058
R6694 GND.n237 GND.n232 15.058
R6695 GND.n102 GND.n98 15.058
R6696 GND.n102 GND.n101 15.058
R6697 GND.n96 GND.n95 15.058
R6698 GND.n91 GND.n90 15.058
R6699 GND.n86 GND.n85 15.058
R6700 GND.n81 GND.n80 15.058
R6701 GND.n76 GND.n75 15.058
R6702 GND.n71 GND.n70 15.058
R6703 GND.n66 GND.n65 15.058
R6704 GND.n61 GND.n60 15.058
R6705 GND.n53 GND.n52 15.058
R6706 GND.n48 GND.n47 15.058
R6707 GND.n43 GND.n42 15.058
R6708 GND.n38 GND.n37 15.058
R6709 GND.n33 GND.n32 15.058
R6710 GND.n28 GND.n27 15.058
R6711 GND.n23 GND.n22 15.058
R6712 GND.n18 GND.n17 15.058
R6713 GND.n13 GND.n12 15.058
R6714 GND.n142 GND.n126 14.634
R6715 GND.n198 GND.n189 14.634
R6716 GND.n230 GND.n225 9.788
R6717 GND.n8 GND.n7 9.788
R6718 GND.n108 GND.n107 9.3
R6719 GND.n102 GND.n100 9.3
R6720 GND.n96 GND.n94 9.3
R6721 GND.n91 GND.n89 9.3
R6722 GND.n86 GND.n84 9.3
R6723 GND.n81 GND.n79 9.3
R6724 GND.n76 GND.n74 9.3
R6725 GND.n71 GND.n69 9.3
R6726 GND.n66 GND.n64 9.3
R6727 GND.n61 GND.n59 9.3
R6728 GND.n56 GND.n55 9.3
R6729 GND.n53 GND.n51 9.3
R6730 GND.n48 GND.n46 9.3
R6731 GND.n43 GND.n41 9.3
R6732 GND.n38 GND.n36 9.3
R6733 GND.n33 GND.n31 9.3
R6734 GND.n28 GND.n26 9.3
R6735 GND.n23 GND.n21 9.3
R6736 GND.n18 GND.n16 9.3
R6737 GND.n13 GND.n11 9.3
R6738 GND.n8 GND.n6 9.3
R6739 GND.n205 GND.n204 9.3
R6740 GND.n370 GND.n369 9.3
R6741 GND.n369 GND.n368 9.3
R6742 GND.n362 GND.n361 9.3
R6743 GND.n361 GND.n360 9.3
R6744 GND.n355 GND.n354 9.3
R6745 GND.n354 GND.n353 9.3
R6746 GND.n348 GND.n347 9.3
R6747 GND.n347 GND.n346 9.3
R6748 GND.n341 GND.n340 9.3
R6749 GND.n340 GND.n339 9.3
R6750 GND.n334 GND.n333 9.3
R6751 GND.n333 GND.n332 9.3
R6752 GND.n327 GND.n326 9.3
R6753 GND.n326 GND.n325 9.3
R6754 GND.n320 GND.n319 9.3
R6755 GND.n319 GND.n318 9.3
R6756 GND.n313 GND.n312 9.3
R6757 GND.n312 GND.n311 9.3
R6758 GND.n306 GND.n305 9.3
R6759 GND.n305 GND.n304 9.3
R6760 GND.n293 GND.n292 9.3
R6761 GND.n292 GND.n291 9.3
R6762 GND.n286 GND.n285 9.3
R6763 GND.n285 GND.n284 9.3
R6764 GND.n279 GND.n278 9.3
R6765 GND.n278 GND.n277 9.3
R6766 GND.n272 GND.n271 9.3
R6767 GND.n271 GND.n270 9.3
R6768 GND.n265 GND.n264 9.3
R6769 GND.n264 GND.n263 9.3
R6770 GND.n258 GND.n257 9.3
R6771 GND.n257 GND.n256 9.3
R6772 GND.n251 GND.n250 9.3
R6773 GND.n250 GND.n249 9.3
R6774 GND.n244 GND.n243 9.3
R6775 GND.n243 GND.n242 9.3
R6776 GND.n237 GND.n236 9.3
R6777 GND.n236 GND.n235 9.3
R6778 GND.n230 GND.n229 9.3
R6779 GND.n229 GND.n228 9.3
R6780 GND.n378 GND.n377 9.3
R6781 GND.n377 GND.n376 9.3
R6782 GND.n164 GND.n162 9.139
R6783 GND.n160 GND.n158 9.139
R6784 GND.n156 GND.n154 9.139
R6785 GND.n152 GND.n150 9.139
R6786 GND.n148 GND.n125 9.139
R6787 GND.n123 GND.n121 9.139
R6788 GND.n119 GND.n117 9.139
R6789 GND.n115 GND.n113 9.139
R6790 GND.n2 GND.n0 9.139
R6791 GND.n221 GND.n219 9.139
R6792 GND.n172 GND.n170 9.139
R6793 GND.n176 GND.n174 9.139
R6794 GND.n180 GND.n178 9.139
R6795 GND.n209 GND.n207 9.139
R6796 GND.n213 GND.n211 9.139
R6797 GND.n217 GND.n215 9.139
R6798 GND.n168 GND.n167 9.139
R6799 GND.n303 GND.n295 7.905
R6800 GND.n300 GND.n299 7.905
R6801 GND.n306 GND.n303 7.152
R6802 GND.n110 GND.n109 4.916
R6803 GND.n380 GND.n379 4.916
R6804 GND.n4 GND.n3 4.65
R6805 GND.n224 GND.n223 4.65
R6806 GND.n173 GND.n172 3.95
R6807 GND.n177 GND.n176 3.95
R6808 GND.n181 GND.n180 3.95
R6809 GND.n210 GND.n209 3.95
R6810 GND.n214 GND.n213 3.95
R6811 GND.n218 GND.n217 3.95
R6812 GND.n161 GND.n160 3.949
R6813 GND.n157 GND.n156 3.949
R6814 GND.n153 GND.n152 3.949
R6815 GND.n149 GND.n148 3.949
R6816 GND.n124 GND.n123 3.949
R6817 GND.n120 GND.n119 3.949
R6818 GND.n116 GND.n115 3.949
R6819 GND.n206 GND.n205 3.932
R6820 GND.n379 GND.n378 3.764
R6821 GND.n109 GND.n108 3.764
R6822 GND.n103 GND.n102 3.216
R6823 GND.n97 GND.n96 3.216
R6824 GND.n92 GND.n91 3.216
R6825 GND.n87 GND.n86 3.216
R6826 GND.n82 GND.n81 3.216
R6827 GND.n77 GND.n76 3.216
R6828 GND.n72 GND.n71 3.216
R6829 GND.n67 GND.n66 3.216
R6830 GND.n62 GND.n61 3.216
R6831 GND.n57 GND.n56 3.216
R6832 GND.n54 GND.n53 3.216
R6833 GND.n49 GND.n48 3.216
R6834 GND.n44 GND.n43 3.216
R6835 GND.n39 GND.n38 3.216
R6836 GND.n34 GND.n33 3.216
R6837 GND.n29 GND.n28 3.216
R6838 GND.n24 GND.n23 3.216
R6839 GND.n19 GND.n18 3.216
R6840 GND.n14 GND.n13 3.216
R6841 GND.n9 GND.n8 3.216
R6842 GND.n371 GND.n370 3.216
R6843 GND.n363 GND.n362 3.216
R6844 GND.n356 GND.n355 3.216
R6845 GND.n349 GND.n348 3.216
R6846 GND.n342 GND.n341 3.216
R6847 GND.n335 GND.n334 3.216
R6848 GND.n328 GND.n327 3.216
R6849 GND.n321 GND.n320 3.216
R6850 GND.n314 GND.n313 3.216
R6851 GND.n307 GND.n306 3.216
R6852 GND.n294 GND.n293 3.216
R6853 GND.n287 GND.n286 3.216
R6854 GND.n280 GND.n279 3.216
R6855 GND.n273 GND.n272 3.216
R6856 GND.n266 GND.n265 3.216
R6857 GND.n259 GND.n258 3.216
R6858 GND.n252 GND.n251 3.216
R6859 GND.n245 GND.n244 3.216
R6860 GND.n238 GND.n237 3.216
R6861 GND.n231 GND.n230 3.216
R6862 GND.n165 GND.n164 3.114
R6863 GND.n222 GND.n221 3.114
R6864 GND.n169 GND.n168 3.114
R6865 GND.n112 GND.n2 3.114
R6866 GND.n379 GND.n373 2.635
R6867 GND.n109 GND.n105 2.635
R6868 GND.n128 GND.n127 2.25
R6869 GND.n142 GND.n128 2.25
R6870 GND.n139 GND.n138 2.25
R6871 GND.n142 GND.n139 2.25
R6872 GND.n130 GND.n129 2.25
R6873 GND.n142 GND.n130 2.25
R6874 GND.n144 GND.n143 2.25
R6875 GND.n137 GND.n136 2.25
R6876 GND.n142 GND.n137 2.25
R6877 GND.n132 GND.n131 2.25
R6878 GND.n142 GND.n132 2.25
R6879 GND.n135 GND.n134 2.25
R6880 GND.n142 GND.n135 2.25
R6881 GND.n191 GND.n190 2.25
R6882 GND.n198 GND.n191 2.25
R6883 GND.n188 GND.n187 2.25
R6884 GND.n198 GND.n188 2.25
R6885 GND.n193 GND.n192 2.25
R6886 GND.n198 GND.n193 2.25
R6887 GND.n200 GND.n199 2.25
R6888 GND.n186 GND.n185 2.25
R6889 GND.n198 GND.n186 2.25
R6890 GND.n195 GND.n194 2.25
R6891 GND.n198 GND.n195 2.25
R6892 GND.n184 GND.n183 2.25
R6893 GND.n198 GND.n184 2.25
R6894 GND.n197 GND.n196 2.25
R6895 GND.n198 GND.n197 2.25
R6896 GND.n141 GND.n140 2.25
R6897 GND.n142 GND.n141 2.25
R6898 GND.n145 GND.n144 2.201
R6899 GND.n201 GND.n200 2.201
R6900 GND.n205 GND.n203 1.129
R6901 GND.n172 GND.n171 1.11
R6902 GND.n176 GND.n175 1.11
R6903 GND.n180 GND.n179 1.11
R6904 GND.n209 GND.n208 1.11
R6905 GND.n213 GND.n212 1.11
R6906 GND.n217 GND.n216 1.11
R6907 GND.n221 GND.n220 1.11
R6908 GND.n164 GND.n163 1.11
R6909 GND.n160 GND.n159 1.11
R6910 GND.n156 GND.n155 1.11
R6911 GND.n152 GND.n151 1.11
R6912 GND.n148 GND.n147 1.11
R6913 GND.n123 GND.n122 1.11
R6914 GND.n119 GND.n118 1.11
R6915 GND.n115 GND.n114 1.11
R6916 GND.n168 GND.n166 1.11
R6917 GND.n2 GND.n1 1.11
R6918 GND.n112 GND.n111 0.265
R6919 GND.n224 GND.n222 0.21
R6920 GND GND.n165 0.16
R6921 GND.n120 GND.n116 0.142
R6922 GND.n124 GND.n120 0.142
R6923 GND.n149 GND.n124 0.142
R6924 GND.n153 GND.n149 0.142
R6925 GND.n157 GND.n153 0.142
R6926 GND.n161 GND.n157 0.142
R6927 GND.n103 GND.n97 0.142
R6928 GND.n97 GND.n92 0.142
R6929 GND.n92 GND.n87 0.142
R6930 GND.n87 GND.n82 0.142
R6931 GND.n82 GND.n77 0.142
R6932 GND.n77 GND.n72 0.142
R6933 GND.n72 GND.n67 0.142
R6934 GND.n67 GND.n62 0.142
R6935 GND.n62 GND.n57 0.142
R6936 GND.n57 GND.n54 0.142
R6937 GND.n54 GND.n49 0.142
R6938 GND.n49 GND.n44 0.142
R6939 GND.n44 GND.n39 0.142
R6940 GND.n39 GND.n34 0.142
R6941 GND.n34 GND.n29 0.142
R6942 GND.n29 GND.n24 0.142
R6943 GND.n24 GND.n19 0.142
R6944 GND.n19 GND.n14 0.142
R6945 GND.n14 GND.n9 0.142
R6946 GND.n9 GND.n4 0.142
R6947 GND.n177 GND.n173 0.142
R6948 GND.n181 GND.n177 0.142
R6949 GND.n206 GND.n181 0.142
R6950 GND.n210 GND.n206 0.142
R6951 GND.n214 GND.n210 0.142
R6952 GND.n218 GND.n214 0.142
R6953 GND.n371 GND.n363 0.142
R6954 GND.n363 GND.n356 0.142
R6955 GND.n356 GND.n349 0.142
R6956 GND.n349 GND.n342 0.142
R6957 GND.n342 GND.n335 0.142
R6958 GND.n335 GND.n328 0.142
R6959 GND.n328 GND.n321 0.142
R6960 GND.n321 GND.n314 0.142
R6961 GND.n314 GND.n307 0.142
R6962 GND.n307 GND.n294 0.142
R6963 GND.n294 GND.n287 0.142
R6964 GND.n287 GND.n280 0.142
R6965 GND.n280 GND.n273 0.142
R6966 GND.n273 GND.n266 0.142
R6967 GND.n266 GND.n259 0.142
R6968 GND.n259 GND.n252 0.142
R6969 GND.n252 GND.n245 0.142
R6970 GND.n245 GND.n238 0.142
R6971 GND.n238 GND.n231 0.142
R6972 GND.n231 GND.n224 0.142
R6973 GND.n222 GND.n218 0.142
R6974 GND.n165 GND.n161 0.141
R6975 GND.n116 GND.n112 0.136
R6976 GND.n173 GND.n169 0.136
R6977 GND.n104 GND.n103 0.125
R6978 GND.n372 GND.n371 0.125
R6979 GND GND.n381 0.114
R6980 GND.n202 GND.n201 0.045
R6981 GND.n147 GND.n146 0.044
R6982 GND.n203 GND.n202 0.044
R6983 GND.n146 GND.n145 0.044
R6984 GND.n110 GND.n104 0.017
R6985 GND.n380 GND.n372 0.017
R6986 GND.n303 GND.n302 0.016
R6987 GND.n302 GND.t0 0.016
R6988 GND.n301 GND.n300 0.016
R6989 GND.t0 GND.n301 0.016
R6990 GND.n111 GND.n110 0.012
R6991 GND.n381 GND.n380 0.012
R6992 GND.n145 GND.n142 0.001
R6993 GND.n201 GND.n198 0.001
C6 VBIAS GND 2.56fF
C7 IND_CT GND 0.27fF
C8 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE GND 4.18fF
C9 VDD GND 30.68fF
C10 VBIAS.n0 GND 0.02fF
C11 VBIAS.n1 GND 0.05fF
C12 VBIAS.n2 GND 0.01fF
C13 VBIAS.n4 GND 0.04fF
C14 VBIAS.n6 GND 0.03fF
C15 VBIAS.n8 GND 0.04fF
C16 VBIAS.n10 GND 0.04fF
C17 VBIAS.n12 GND 0.01fF
C18 VBIAS.n14 GND 0.02fF
C19 VBIAS.n16 GND 0.03fF
C20 VBIAS.n18 GND 0.08fF
C21 VBIAS.n20 GND 0.01fF
C22 VBIAS.n22 GND 0.01fF
C23 VBIAS.n24 GND 0.01fF
C24 VBIAS.n25 GND 0.04fF
C25 VBIAS.n26 GND 0.02fF
C26 VBIAS.n27 GND 0.01fF
C27 VBIAS.n28 GND 0.01fF
C28 VBIAS.n30 GND 0.02fF
C29 VBIAS.n32 GND 0.03fF
C30 VBIAS.n34 GND 0.02fF
C31 VBIAS.n36 GND 0.01fF
C32 VBIAS.n38 GND 0.04fF
C33 VBIAS.n40 GND 0.04fF
C34 VBIAS.n43 GND 0.01fF
C35 VBIAS.n44 GND 0.05fF
C36 VBIAS.n45 GND 0.02fF
C37 VBIAS.n46 GND 0.01fF
C38 VBIAS.n48 GND 0.01fF
C39 VBIAS.n50 GND 0.01fF
C40 VBIAS.n52 GND 0.01fF
C41 VBIAS.n53 GND 0.09fF
C42 VBIAS.n54 GND 0.01fF
C43 VBIAS.n55 GND 0.05fF
C44 VBIAS.n56 GND 0.01fF
C45 VBIAS.n58 GND 0.01fF
C46 VBIAS.n60 GND 0.03fF
C47 VBIAS.n61 GND 0.03fF
C48 VBIAS.t0 GND 0.11fF $ **FLOATING
C49 VBIAS.n63 GND 0.01fF
C50 VBIAS.n65 GND 0.01fF
C51 VBIAS.n67 GND 0.01fF
C52 VBIAS.n69 GND 0.01fF
C53 VBIAS.n70 GND 0.03fF
C54 VBIAS.n71 GND 0.04fF
C55 VBIAS.n72 GND 0.01fF
C56 VBIAS.n74 GND 0.01fF
C57 VBIAS.n76 GND 0.01fF
C58 VBIAS.n77 GND 0.05fF
C59 VBIAS.n78 GND 0.91fF
C60 VBIAS.n80 GND 0.11fF
C61 IND_CT.n0 GND 0.00fF
C62 IND_CT.n1 GND 0.01fF
C63 IND_CT.n2 GND 0.01fF
C64 IND_CT.n3 GND 0.01fF
C65 IND_CT.n4 GND 0.00fF
C66 IND_CT.n5 GND 0.00fF
C67 IND_CT.n6 GND 0.00fF
C68 IND_CT.n7 GND 0.00fF
C69 IND_CT.n8 GND 0.00fF
C70 IND_CT.n9 GND 0.01fF
C71 IND_CT.n10 GND 0.01fF
C72 IND_CT.n11 GND 0.01fF
C73 IND_CT.n12 GND 0.01fF
C74 IND_CT.n13 GND 0.01fF
C75 IND_CT.n14 GND 0.01fF
C76 IND_CT.n15 GND 0.01fF
C77 IND_CT.n16 GND 0.00fF
C78 IND_CT.n17 GND 0.01fF
C79 IND_CT.t10 GND 0.11fF $ **FLOATING
C80 IND_CT.t13 GND 0.11fF $ **FLOATING
C81 IND_CT.n18 GND 0.28fF
C82 IND_CT.n19 GND 0.11fF
C83 IND_CT.n20 GND 0.19fF
C84 IND_CT.n21 GND 0.12fF
C85 IND_CT.n22 GND 0.01fF
C86 IND_CT.n23 GND 0.04fF
C87 IND_CT.n24 GND 0.01fF
C88 IND_CT.n25 GND 0.05fF
C89 IND_CT.n26 GND 0.02fF
C90 IND_CT.n27 GND 0.04fF
C91 IND_CT.n28 GND 0.00fF
C92 IND_CT.n29 GND 0.02fF
C93 IND_CT.n30 GND 0.02fF
C94 IND_CT.n31 GND 0.00fF
C95 IND_CT.n32 GND 0.01fF
C96 IND_CT.n33 GND 0.01fF
C97 IND_CT.n34 GND 0.00fF
C98 IND_CT.n35 GND 0.01fF
C99 IND_CT.n36 GND 0.01fF
C100 IND_CT.n37 GND 0.01fF
C101 IND_CT.n38 GND 0.01fF
C102 IND_CT.n39 GND 0.00fF
C103 IND_CT.n40 GND 0.01fF
C104 IND_CT.n41 GND 0.01fF
C105 IND_CT.n42 GND 0.00fF
C106 IND_CT.n43 GND 0.01fF
C107 IND_CT.n44 GND 0.01fF
C108 IND_CT.n45 GND 0.00fF
C109 IND_CT.n46 GND 0.00fF
C110 IND_CT.n47 GND 0.01fF
C111 IND_CT.n48 GND 0.01fF
C112 IND_CT.n49 GND 0.06fF
C113 IND_CT.n50 GND 0.26fF
C114 IND_CT.n51 GND 0.25fF
C115 IND_CT.n52 GND 0.26fF
C116 IND_CT.n53 GND 0.00fF
C117 IND_CT.n54 GND 0.25fF
C118 IND_CT.n55 GND 0.86fF
C119 IND_CT.n56 GND 0.00fF
C120 IND_CT.n57 GND 0.25fF
C121 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/DRAIN GND 0.01fF
C122 IND_CT.n59 GND 0.04fF
C123 IND_CT.n60 GND 0.04fF
C124 IND_CT.n61 GND 0.02fF
C125 IND_CT.n63 GND 0.02fF
C126 IND_CT.n64 GND 0.03fF
C127 IND_CT.n65 GND 0.04fF
C128 IND_CT.n66 GND 0.03fF
C129 IND_CT.n67 GND 0.04fF
C130 IND_CT.n68 GND 0.04fF
C131 IND_CT.n69 GND 0.03fF
C132 IND_CT.n70 GND 0.02fF
C133 IND_CT.n71 GND 0.01fF
C134 IND_CT.n72 GND 0.02fF
C135 IND_CT.n73 GND 0.03fF
C136 IND_CT.n74 GND 0.03fF
C137 IND_CT.n75 GND 0.04fF
C138 IND_CT.n76 GND 0.03fF
C139 IND_CT.n77 GND 0.04fF
C140 IND_CT.n78 GND 0.01fF
C141 IND_CT.t6 GND 0.11fF $ **FLOATING
C142 IND_CT.t12 GND 0.11fF $ **FLOATING
C143 IND_CT.n79 GND 0.28fF
C144 IND_CT.n80 GND 0.12fF
C145 IND_CT.n81 GND 0.00fF
C146 IND_CT.n82 GND 0.01fF
C147 IND_CT.n83 GND 0.02fF
C148 IND_CT.n84 GND 0.02fF
C149 IND_CT.n85 GND 0.00fF
C150 IND_CT.n86 GND 0.01fF
C151 IND_CT.n87 GND 0.01fF
C152 IND_CT.n88 GND 0.01fF
C153 IND_CT.n89 GND 0.01fF
C154 IND_CT.n90 GND 0.00fF
C155 IND_CT.n91 GND 0.01fF
C156 IND_CT.n92 GND 0.01fF
C157 IND_CT.n93 GND 0.01fF
C158 IND_CT.n94 GND 0.01fF
C159 IND_CT.n95 GND 0.01fF
C160 IND_CT.n96 GND 0.00fF
C161 IND_CT.n97 GND 0.00fF
C162 IND_CT.n98 GND 0.01fF
C163 IND_CT.n99 GND 0.01fF
C164 IND_CT.n100 GND 0.01fF
C165 IND_CT.n101 GND 0.01fF
C166 IND_CT.n102 GND 0.01fF
C167 IND_CT.n103 GND 0.01fF
C168 IND_CT.n104 GND 0.00fF
C169 IND_CT.n105 GND 0.00fF
C170 IND_CT.n106 GND 0.00fF
C171 IND_CT.n107 GND 0.00fF
C172 IND_CT.n108 GND 0.00fF
C173 IND_CT.n109 GND 0.00fF
C174 IND_CT.n110 GND 0.01fF
C175 IND_CT.n111 GND 0.01fF
C176 IND_CT.n112 GND 0.01fF
C177 IND_CT.n113 GND 0.01fF
C178 IND_CT.n114 GND 0.01fF
C179 IND_CT.n115 GND 0.01fF
C180 IND_CT.n116 GND 0.00fF
C181 IND_CT.n117 GND 0.18fF
C182 IND_CT.n118 GND 0.14fF
C183 IND_CT.n119 GND 0.04fF
C184 IND_CT.n120 GND 0.01fF
C185 IND_CT.n121 GND 0.04fF
C186 IND_CT.n122 GND 0.03fF
C187 IND_CT.n123 GND 0.04fF
C188 IND_CT.n124 GND 0.01fF
C189 IND_CT.t15 GND 0.11fF $ **FLOATING
C190 IND_CT.t1 GND 0.11fF $ **FLOATING
C191 IND_CT.n125 GND 0.28fF
C192 IND_CT.n126 GND 0.12fF
C193 IND_CT.n127 GND 0.00fF
C194 IND_CT.n128 GND 0.01fF
C195 IND_CT.n129 GND 0.00fF
C196 IND_CT.n130 GND 0.02fF
C197 IND_CT.n131 GND 0.02fF
C198 IND_CT.n132 GND 0.01fF
C199 IND_CT.n133 GND 0.01fF
C200 IND_CT.n134 GND 0.01fF
C201 IND_CT.n135 GND 0.01fF
C202 IND_CT.n136 GND 0.00fF
C203 IND_CT.n137 GND 0.01fF
C204 IND_CT.n138 GND 0.01fF
C205 IND_CT.n139 GND 0.01fF
C206 IND_CT.n140 GND 0.00fF
C207 IND_CT.n141 GND 0.01fF
C208 IND_CT.n142 GND 0.01fF
C209 IND_CT.n143 GND 0.00fF
C210 IND_CT.n144 GND 0.00fF
C211 IND_CT.n145 GND 0.01fF
C212 IND_CT.n146 GND 0.01fF
C213 IND_CT.n147 GND 0.01fF
C214 IND_CT.n148 GND 0.01fF
C215 IND_CT.n149 GND 0.01fF
C216 IND_CT.n150 GND 0.01fF
C217 IND_CT.n151 GND 0.00fF
C218 IND_CT.n152 GND 0.00fF
C219 IND_CT.n153 GND 0.00fF
C220 IND_CT.n154 GND 0.00fF
C221 IND_CT.n155 GND 0.00fF
C222 IND_CT.n156 GND 0.01fF
C223 IND_CT.n157 GND 0.01fF
C224 IND_CT.n158 GND 0.01fF
C225 IND_CT.n159 GND 0.01fF
C226 IND_CT.n160 GND 0.01fF
C227 IND_CT.n161 GND 0.01fF
C228 IND_CT.n162 GND 0.00fF
C229 IND_CT.n163 GND 0.18fF
C230 IND_CT.n164 GND 0.14fF
C231 IND_CT.n165 GND 0.04fF
C232 IND_CT.n166 GND 0.01fF
C233 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/DRAIN GND 0.01fF
C234 IND_CT.n167 GND 0.04fF
C235 IND_CT.n168 GND 0.04fF
C236 IND_CT.n169 GND 0.02fF
C237 IND_CT.n171 GND 0.02fF
C238 IND_CT.n172 GND 0.03fF
C239 IND_CT.n173 GND 0.04fF
C240 IND_CT.n174 GND 0.03fF
C241 IND_CT.n175 GND 0.04fF
C242 IND_CT.n176 GND 0.04fF
C243 IND_CT.n177 GND 0.03fF
C244 IND_CT.n178 GND 0.02fF
C245 IND_CT.n179 GND 0.01fF
C246 IND_CT.n180 GND 0.02fF
C247 IND_CT.n181 GND 0.03fF
C248 IND_CT.n182 GND 0.03fF
C249 IND_CT.n183 GND 0.04fF
C250 IND_CT.n184 GND 0.03fF
C251 IND_CT.n185 GND 0.04fF
C252 IND_CT.n186 GND 0.01fF
C253 IND_CT.t5 GND 0.11fF $ **FLOATING
C254 IND_CT.t14 GND 0.11fF $ **FLOATING
C255 IND_CT.n187 GND 0.28fF
C256 IND_CT.n188 GND 0.12fF
C257 IND_CT.n189 GND 0.00fF
C258 IND_CT.n190 GND 0.01fF
C259 IND_CT.n191 GND 0.02fF
C260 IND_CT.n192 GND 0.02fF
C261 IND_CT.n193 GND 0.00fF
C262 IND_CT.n194 GND 0.01fF
C263 IND_CT.n195 GND 0.01fF
C264 IND_CT.n196 GND 0.01fF
C265 IND_CT.n197 GND 0.01fF
C266 IND_CT.n198 GND 0.00fF
C267 IND_CT.n199 GND 0.01fF
C268 IND_CT.n200 GND 0.01fF
C269 IND_CT.n201 GND 0.01fF
C270 IND_CT.n202 GND 0.01fF
C271 IND_CT.n203 GND 0.01fF
C272 IND_CT.n204 GND 0.00fF
C273 IND_CT.n205 GND 0.00fF
C274 IND_CT.n206 GND 0.01fF
C275 IND_CT.n207 GND 0.01fF
C276 IND_CT.n208 GND 0.01fF
C277 IND_CT.n209 GND 0.01fF
C278 IND_CT.n210 GND 0.01fF
C279 IND_CT.n211 GND 0.01fF
C280 IND_CT.n212 GND 0.00fF
C281 IND_CT.n213 GND 0.00fF
C282 IND_CT.n214 GND 0.00fF
C283 IND_CT.n215 GND 0.00fF
C284 IND_CT.n216 GND 0.00fF
C285 IND_CT.n217 GND 0.00fF
C286 IND_CT.n218 GND 0.01fF
C287 IND_CT.n219 GND 0.01fF
C288 IND_CT.n220 GND 0.01fF
C289 IND_CT.n221 GND 0.01fF
C290 IND_CT.n222 GND 0.01fF
C291 IND_CT.n223 GND 0.01fF
C292 IND_CT.n224 GND 0.00fF
C293 IND_CT.n225 GND 0.18fF
C294 IND_CT.n226 GND 0.14fF
C295 IND_CT.n227 GND 0.04fF
C296 IND_CT.n228 GND 0.01fF
C297 IND_CT.n229 GND 0.04fF
C298 IND_CT.n230 GND 0.03fF
C299 IND_CT.n231 GND 0.04fF
C300 IND_CT.n232 GND 0.01fF
C301 IND_CT.t3 GND 0.11fF $ **FLOATING
C302 IND_CT.t8 GND 0.11fF $ **FLOATING
C303 IND_CT.n233 GND 0.28fF
C304 IND_CT.n234 GND 0.12fF
C305 IND_CT.n235 GND 0.00fF
C306 IND_CT.n236 GND 0.01fF
C307 IND_CT.n237 GND 0.00fF
C308 IND_CT.n238 GND 0.02fF
C309 IND_CT.n239 GND 0.02fF
C310 IND_CT.n240 GND 0.01fF
C311 IND_CT.n241 GND 0.01fF
C312 IND_CT.n242 GND 0.01fF
C313 IND_CT.n243 GND 0.01fF
C314 IND_CT.n244 GND 0.00fF
C315 IND_CT.n245 GND 0.01fF
C316 IND_CT.n246 GND 0.01fF
C317 IND_CT.n247 GND 0.01fF
C318 IND_CT.n248 GND 0.00fF
C319 IND_CT.n249 GND 0.01fF
C320 IND_CT.n250 GND 0.01fF
C321 IND_CT.n251 GND 0.00fF
C322 IND_CT.n252 GND 0.00fF
C323 IND_CT.n253 GND 0.01fF
C324 IND_CT.n254 GND 0.01fF
C325 IND_CT.n255 GND 0.01fF
C326 IND_CT.n256 GND 0.01fF
C327 IND_CT.n257 GND 0.01fF
C328 IND_CT.n258 GND 0.01fF
C329 IND_CT.n259 GND 0.00fF
C330 IND_CT.n260 GND 0.00fF
C331 IND_CT.n261 GND 0.00fF
C332 IND_CT.n262 GND 0.00fF
C333 IND_CT.n263 GND 0.00fF
C334 IND_CT.n264 GND 0.01fF
C335 IND_CT.n265 GND 0.01fF
C336 IND_CT.n266 GND 0.01fF
C337 IND_CT.n267 GND 0.01fF
C338 IND_CT.n268 GND 0.01fF
C339 IND_CT.n269 GND 0.01fF
C340 IND_CT.n270 GND 0.00fF
C341 IND_CT.n271 GND 0.18fF
C342 IND_CT.n272 GND 0.14fF
C343 IND_CT.n273 GND 0.04fF
C344 IND_CT.n274 GND 0.01fF
C345 IND_CT.n275 GND 0.19fF
C346 IND_CT.n276 GND 0.13fF
C347 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/DRAIN GND 0.01fF
C348 IND_CT.n278 GND 0.04fF
C349 IND_CT.n279 GND 0.04fF
C350 IND_CT.n280 GND 0.02fF
C351 IND_CT.n282 GND 0.02fF
C352 IND_CT.n283 GND 0.03fF
C353 IND_CT.n284 GND 0.04fF
C354 IND_CT.n285 GND 0.03fF
C355 IND_CT.n286 GND 0.04fF
C356 IND_CT.n287 GND 0.04fF
C357 IND_CT.n288 GND 0.03fF
C358 IND_CT.n289 GND 0.02fF
C359 IND_CT.n290 GND 0.03fF
C360 IND_CT.n291 GND 0.03fF
C361 IND_CT.n292 GND 0.03fF
C362 IND_CT.n293 GND 0.01fF
C363 IND_CT.n294 GND 0.09fF
C364 IND_CT.n296 GND 0.13fF
C365 IND_CT.n297 GND 0.45fF
C366 IND_CT.n298 GND 0.45fF
C367 IND_CT.n299 GND 0.13fF
C368 IND_CT.n301 GND 0.09fF
C369 IND_CT.n303 GND 0.13fF
C370 IND_CT.n304 GND 1.08fF
C371 IND_CT.n305 GND 1.08fF
C372 IND_CT.n306 GND 0.13fF
C373 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/DRAIN GND 0.01fF
C374 IND_CT.n308 GND 0.04fF
C375 IND_CT.n309 GND 0.04fF
C376 IND_CT.n310 GND 0.02fF
C377 IND_CT.n312 GND 0.02fF
C378 IND_CT.n313 GND 0.03fF
C379 IND_CT.n314 GND 0.04fF
C380 IND_CT.n315 GND 0.03fF
C381 IND_CT.n316 GND 0.04fF
C382 IND_CT.n317 GND 0.04fF
C383 IND_CT.n318 GND 0.03fF
C384 IND_CT.n319 GND 0.02fF
C385 IND_CT.n320 GND 0.03fF
C386 IND_CT.n321 GND 0.03fF
C387 IND_CT.n322 GND 0.03fF
C388 IND_CT.n323 GND 0.01fF
C389 IND_CT.n324 GND 0.09fF
C390 IND_CT.n326 GND 0.13fF
C391 IND_CT.n327 GND 0.45fF
C392 IND_CT.n328 GND 0.45fF
C393 IND_CT.n329 GND 0.13fF
C394 IND_CT.n331 GND 0.09fF
C395 IND_CT.n333 GND 0.13fF
C396 IND_CT.n334 GND 0.44fF
C397 IND_CT.n335 GND 0.48fF
C398 IND_CT.n337 GND 0.25fF
C399 IND_CT.n338 GND 0.26fF
C400 IND_CT.n339 GND 1.36fF
C401 IND_CT.n340 GND 1.36fF
C402 IND_CT.n342 GND 0.48fF
C403 IND_CT.n343 GND 0.44fF
C404 IND_CT.n344 GND 0.13fF
C405 IND_CT.n346 GND 0.00fF
C406 IND_CT.n347 GND 0.00fF
C407 IND_CT.n348 GND 0.02fF
C408 IND_CT.n349 GND 0.02fF
C409 IND_CT.n350 GND 0.01fF
C410 IND_CT.n351 GND 0.01fF
C411 IND_CT.n352 GND 0.00fF
C412 IND_CT.n353 GND 0.01fF
C413 IND_CT.n354 GND 0.01fF
C414 IND_CT.n355 GND 0.01fF
C415 IND_CT.n356 GND 0.01fF
C416 IND_CT.n357 GND 0.00fF
C417 IND_CT.n358 GND 0.01fF
C418 IND_CT.n359 GND 0.01fF
C419 IND_CT.n360 GND 0.00fF
C420 IND_CT.n361 GND 0.01fF
C421 IND_CT.n362 GND 0.01fF
C422 IND_CT.n363 GND 0.00fF
C423 IND_CT.n364 GND 0.00fF
C424 IND_CT.n365 GND 0.01fF
C425 IND_CT.n366 GND 0.01fF
C426 IND_CT.n367 GND 0.06fF
C427 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/DRAIN GND 0.02fF
C428 IND_CT.n368 GND 0.04fF
C429 IND_CT.n369 GND 0.04fF
C430 IND_CT.n370 GND 0.03fF
C431 IND_CT.n372 GND 0.02fF
C432 IND_CT.n373 GND 0.03fF
C433 IND_CT.n374 GND 0.02fF
C434 IND_CT.n375 GND 0.02fF
C435 IND_CT.n376 GND 0.02fF
C436 IND_CT.n377 GND 0.04fF
C437 IND_CT.n378 GND 0.03fF
C438 IND_CT.n379 GND 0.03fF
C439 IND_CT.n380 GND 0.03fF
C440 IND_CT.n381 GND 0.04fF
C441 IND_CT.n383 GND 0.04fF
C442 IND_CT.n384 GND 0.02fF
C443 IND_CT.n385 GND 0.05fF
C444 IND_CT.n386 GND 0.01fF
C445 IND_CT.t9 GND 0.11fF $ **FLOATING
C446 IND_CT.t11 GND 0.11fF $ **FLOATING
C447 IND_CT.n387 GND 0.28fF
C448 IND_CT.n388 GND 0.12fF
C449 IND_CT.n389 GND 0.01fF
C450 IND_CT.n390 GND 0.01fF
C451 IND_CT.n391 GND 0.01fF
C452 IND_CT.n392 GND 0.00fF
C453 IND_CT.n393 GND 0.00fF
C454 IND_CT.n394 GND 0.00fF
C455 IND_CT.n395 GND 0.00fF
C456 IND_CT.n396 GND 0.00fF
C457 IND_CT.n397 GND 0.00fF
C458 IND_CT.n398 GND 0.01fF
C459 IND_CT.n399 GND 0.01fF
C460 IND_CT.n400 GND 0.01fF
C461 IND_CT.n401 GND 0.01fF
C462 IND_CT.n402 GND 0.01fF
C463 IND_CT.n403 GND 0.01fF
C464 IND_CT.n404 GND 0.01fF
C465 IND_CT.n405 GND 0.00fF
C466 IND_CT.n406 GND 0.19fF
C467 IND_CT.n407 GND 0.12fF
C468 IND_CT.n408 GND 0.01fF
C469 IND_CT.n409 GND 0.04fF
C470 IND_CT.n410 GND 0.01fF
C471 IND_CT.n411 GND 0.09fF
C472 IND_CT.n413 GND 0.13fF
C473 IND_CT.n414 GND 0.45fF
C474 IND_CT.n415 GND 0.45fF
C475 IND_CT.n416 GND 0.13fF
C476 IND_CT.n418 GND 0.04fF
C477 IND_CT.n419 GND 0.02fF
C478 IND_CT.n420 GND 0.05fF
C479 IND_CT.n421 GND 0.01fF
C480 IND_CT.t7 GND 0.11fF $ **FLOATING
C481 IND_CT.t2 GND 0.11fF $ **FLOATING
C482 IND_CT.n422 GND 0.28fF
C483 IND_CT.n423 GND 0.12fF
C484 IND_CT.n424 GND 0.00fF
C485 IND_CT.n425 GND 0.01fF
C486 IND_CT.n426 GND 0.01fF
C487 IND_CT.n427 GND 0.01fF
C488 IND_CT.n428 GND 0.00fF
C489 IND_CT.n429 GND 0.00fF
C490 IND_CT.n430 GND 0.00fF
C491 IND_CT.n431 GND 0.00fF
C492 IND_CT.n432 GND 0.00fF
C493 IND_CT.n433 GND 0.01fF
C494 IND_CT.n434 GND 0.01fF
C495 IND_CT.n435 GND 0.01fF
C496 IND_CT.n436 GND 0.01fF
C497 IND_CT.n437 GND 0.01fF
C498 IND_CT.n438 GND 0.01fF
C499 IND_CT.n439 GND 0.01fF
C500 IND_CT.n440 GND 0.00fF
C501 IND_CT.n441 GND 0.19fF
C502 IND_CT.n442 GND 0.12fF
C503 IND_CT.n443 GND 0.01fF
C504 IND_CT.n444 GND 0.04fF
C505 IND_CT.n445 GND 0.01fF
C506 IND_CT.n446 GND 0.00fF
C507 IND_CT.n447 GND 0.00fF
C508 IND_CT.n448 GND 0.02fF
C509 IND_CT.n449 GND 0.02fF
C510 IND_CT.n450 GND 0.01fF
C511 IND_CT.n451 GND 0.01fF
C512 IND_CT.n452 GND 0.00fF
C513 IND_CT.n453 GND 0.01fF
C514 IND_CT.n454 GND 0.01fF
C515 IND_CT.n455 GND 0.01fF
C516 IND_CT.n456 GND 0.01fF
C517 IND_CT.n457 GND 0.00fF
C518 IND_CT.n458 GND 0.01fF
C519 IND_CT.n459 GND 0.01fF
C520 IND_CT.n460 GND 0.00fF
C521 IND_CT.n461 GND 0.01fF
C522 IND_CT.n462 GND 0.01fF
C523 IND_CT.n463 GND 0.00fF
C524 IND_CT.n464 GND 0.00fF
C525 IND_CT.n465 GND 0.01fF
C526 IND_CT.n466 GND 0.01fF
C527 IND_CT.n467 GND 0.06fF
C528 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/DRAIN GND 0.02fF
C529 IND_CT.n468 GND 0.04fF
C530 IND_CT.n469 GND 0.04fF
C531 IND_CT.n470 GND 0.03fF
C532 IND_CT.n472 GND 0.02fF
C533 IND_CT.n473 GND 0.02fF
C534 IND_CT.n474 GND 0.03fF
C535 IND_CT.n475 GND 0.02fF
C536 IND_CT.n476 GND 0.02fF
C537 IND_CT.n477 GND 0.04fF
C538 IND_CT.n478 GND 0.03fF
C539 IND_CT.n479 GND 0.03fF
C540 IND_CT.n480 GND 0.03fF
C541 IND_CT.n481 GND 0.04fF
C542 IND_CT.n483 GND 0.09fF
C543 IND_CT.n485 GND 0.13fF
C544 IND_CT.n486 GND 1.08fF
C545 IND_CT.n487 GND 1.08fF
C546 IND_CT.n488 GND 0.13fF
C547 IND_CT.n490 GND 0.00fF
C548 IND_CT.n491 GND 0.00fF
C549 IND_CT.n492 GND 0.02fF
C550 IND_CT.n493 GND 0.02fF
C551 IND_CT.n494 GND 0.01fF
C552 IND_CT.n495 GND 0.01fF
C553 IND_CT.n496 GND 0.00fF
C554 IND_CT.n497 GND 0.01fF
C555 IND_CT.n498 GND 0.01fF
C556 IND_CT.n499 GND 0.01fF
C557 IND_CT.n500 GND 0.01fF
C558 IND_CT.n501 GND 0.00fF
C559 IND_CT.n502 GND 0.01fF
C560 IND_CT.n503 GND 0.01fF
C561 IND_CT.n504 GND 0.00fF
C562 IND_CT.n505 GND 0.01fF
C563 IND_CT.n506 GND 0.01fF
C564 IND_CT.n507 GND 0.00fF
C565 IND_CT.n508 GND 0.00fF
C566 IND_CT.n509 GND 0.01fF
C567 IND_CT.n510 GND 0.01fF
C568 IND_CT.n511 GND 0.06fF
C569 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/DRAIN GND 0.02fF
C570 IND_CT.n512 GND 0.04fF
C571 IND_CT.n513 GND 0.04fF
C572 IND_CT.n514 GND 0.03fF
C573 IND_CT.n516 GND 0.02fF
C574 IND_CT.n517 GND 0.03fF
C575 IND_CT.n518 GND 0.02fF
C576 IND_CT.n519 GND 0.02fF
C577 IND_CT.n520 GND 0.02fF
C578 IND_CT.n521 GND 0.04fF
C579 IND_CT.n522 GND 0.03fF
C580 IND_CT.n523 GND 0.03fF
C581 IND_CT.n524 GND 0.03fF
C582 IND_CT.n525 GND 0.04fF
C583 IND_CT.n527 GND 0.04fF
C584 IND_CT.n528 GND 0.02fF
C585 IND_CT.n529 GND 0.05fF
C586 IND_CT.n530 GND 0.01fF
C587 IND_CT.t4 GND 0.11fF $ **FLOATING
C588 IND_CT.t0 GND 0.11fF $ **FLOATING
C589 IND_CT.n531 GND 0.28fF
C590 IND_CT.n532 GND 0.12fF
C591 IND_CT.n533 GND 0.01fF
C592 IND_CT.n534 GND 0.01fF
C593 IND_CT.n535 GND 0.01fF
C594 IND_CT.n536 GND 0.00fF
C595 IND_CT.n537 GND 0.00fF
C596 IND_CT.n538 GND 0.00fF
C597 IND_CT.n539 GND 0.00fF
C598 IND_CT.n540 GND 0.00fF
C599 IND_CT.n541 GND 0.00fF
C600 IND_CT.n542 GND 0.01fF
C601 IND_CT.n543 GND 0.01fF
C602 IND_CT.n544 GND 0.01fF
C603 IND_CT.n545 GND 0.01fF
C604 IND_CT.n546 GND 0.01fF
C605 IND_CT.n547 GND 0.01fF
C606 IND_CT.n548 GND 0.01fF
C607 IND_CT.n549 GND 0.00fF
C608 IND_CT.n550 GND 0.19fF
C609 IND_CT.n551 GND 0.12fF
C610 IND_CT.n552 GND 0.01fF
C611 IND_CT.n553 GND 0.04fF
C612 IND_CT.n554 GND 0.01fF
C613 IND_CT.n555 GND 0.09fF
C614 IND_CT.n557 GND 0.13fF
C615 IND_CT.n558 GND 0.45fF
C616 IND_CT.n559 GND 0.45fF
C617 IND_CT.n560 GND 0.13fF
C618 IND_CT.n562 GND 0.19fF
C619 IND_CT.n563 GND 0.13fF
C620 IND_CT.n565 GND 0.09fF
C621 IND_CT.n567 GND 0.04fF
C622 IND_CT.n568 GND 0.03fF
C623 IND_CT.n569 GND 0.03fF
C624 IND_CT.n570 GND 0.03fF
C625 IND_CT.n571 GND 0.04fF
C626 IND_CT.n572 GND 0.02fF
C627 IND_CT.n573 GND 0.02fF
C628 IND_CT.n574 GND 0.02fF
C629 IND_CT.n575 GND 0.03fF
C630 IND_CT.n576 GND 0.02fF
C631 IND_CT.n578 GND 0.03fF
C632 IND_CT.n579 GND 0.04fF
C633 IND_CT.n580 GND 0.04fF
C634 VDD.n0 GND 0.01fF
C635 VDD.n1 GND 0.01fF
C636 VDD.n2 GND 0.00fF
C637 VDD.n3 GND 0.00fF
C638 VDD.n4 GND 0.00fF
C639 VDD.n5 GND 0.00fF
C640 VDD.n6 GND 0.00fF
C641 VDD.n7 GND 0.00fF
C642 VDD.n8 GND 0.00fF
C643 VDD.n9 GND 0.00fF
C644 VDD.n10 GND 0.00fF
C645 VDD.n11 GND 0.00fF
C646 VDD.n12 GND 0.00fF
C647 VDD.n13 GND 0.00fF
C648 VDD.n14 GND 0.00fF
C649 VDD.n15 GND 0.00fF
C650 VDD.n16 GND 0.00fF
C651 VDD.n17 GND 0.00fF
C652 VDD.n18 GND 0.00fF
C653 VDD.n19 GND 0.00fF
C654 VDD.n20 GND 0.00fF
C655 VDD.t60 GND 0.04fF $ **FLOATING
C656 VDD.n21 GND 0.13fF
C657 VDD.n22 GND 0.00fF
C658 VDD.n23 GND 0.04fF
C659 VDD.n24 GND 0.07fF
C660 VDD.n25 GND 0.00fF
C661 VDD.n26 GND 0.00fF
C662 VDD.n27 GND 0.00fF
C663 VDD.n28 GND 0.00fF
C664 VDD.n29 GND 0.00fF
C665 VDD.n30 GND 0.00fF
C666 VDD.n31 GND 0.00fF
C667 VDD.n32 GND 0.00fF
C668 VDD.n33 GND 0.00fF
C669 VDD.n34 GND 0.00fF
C670 VDD.n35 GND 0.00fF
C671 VDD.n36 GND 0.00fF
C672 VDD.n37 GND 0.00fF
C673 VDD.n38 GND 0.00fF
C674 VDD.n39 GND 0.00fF
C675 VDD.n40 GND 0.00fF
C676 VDD.n41 GND 0.00fF
C677 VDD.n42 GND 0.02fF
C678 VDD.n43 GND 0.01fF
C679 VDD.n44 GND 0.01fF
C680 VDD.n46 GND 0.01fF
C681 VDD.n47 GND 0.01fF
C682 VDD.n48 GND 0.01fF
C683 VDD.n50 GND 0.01fF
C684 VDD.n51 GND 0.01fF
C685 VDD.n52 GND 0.01fF
C686 VDD.n53 GND 0.01fF
C687 VDD.n54 GND 0.01fF
C688 VDD.n55 GND 0.01fF
C689 VDD.n56 GND 0.01fF
C690 VDD.n57 GND 0.09fF
C691 VDD.n58 GND 0.09fF
C692 VDD.n59 GND 0.01fF
C693 VDD.n60 GND 0.03fF
C694 VDD.n61 GND 0.01fF
C695 VDD.n62 GND 0.01fF
C696 VDD.n63 GND 0.01fF
C697 VDD.n64 GND 0.00fF
C698 VDD.n65 GND 0.00fF
C699 VDD.n66 GND 0.01fF
C700 VDD.n67 GND 0.01fF
C701 VDD.n68 GND 0.01fF
C702 VDD.n69 GND 0.01fF
C703 VDD.n70 GND 0.03fF
C704 VDD.n71 GND 0.01fF
C705 VDD.n72 GND 0.00fF
C706 VDD.n73 GND 0.01fF
C707 VDD.n74 GND 0.01fF
C708 VDD.n75 GND 0.04fF
C709 VDD.n76 GND 0.05fF
C710 VDD.n77 GND 0.04fF
C711 VDD.n78 GND 0.04fF
C712 VDD.n80 GND 0.05fF
C713 VDD.n81 GND 0.03fF
C714 VDD.n82 GND 0.02fF
C715 VDD.n83 GND 0.03fF
C716 VDD.n84 GND 0.00fF
C717 VDD.n85 GND 0.01fF
C718 VDD.n86 GND 0.01fF
C719 VDD.n87 GND 0.01fF
C720 VDD.n88 GND 0.03fF
C721 VDD.n89 GND 0.01fF
C722 VDD.n90 GND 0.00fF
C723 VDD.n91 GND 0.01fF
C724 VDD.n92 GND 0.01fF
C725 VDD.n93 GND 0.05fF
C726 VDD.n94 GND 0.03fF
C727 VDD.n95 GND 0.02fF
C728 VDD.n96 GND 0.03fF
C729 VDD.n97 GND 0.05fF
C730 VDD.n98 GND 0.02fF
C731 VDD.n99 GND 0.03fF
C732 VDD.n100 GND 0.02fF
C733 VDD.n101 GND 0.03fF
C734 VDD.n102 GND 0.00fF
C735 VDD.n103 GND 0.01fF
C736 VDD.n104 GND 0.00fF
C737 VDD.n105 GND 0.01fF
C738 VDD.n106 GND 0.01fF
C739 VDD.n107 GND 0.01fF
C740 VDD.n108 GND 0.04fF
C741 VDD.n109 GND 0.01fF
C742 VDD.n110 GND 0.01fF
C743 VDD.n111 GND 0.05fF
C744 VDD.n112 GND 0.03fF
C745 VDD.n113 GND 0.00fF
C746 VDD.n114 GND 0.01fF
C747 VDD.n115 GND 0.00fF
C748 VDD.n116 GND 0.01fF
C749 VDD.n117 GND 0.01fF
C750 VDD.n118 GND 0.01fF
C751 VDD.n119 GND 0.04fF
C752 VDD.n120 GND 0.01fF
C753 VDD.n121 GND 0.01fF
C754 VDD.n122 GND 0.02fF
C755 VDD.n123 GND 0.03fF
C756 VDD.n124 GND 0.05fF
C757 VDD.n126 GND 0.03fF
C758 VDD.n127 GND 0.00fF
C759 VDD.n128 GND 0.01fF
C760 VDD.n129 GND 0.01fF
C761 VDD.n130 GND 0.01fF
C762 VDD.n131 GND 0.01fF
C763 VDD.n132 GND 0.03fF
C764 VDD.n133 GND 0.01fF
C765 VDD.n134 GND 0.03fF
C766 VDD.n135 GND 0.01fF
C767 VDD.n136 GND 0.01fF
C768 VDD.n137 GND 0.01fF
C769 VDD.n138 GND 0.00fF
C770 VDD.n139 GND 0.00fF
C771 VDD.n140 GND 0.01fF
C772 VDD.n141 GND 0.01fF
C773 VDD.n142 GND 0.05fF
C774 VDD.n143 GND 0.04fF
C775 VDD.n144 GND 0.04fF
C776 VDD.n145 GND 0.05fF
C777 VDD.n146 GND 0.07fF
C778 VDD.n147 GND 0.02fF
C779 VDD.n148 GND 0.03fF
C780 VDD.n149 GND 0.00fF
C781 VDD.n150 GND 0.01fF
C782 VDD.n151 GND 0.01fF
C783 VDD.n152 GND 0.05fF
C784 VDD.n153 GND 0.02fF
C785 VDD.n154 GND 0.01fF
C786 VDD.n155 GND 0.05fF
C787 VDD.n156 GND 0.02fF
C788 VDD.n157 GND 0.03fF
C789 VDD.n158 GND 0.00fF
C790 VDD.n159 GND 0.01fF
C791 VDD.n160 GND 0.01fF
C792 VDD.n161 GND 0.00fF
C793 VDD.n162 GND 0.00fF
C794 VDD.n163 GND 0.00fF
C795 VDD.n164 GND 0.01fF
C796 VDD.n165 GND 0.01fF
C797 VDD.n166 GND 0.03fF
C798 VDD.n167 GND 0.01fF
C799 VDD.n168 GND 0.01fF
C800 VDD.n169 GND 0.00fF
C801 VDD.n170 GND 0.00fF
C802 VDD.n171 GND 0.00fF
C803 VDD.n172 GND 0.00fF
C804 VDD.n173 GND 0.00fF
C805 VDD.n174 GND 0.00fF
C806 VDD.n175 GND 0.00fF
C807 VDD.n176 GND 0.00fF
C808 VDD.n177 GND 0.00fF
C809 VDD.n178 GND 0.00fF
C810 VDD.n179 GND 0.00fF
C811 VDD.n180 GND 0.00fF
C812 VDD.n181 GND 0.00fF
C813 VDD.n182 GND 0.00fF
C814 VDD.n183 GND 0.00fF
C815 VDD.n184 GND 0.00fF
C816 VDD.n185 GND 0.00fF
C817 VDD.n186 GND 0.00fF
C818 VDD.n187 GND 0.00fF
C819 VDD.n188 GND 0.00fF
C820 VDD.n189 GND 0.00fF
C821 VDD.n190 GND 0.00fF
C822 VDD.n191 GND 0.00fF
C823 VDD.n192 GND 0.00fF
C824 VDD.n193 GND 0.00fF
C825 VDD.n194 GND 0.00fF
C826 VDD.n195 GND 0.00fF
C827 VDD.n196 GND 0.00fF
C828 VDD.n197 GND 0.00fF
C829 VDD.n198 GND 0.00fF
C830 VDD.n199 GND 0.00fF
C831 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/DRAIN GND 0.00fF
C832 VDD.n200 GND 0.01fF
C833 VDD.n201 GND 0.01fF
C834 VDD.n202 GND 0.01fF
C835 VDD.n203 GND 0.02fF
C836 VDD.n204 GND 0.02fF
C837 VDD.n205 GND 0.01fF
C838 VDD.n206 GND 0.01fF
C839 VDD.n207 GND 0.02fF
C840 VDD.n208 GND 0.02fF
C841 VDD.n209 GND 0.01fF
C842 VDD.n210 GND 0.03fF
C843 VDD.n211 GND 0.03fF
C844 VDD.n212 GND 0.04fF
C845 VDD.n213 GND 0.00fF
C846 VDD.n214 GND 0.00fF
C847 VDD.n215 GND 0.00fF
C848 VDD.n216 GND 0.00fF
C849 VDD.n217 GND 0.00fF
C850 VDD.n218 GND 0.01fF
C851 VDD.n219 GND 0.00fF
C852 VDD.n220 GND 0.01fF
C853 VDD.n221 GND 0.00fF
C854 VDD.n222 GND 0.00fF
C855 VDD.n223 GND 0.00fF
C856 VDD.n224 GND 0.00fF
C857 VDD.n225 GND 0.01fF
C858 VDD.n226 GND 0.00fF
C859 VDD.n227 GND 0.01fF
C860 VDD.n228 GND 0.00fF
C861 VDD.n229 GND 0.00fF
C862 VDD.n230 GND 0.00fF
C863 VDD.n231 GND 0.00fF
C864 VDD.n232 GND 0.01fF
C865 VDD.n233 GND 0.00fF
C866 VDD.n234 GND 0.01fF
C867 VDD.n235 GND 0.00fF
C868 VDD.n236 GND 0.00fF
C869 VDD.n237 GND 0.00fF
C870 VDD.n238 GND 0.00fF
C871 VDD.n239 GND 0.01fF
C872 VDD.n240 GND 0.00fF
C873 VDD.n241 GND 0.01fF
C874 VDD.n242 GND 0.00fF
C875 VDD.n243 GND 0.00fF
C876 VDD.n244 GND 0.07fF
C877 VDD.t32 GND 0.04fF $ **FLOATING
C878 VDD.n245 GND 0.07fF
C879 VDD.n246 GND 0.01fF
C880 VDD.n247 GND 0.01fF
C881 VDD.n248 GND 0.01fF
C882 VDD.n249 GND 0.01fF
C883 VDD.n250 GND 0.03fF
C884 VDD.n251 GND 0.01fF
C885 VDD.n252 GND 0.01fF
C886 VDD.n253 GND 0.63fF
C887 VDD.n254 GND 0.02fF
C888 VDD.n255 GND 0.01fF
C889 VDD.n256 GND 0.02fF
C890 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/BULK GND 0.01fF
C891 VDD.n257 GND 0.01fF
C892 VDD.n258 GND 0.01fF
C893 VDD.n259 GND 0.00fF
C894 VDD.n261 GND 0.00fF
C895 VDD.n262 GND 0.00fF
C896 VDD.n263 GND 0.00fF
C897 VDD.n264 GND 0.00fF
C898 VDD.n265 GND 0.00fF
C899 VDD.n266 GND 0.01fF
C900 VDD.n267 GND 0.01fF
C901 VDD.n268 GND 0.00fF
C902 VDD.n270 GND 0.01fF
C903 VDD.n272 GND 0.00fF
C904 VDD.n273 GND 0.00fF
C905 VDD.n274 GND 0.00fF
C906 VDD.n275 GND 0.00fF
C907 VDD.n276 GND 0.00fF
C908 VDD.n277 GND 0.00fF
C909 VDD.n278 GND 0.01fF
C910 VDD.n280 GND 0.01fF
C911 VDD.n281 GND 0.02fF
C912 VDD.n282 GND 0.01fF
C913 VDD.n283 GND 0.02fF
C914 VDD.n284 GND 0.01fF
C915 VDD.n285 GND 0.02fF
C916 VDD.n287 GND 0.01fF
C917 VDD.n289 GND 0.00fF
C918 VDD.n290 GND 0.00fF
C919 VDD.n291 GND 0.00fF
C920 VDD.n292 GND 0.01fF
C921 VDD.n293 GND 0.00fF
C922 VDD.n294 GND 0.00fF
C923 VDD.n295 GND 0.02fF
C924 VDD.n296 GND 0.01fF
C925 VDD.n297 GND 0.03fF
C926 VDD.n299 GND 0.01fF
C927 VDD.n301 GND 0.00fF
C928 VDD.n302 GND 0.00fF
C929 VDD.n303 GND 0.00fF
C930 VDD.n304 GND 0.00fF
C931 VDD.n305 GND 0.00fF
C932 VDD.n306 GND 0.00fF
C933 VDD.n307 GND 0.01fF
C934 VDD.n308 GND 0.01fF
C935 VDD.n310 GND 0.00fF
C936 VDD.n311 GND 0.00fF
C937 VDD.n312 GND 0.00fF
C938 VDD.n313 GND 0.00fF
C939 VDD.n314 GND 0.00fF
C940 VDD.n315 GND 0.00fF
C941 VDD.n316 GND 0.01fF
C942 VDD.n317 GND 0.00fF
C943 VDD.n318 GND 0.00fF
C944 VDD.n319 GND 0.00fF
C945 VDD.n320 GND 0.00fF
C946 VDD.n321 GND 0.00fF
C947 VDD.n322 GND 0.01fF
C948 VDD.n323 GND 0.01fF
C949 VDD.n324 GND 0.00fF
C950 VDD.n326 GND 0.00fF
C951 VDD.n327 GND 0.00fF
C952 VDD.n328 GND 0.00fF
C953 VDD.n329 GND 0.00fF
C954 VDD.n330 GND 0.00fF
C955 VDD.n331 GND 0.01fF
C956 VDD.n332 GND 0.01fF
C957 VDD.n333 GND 0.00fF
C958 VDD.n335 GND 0.35fF
C959 VDD.n336 GND 0.02fF
C960 VDD.n337 GND 0.00fF
C961 VDD.n338 GND 0.00fF
C962 VDD.n339 GND 0.00fF
C963 VDD.n340 GND 0.00fF
C964 VDD.n341 GND 0.02fF
C965 VDD.n342 GND 0.01fF
C966 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/BULK GND 0.01fF
C967 VDD.n343 GND 0.01fF
C968 VDD.n345 GND 0.00fF
C969 VDD.n346 GND 0.01fF
C970 VDD.n347 GND 0.00fF
C971 VDD.n348 GND 0.00fF
C972 VDD.n349 GND 0.00fF
C973 VDD.n350 GND 0.00fF
C974 VDD.n351 GND 0.00fF
C975 VDD.n352 GND 0.01fF
C976 VDD.n353 GND 0.01fF
C977 VDD.n354 GND 0.00fF
C978 VDD.n356 GND 0.01fF
C979 VDD.n358 GND 0.00fF
C980 VDD.n359 GND 0.00fF
C981 VDD.n360 GND 0.00fF
C982 VDD.n361 GND 0.00fF
C983 VDD.n362 GND 0.00fF
C984 VDD.n363 GND 0.00fF
C985 VDD.n364 GND 0.01fF
C986 VDD.n366 GND 0.00fF
C987 VDD.n367 GND 0.00fF
C988 VDD.n368 GND 0.00fF
C989 VDD.n369 GND 0.00fF
C990 VDD.n370 GND 0.00fF
C991 VDD.n371 GND 0.01fF
C992 VDD.n372 GND 0.01fF
C993 VDD.n373 GND 0.00fF
C994 VDD.n376 GND 0.01fF
C995 VDD.n377 GND 0.00fF
C996 VDD.n378 GND 0.00fF
C997 VDD.n379 GND 0.00fF
C998 VDD.n380 GND 0.00fF
C999 VDD.n381 GND 0.00fF
C1000 VDD.n382 GND 0.00fF
C1001 VDD.n383 GND 0.01fF
C1002 VDD.n385 GND 0.01fF
C1003 VDD.n387 GND 0.00fF
C1004 VDD.n388 GND 0.00fF
C1005 VDD.n389 GND 0.00fF
C1006 VDD.n390 GND 0.00fF
C1007 VDD.n391 GND 0.00fF
C1008 VDD.n392 GND 0.00fF
C1009 VDD.n393 GND 0.01fF
C1010 VDD.n395 GND 0.01fF
C1011 VDD.n396 GND 0.00fF
C1012 VDD.n397 GND 0.00fF
C1013 VDD.n398 GND 0.00fF
C1014 VDD.n399 GND 0.00fF
C1015 VDD.n400 GND 0.00fF
C1016 VDD.n401 GND 0.00fF
C1017 VDD.n402 GND 0.01fF
C1018 VDD.n404 GND 0.01fF
C1019 VDD.n406 GND 0.00fF
C1020 VDD.n407 GND 0.00fF
C1021 VDD.n408 GND 0.00fF
C1022 VDD.n409 GND 0.01fF
C1023 VDD.n410 GND 0.00fF
C1024 VDD.n411 GND 0.00fF
C1025 VDD.n412 GND 0.02fF
C1026 VDD.n413 GND 0.01fF
C1027 VDD.n414 GND 0.03fF
C1028 VDD.n416 GND 0.01fF
C1029 VDD.n417 GND 0.02fF
C1030 VDD.n418 GND 0.01fF
C1031 VDD.n419 GND 0.02fF
C1032 VDD.n421 GND 0.01fF
C1033 VDD.n422 GND 0.02fF
C1034 VDD.n425 GND 0.35fF
C1035 VDD.n427 GND 0.02fF
C1036 VDD.n428 GND 0.01fF
C1037 VDD.n429 GND 0.00fF
C1038 VDD.n430 GND 0.00fF
C1039 VDD.n431 GND 0.00fF
C1040 VDD.n432 GND 0.00fF
C1041 VDD.n433 GND 0.01fF
C1042 VDD.n434 GND 0.00fF
C1043 VDD.n435 GND 0.00fF
C1044 VDD.n436 GND 0.01fF
C1045 VDD.n437 GND 0.01fF
C1046 VDD.n438 GND 0.00fF
C1047 VDD.n439 GND 0.01fF
C1048 VDD.n440 GND 0.01fF
C1049 VDD.n441 GND 0.00fF
C1050 VDD.n442 GND 0.01fF
C1051 VDD.n443 GND 0.01fF
C1052 VDD.n444 GND 0.00fF
C1053 VDD.n445 GND 0.01fF
C1054 VDD.n446 GND 0.01fF
C1055 VDD.n447 GND 0.00fF
C1056 VDD.n448 GND 0.01fF
C1057 VDD.n449 GND 0.01fF
C1058 VDD.n450 GND 0.00fF
C1059 VDD.n451 GND 0.01fF
C1060 VDD.n452 GND 0.01fF
C1061 VDD.n453 GND 0.00fF
C1062 VDD.n454 GND 0.01fF
C1063 VDD.n455 GND 0.01fF
C1064 VDD.n456 GND 0.00fF
C1065 VDD.n457 GND 0.01fF
C1066 VDD.t33 GND 0.04fF $ **FLOATING
C1067 VDD.n458 GND 0.11fF
C1068 VDD.n459 GND 0.01fF
C1069 VDD.n460 GND 0.00fF
C1070 VDD.n461 GND 0.02fF
C1071 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/SOURCE GND 0.01fF
C1072 VDD.n462 GND 0.02fF
C1073 VDD.n463 GND 0.01fF
C1074 VDD.n464 GND 0.03fF
C1075 VDD.n465 GND 0.03fF
C1076 VDD.n466 GND 0.01fF
C1077 VDD.n467 GND 0.02fF
C1078 VDD.n468 GND 0.02fF
C1079 VDD.n469 GND 0.01fF
C1080 VDD.n470 GND 0.01fF
C1081 VDD.n471 GND 0.02fF
C1082 VDD.n472 GND 0.02fF
C1083 VDD.n473 GND 0.01fF
C1084 VDD.n474 GND 0.01fF
C1085 VDD.n475 GND 0.00fF
C1086 VDD.n476 GND 0.00fF
C1087 VDD.n477 GND 0.00fF
C1088 VDD.n478 GND 0.00fF
C1089 VDD.n479 GND 0.00fF
C1090 VDD.n480 GND 0.00fF
C1091 VDD.n481 GND 0.00fF
C1092 VDD.n482 GND 0.00fF
C1093 VDD.n483 GND 0.00fF
C1094 VDD.n484 GND 0.00fF
C1095 VDD.n485 GND 0.00fF
C1096 VDD.n486 GND 0.00fF
C1097 VDD.n487 GND 0.00fF
C1098 VDD.n488 GND 0.00fF
C1099 VDD.n489 GND 0.00fF
C1100 VDD.n490 GND 0.00fF
C1101 VDD.n491 GND 0.00fF
C1102 VDD.n492 GND 0.00fF
C1103 VDD.n493 GND 0.00fF
C1104 VDD.n494 GND 0.00fF
C1105 VDD.n495 GND 0.00fF
C1106 VDD.n496 GND 0.00fF
C1107 VDD.n497 GND 0.00fF
C1108 VDD.n498 GND 0.00fF
C1109 VDD.n499 GND 0.00fF
C1110 VDD.n500 GND 0.00fF
C1111 VDD.n501 GND 0.00fF
C1112 VDD.n502 GND 0.00fF
C1113 VDD.n503 GND 0.00fF
C1114 VDD.n504 GND 0.00fF
C1115 VDD.n505 GND 0.00fF
C1116 VDD.n506 GND 0.00fF
C1117 VDD.n507 GND 0.00fF
C1118 VDD.n508 GND 0.00fF
C1119 VDD.n509 GND 0.00fF
C1120 VDD.n510 GND 0.00fF
C1121 VDD.n511 GND 0.00fF
C1122 VDD.n512 GND 0.00fF
C1123 VDD.n513 GND 0.01fF
C1124 VDD.n514 GND 0.00fF
C1125 VDD.n515 GND 0.01fF
C1126 VDD.n516 GND 0.00fF
C1127 VDD.n517 GND 0.00fF
C1128 VDD.n518 GND 0.00fF
C1129 VDD.n519 GND 0.00fF
C1130 VDD.n520 GND 0.01fF
C1131 VDD.n521 GND 0.00fF
C1132 VDD.n522 GND 0.01fF
C1133 VDD.n523 GND 0.00fF
C1134 VDD.n524 GND 0.00fF
C1135 VDD.n525 GND 0.00fF
C1136 VDD.n526 GND 0.00fF
C1137 VDD.n527 GND 0.01fF
C1138 VDD.n528 GND 0.00fF
C1139 VDD.n529 GND 0.01fF
C1140 VDD.n530 GND 0.00fF
C1141 VDD.n531 GND 0.00fF
C1142 VDD.n532 GND 0.00fF
C1143 VDD.n533 GND 0.00fF
C1144 VDD.n534 GND 0.01fF
C1145 VDD.n535 GND 0.00fF
C1146 VDD.n536 GND 0.01fF
C1147 VDD.n537 GND 0.00fF
C1148 VDD.n538 GND 0.00fF
C1149 VDD.n539 GND 0.01fF
C1150 VDD.n540 GND 0.01fF
C1151 VDD.n541 GND 0.04fF
C1152 VDD.n542 GND 0.01fF
C1153 VDD.n543 GND 0.01fF
C1154 VDD.n544 GND 0.01fF
C1155 VDD.n545 GND 0.00fF
C1156 VDD.n546 GND 0.00fF
C1157 VDD.n547 GND 0.01fF
C1158 VDD.n548 GND 0.00fF
C1159 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/GATE GND 0.04fF
C1160 VDD.n549 GND 0.04fF
C1161 VDD.n550 GND 0.02fF
C1162 VDD.n551 GND 0.02fF
C1163 VDD.n552 GND 0.02fF
C1164 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/BULK GND 0.01fF
C1165 VDD.n553 GND 0.01fF
C1166 VDD.n554 GND 0.00fF
C1167 VDD.n555 GND 0.00fF
C1168 VDD.n556 GND 0.00fF
C1169 VDD.n557 GND 0.00fF
C1170 VDD.n558 GND 0.00fF
C1171 VDD.n559 GND 0.01fF
C1172 VDD.n561 GND 0.00fF
C1173 VDD.n562 GND 0.01fF
C1174 VDD.n563 GND 0.00fF
C1175 VDD.n564 GND 0.01fF
C1176 VDD.n565 GND 0.00fF
C1177 VDD.n566 GND 0.01fF
C1178 VDD.n567 GND 0.00fF
C1179 VDD.n568 GND 0.00fF
C1180 VDD.n569 GND 0.00fF
C1181 VDD.n570 GND 0.00fF
C1182 VDD.n571 GND 0.01fF
C1183 VDD.n572 GND 0.00fF
C1184 VDD.n574 GND 0.01fF
C1185 VDD.n575 GND 0.00fF
C1186 VDD.n576 GND 0.01fF
C1187 VDD.n577 GND 0.00fF
C1188 VDD.n578 GND 0.01fF
C1189 VDD.n579 GND 0.00fF
C1190 VDD.n580 GND 0.00fF
C1191 VDD.n581 GND 0.00fF
C1192 VDD.n582 GND 0.00fF
C1193 VDD.n583 GND 0.01fF
C1194 VDD.n585 GND 0.00fF
C1195 VDD.n587 GND 0.01fF
C1196 VDD.n588 GND 0.00fF
C1197 VDD.n589 GND 0.01fF
C1198 VDD.n590 GND 0.00fF
C1199 VDD.n591 GND 0.01fF
C1200 VDD.n592 GND 0.00fF
C1201 VDD.n593 GND 0.00fF
C1202 VDD.n594 GND 0.00fF
C1203 VDD.n595 GND 0.00fF
C1204 VDD.n596 GND 0.01fF
C1205 VDD.n597 GND 0.00fF
C1206 VDD.n599 GND 0.01fF
C1207 VDD.n600 GND 0.00fF
C1208 VDD.n601 GND 0.01fF
C1209 VDD.n602 GND 0.00fF
C1210 VDD.n603 GND 0.00fF
C1211 VDD.n605 GND 0.01fF
C1212 VDD.n606 GND 0.00fF
C1213 VDD.n608 GND 0.01fF
C1214 VDD.n609 GND 0.00fF
C1215 VDD.n610 GND 0.01fF
C1216 VDD.n611 GND 0.00fF
C1217 VDD.n612 GND 0.00fF
C1218 VDD.n613 GND 0.00fF
C1219 VDD.n614 GND 0.01fF
C1220 VDD.n615 GND 0.00fF
C1221 VDD.n616 GND 0.00fF
C1222 VDD.n617 GND 0.01fF
C1223 VDD.n619 GND 0.00fF
C1224 VDD.n621 GND 0.01fF
C1225 VDD.n622 GND 0.00fF
C1226 VDD.n623 GND 0.01fF
C1227 VDD.n624 GND 0.00fF
C1228 VDD.n625 GND 0.00fF
C1229 VDD.n626 GND 0.00fF
C1230 VDD.n627 GND 0.01fF
C1231 VDD.n628 GND 0.00fF
C1232 VDD.n629 GND 0.00fF
C1233 VDD.n630 GND 0.01fF
C1234 VDD.n631 GND 0.00fF
C1235 VDD.n633 GND 0.01fF
C1236 VDD.n634 GND 0.00fF
C1237 VDD.n635 GND 0.01fF
C1238 VDD.n636 GND 0.00fF
C1239 VDD.n637 GND 0.00fF
C1240 VDD.n638 GND 0.00fF
C1241 VDD.n639 GND 0.01fF
C1242 VDD.n640 GND 0.00fF
C1243 VDD.n641 GND 0.00fF
C1244 VDD.n642 GND 0.01fF
C1245 VDD.n644 GND 0.00fF
C1246 VDD.n645 GND 0.01fF
C1247 VDD.n646 GND 0.00fF
C1248 VDD.n647 GND 0.01fF
C1249 VDD.n648 GND 0.00fF
C1250 VDD.n649 GND 0.00fF
C1251 VDD.n650 GND 0.01fF
C1252 VDD.n651 GND 0.01fF
C1253 VDD.n652 GND 0.02fF
C1254 VDD.n653 GND 0.01fF
C1255 VDD.n654 GND 0.02fF
C1256 VDD.n655 GND 0.02fF
C1257 VDD.n656 GND 0.01fF
C1258 VDD.n657 GND 0.02fF
C1259 VDD.n658 GND 0.01fF
C1260 VDD.n659 GND 0.02fF
C1261 VDD.n660 GND 0.01fF
C1262 VDD.n661 GND 0.01fF
C1263 VDD.n662 GND 0.01fF
C1264 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/BULK GND 0.01fF
C1265 VDD.n663 GND 0.01fF
C1266 VDD.n664 GND 0.01fF
C1267 VDD.n665 GND 0.00fF
C1268 VDD.n667 GND 0.00fF
C1269 VDD.n668 GND 0.00fF
C1270 VDD.n669 GND 0.00fF
C1271 VDD.n670 GND 0.00fF
C1272 VDD.n671 GND 0.00fF
C1273 VDD.n672 GND 0.01fF
C1274 VDD.n673 GND 0.01fF
C1275 VDD.n674 GND 0.00fF
C1276 VDD.n676 GND 0.01fF
C1277 VDD.n678 GND 0.00fF
C1278 VDD.n679 GND 0.00fF
C1279 VDD.n680 GND 0.00fF
C1280 VDD.n681 GND 0.00fF
C1281 VDD.n682 GND 0.00fF
C1282 VDD.n683 GND 0.00fF
C1283 VDD.n684 GND 0.01fF
C1284 VDD.n687 GND 0.01fF
C1285 VDD.n688 GND 0.02fF
C1286 VDD.n689 GND 0.01fF
C1287 VDD.n690 GND 0.02fF
C1288 VDD.n691 GND 0.01fF
C1289 VDD.n692 GND 0.02fF
C1290 VDD.n694 GND 0.01fF
C1291 VDD.n696 GND 0.00fF
C1292 VDD.n697 GND 0.00fF
C1293 VDD.n698 GND 0.00fF
C1294 VDD.n699 GND 0.01fF
C1295 VDD.n700 GND 0.00fF
C1296 VDD.n701 GND 0.00fF
C1297 VDD.n702 GND 0.02fF
C1298 VDD.n703 GND 0.01fF
C1299 VDD.n704 GND 0.03fF
C1300 VDD.n706 GND 0.01fF
C1301 VDD.n708 GND 0.00fF
C1302 VDD.n709 GND 0.00fF
C1303 VDD.n710 GND 0.00fF
C1304 VDD.n711 GND 0.00fF
C1305 VDD.n712 GND 0.00fF
C1306 VDD.n713 GND 0.00fF
C1307 VDD.n714 GND 0.01fF
C1308 VDD.n715 GND 0.01fF
C1309 VDD.n717 GND 0.00fF
C1310 VDD.n718 GND 0.00fF
C1311 VDD.n719 GND 0.00fF
C1312 VDD.n720 GND 0.00fF
C1313 VDD.n721 GND 0.00fF
C1314 VDD.n722 GND 0.00fF
C1315 VDD.n723 GND 0.01fF
C1316 VDD.n724 GND 0.00fF
C1317 VDD.n725 GND 0.00fF
C1318 VDD.n726 GND 0.00fF
C1319 VDD.n727 GND 0.00fF
C1320 VDD.n728 GND 0.00fF
C1321 VDD.n729 GND 0.01fF
C1322 VDD.n730 GND 0.01fF
C1323 VDD.n731 GND 0.00fF
C1324 VDD.n733 GND 0.00fF
C1325 VDD.n734 GND 0.00fF
C1326 VDD.n735 GND 0.00fF
C1327 VDD.n736 GND 0.00fF
C1328 VDD.n737 GND 0.00fF
C1329 VDD.n738 GND 0.01fF
C1330 VDD.n739 GND 0.01fF
C1331 VDD.n740 GND 0.00fF
C1332 VDD.n742 GND 0.35fF
C1333 VDD.n743 GND 0.02fF
C1334 VDD.n744 GND 0.01fF
C1335 VDD.n745 GND 0.01fF
C1336 VDD.n746 GND 0.00fF
C1337 VDD.n747 GND 0.00fF
C1338 VDD.n748 GND 0.00fF
C1339 VDD.n749 GND 0.01fF
C1340 VDD.n750 GND 0.01fF
C1341 VDD.n751 GND 0.03fF
C1342 VDD.n752 GND 0.01fF
C1343 VDD.n753 GND 0.01fF
C1344 VDD.n754 GND 0.00fF
C1345 VDD.n755 GND 0.00fF
C1346 VDD.n756 GND 0.00fF
C1347 VDD.n757 GND 0.00fF
C1348 VDD.n758 GND 0.00fF
C1349 VDD.n759 GND 0.00fF
C1350 VDD.n760 GND 0.00fF
C1351 VDD.n761 GND 0.00fF
C1352 VDD.n762 GND 0.00fF
C1353 VDD.n763 GND 0.00fF
C1354 VDD.n764 GND 0.00fF
C1355 VDD.n765 GND 0.00fF
C1356 VDD.n766 GND 0.00fF
C1357 VDD.n767 GND 0.00fF
C1358 VDD.n768 GND 0.00fF
C1359 VDD.n769 GND 0.00fF
C1360 VDD.n770 GND 0.00fF
C1361 VDD.n771 GND 0.00fF
C1362 VDD.n772 GND 0.00fF
C1363 VDD.n773 GND 0.00fF
C1364 VDD.n774 GND 0.00fF
C1365 VDD.n775 GND 0.00fF
C1366 VDD.n776 GND 0.00fF
C1367 VDD.n777 GND 0.00fF
C1368 VDD.n778 GND 0.00fF
C1369 VDD.n779 GND 0.00fF
C1370 VDD.n780 GND 0.00fF
C1371 VDD.n781 GND 0.00fF
C1372 VDD.n782 GND 0.00fF
C1373 VDD.n783 GND 0.00fF
C1374 VDD.n784 GND 0.00fF
C1375 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/DRAIN GND 0.00fF
C1376 VDD.n785 GND 0.01fF
C1377 VDD.n786 GND 0.01fF
C1378 VDD.n787 GND 0.01fF
C1379 VDD.n788 GND 0.02fF
C1380 VDD.n789 GND 0.02fF
C1381 VDD.n790 GND 0.01fF
C1382 VDD.n791 GND 0.01fF
C1383 VDD.n792 GND 0.02fF
C1384 VDD.n793 GND 0.02fF
C1385 VDD.n794 GND 0.01fF
C1386 VDD.n795 GND 0.03fF
C1387 VDD.n796 GND 0.03fF
C1388 VDD.n797 GND 0.04fF
C1389 VDD.n798 GND 0.00fF
C1390 VDD.n799 GND 0.00fF
C1391 VDD.n800 GND 0.00fF
C1392 VDD.n801 GND 0.00fF
C1393 VDD.n802 GND 0.00fF
C1394 VDD.n803 GND 0.01fF
C1395 VDD.n804 GND 0.00fF
C1396 VDD.n805 GND 0.01fF
C1397 VDD.n806 GND 0.00fF
C1398 VDD.n807 GND 0.00fF
C1399 VDD.n808 GND 0.00fF
C1400 VDD.n809 GND 0.00fF
C1401 VDD.n810 GND 0.01fF
C1402 VDD.n811 GND 0.00fF
C1403 VDD.n812 GND 0.01fF
C1404 VDD.n813 GND 0.00fF
C1405 VDD.n814 GND 0.00fF
C1406 VDD.n815 GND 0.00fF
C1407 VDD.n816 GND 0.00fF
C1408 VDD.n817 GND 0.01fF
C1409 VDD.n818 GND 0.00fF
C1410 VDD.n819 GND 0.01fF
C1411 VDD.n820 GND 0.00fF
C1412 VDD.n821 GND 0.00fF
C1413 VDD.n822 GND 0.00fF
C1414 VDD.n823 GND 0.00fF
C1415 VDD.n824 GND 0.01fF
C1416 VDD.n825 GND 0.00fF
C1417 VDD.n826 GND 0.01fF
C1418 VDD.n827 GND 0.00fF
C1419 VDD.n828 GND 0.00fF
C1420 VDD.t19 GND 0.04fF $ **FLOATING
C1421 VDD.n829 GND 0.07fF
C1422 VDD.n830 GND 0.01fF
C1423 VDD.n831 GND 0.01fF
C1424 VDD.n832 GND 0.01fF
C1425 VDD.n833 GND 0.00fF
C1426 VDD.n834 GND 0.01fF
C1427 VDD.n835 GND 0.03fF
C1428 VDD.n836 GND 0.07fF
C1429 VDD.n837 GND 0.37fF
C1430 VDD.n839 GND 0.10fF
C1431 VDD.n840 GND 0.03fF
C1432 VDD.n841 GND 0.02fF
C1433 VDD.n842 GND 0.03fF
C1434 VDD.n843 GND 0.00fF
C1435 VDD.n844 GND 0.01fF
C1436 VDD.n845 GND 0.01fF
C1437 VDD.n846 GND 0.01fF
C1438 VDD.n847 GND 0.03fF
C1439 VDD.n848 GND 0.01fF
C1440 VDD.n849 GND 0.00fF
C1441 VDD.n850 GND 0.01fF
C1442 VDD.n851 GND 0.01fF
C1443 VDD.n852 GND 0.05fF
C1444 VDD.n854 GND 0.05fF
C1445 VDD.n855 GND 0.04fF
C1446 VDD.n856 GND 0.04fF
C1447 VDD.n857 GND 0.01fF
C1448 VDD.n858 GND 0.00fF
C1449 VDD.n859 GND 0.00fF
C1450 VDD.n860 GND 0.01fF
C1451 VDD.n861 GND 0.01fF
C1452 VDD.n862 GND 0.01fF
C1453 VDD.n863 GND 0.01fF
C1454 VDD.n864 GND 0.03fF
C1455 VDD.n865 GND 0.01fF
C1456 VDD.n866 GND 0.00fF
C1457 VDD.n867 GND 0.01fF
C1458 VDD.n868 GND 0.01fF
C1459 VDD.n869 GND 0.02fF
C1460 VDD.n870 GND 0.03fF
C1461 VDD.n871 GND 0.05fF
C1462 VDD.n872 GND 0.03fF
C1463 VDD.n873 GND 0.00fF
C1464 VDD.n874 GND 0.01fF
C1465 VDD.n875 GND 0.01fF
C1466 VDD.n876 GND 0.01fF
C1467 VDD.n877 GND 0.01fF
C1468 VDD.n878 GND 0.03fF
C1469 VDD.n879 GND 0.01fF
C1470 VDD.n880 GND 0.03fF
C1471 VDD.n881 GND 0.01fF
C1472 VDD.n882 GND 0.01fF
C1473 VDD.n883 GND 0.01fF
C1474 VDD.n884 GND 0.00fF
C1475 VDD.n885 GND 0.00fF
C1476 VDD.n886 GND 0.01fF
C1477 VDD.n887 GND 0.01fF
C1478 VDD.n888 GND 0.04fF
C1479 VDD.n889 GND 0.04fF
C1480 VDD.n890 GND 0.05fF
C1481 VDD.n891 GND 0.10fF
C1482 VDD.n893 GND 1.52fF
C1483 VDD.n894 GND 1.53fF
C1484 VDD.n895 GND 0.07fF
C1485 VDD.n896 GND 0.03fF
C1486 VDD.n897 GND 0.01fF
C1487 VDD.n898 GND 0.05fF
C1488 VDD.n899 GND 0.02fF
C1489 VDD.n900 GND 0.00fF
C1490 VDD.n901 GND 0.01fF
C1491 VDD.n902 GND 0.01fF
C1492 VDD.n903 GND 0.05fF
C1493 VDD.n905 GND 0.02fF
C1494 VDD.n906 GND 0.03fF
C1495 VDD.n907 GND 0.00fF
C1496 VDD.n908 GND 0.01fF
C1497 VDD.n909 GND 0.01fF
C1498 VDD.n910 GND 0.01fF
C1499 VDD.n911 GND 0.04fF
C1500 VDD.n912 GND 0.01fF
C1501 VDD.n913 GND 0.00fF
C1502 VDD.n914 GND 0.01fF
C1503 VDD.n915 GND 0.01fF
C1504 VDD.n916 GND 0.02fF
C1505 VDD.n917 GND 0.03fF
C1506 VDD.n918 GND 0.05fF
C1507 VDD.n919 GND 0.10fF
C1508 VDD.n920 GND 0.05fF
C1509 VDD.n921 GND 0.01fF
C1510 VDD.n922 GND 0.02fF
C1511 VDD.n923 GND 0.02fF
C1512 VDD.n924 GND 0.02fF
C1513 VDD.n925 GND 0.01fF
C1514 VDD.n927 GND 0.02fF
C1515 VDD.n928 GND 0.01fF
C1516 VDD.n929 GND 0.01fF
C1517 VDD.n930 GND 0.01fF
C1518 VDD.n931 GND 0.00fF
C1519 VDD.n932 GND 0.00fF
C1520 VDD.n933 GND 0.00fF
C1521 VDD.n934 GND 0.01fF
C1522 VDD.n935 GND 0.01fF
C1523 VDD.n936 GND 0.00fF
C1524 VDD.n937 GND 0.00fF
C1525 VDD.n938 GND 0.00fF
C1526 VDD.n939 GND 0.00fF
C1527 VDD.n940 GND 0.00fF
C1528 VDD.n941 GND 0.00fF
C1529 VDD.n942 GND 0.00fF
C1530 VDD.n943 GND 0.00fF
C1531 VDD.n944 GND 0.00fF
C1532 VDD.n945 GND 0.00fF
C1533 VDD.n946 GND 0.00fF
C1534 VDD.n947 GND 0.00fF
C1535 VDD.n948 GND 0.00fF
C1536 VDD.n949 GND 0.00fF
C1537 VDD.n950 GND 0.00fF
C1538 VDD.n951 GND 0.00fF
C1539 VDD.n952 GND 0.00fF
C1540 VDD.n953 GND 0.00fF
C1541 VDD.n954 GND 0.00fF
C1542 VDD.n955 GND 0.00fF
C1543 VDD.n956 GND 0.00fF
C1544 VDD.n957 GND 0.00fF
C1545 VDD.n958 GND 0.00fF
C1546 VDD.n959 GND 0.00fF
C1547 VDD.n960 GND 0.00fF
C1548 VDD.n961 GND 0.00fF
C1549 VDD.n962 GND 0.00fF
C1550 VDD.n963 GND 0.00fF
C1551 VDD.n964 GND 0.00fF
C1552 VDD.n965 GND 0.00fF
C1553 VDD.n966 GND 0.00fF
C1554 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/DRAIN GND 0.00fF
C1555 VDD.n967 GND 0.01fF
C1556 VDD.n968 GND 0.01fF
C1557 VDD.n969 GND 0.01fF
C1558 VDD.n970 GND 0.02fF
C1559 VDD.n971 GND 0.02fF
C1560 VDD.n972 GND 0.01fF
C1561 VDD.n973 GND 0.01fF
C1562 VDD.n974 GND 0.02fF
C1563 VDD.n975 GND 0.02fF
C1564 VDD.n976 GND 0.01fF
C1565 VDD.n977 GND 0.03fF
C1566 VDD.n978 GND 0.03fF
C1567 VDD.n979 GND 0.04fF
C1568 VDD.n980 GND 0.00fF
C1569 VDD.n981 GND 0.00fF
C1570 VDD.n982 GND 0.00fF
C1571 VDD.n983 GND 0.00fF
C1572 VDD.n984 GND 0.00fF
C1573 VDD.n985 GND 0.01fF
C1574 VDD.n986 GND 0.00fF
C1575 VDD.n987 GND 0.01fF
C1576 VDD.n988 GND 0.00fF
C1577 VDD.n989 GND 0.00fF
C1578 VDD.n990 GND 0.00fF
C1579 VDD.n991 GND 0.00fF
C1580 VDD.n992 GND 0.01fF
C1581 VDD.n993 GND 0.00fF
C1582 VDD.n994 GND 0.01fF
C1583 VDD.n995 GND 0.00fF
C1584 VDD.n996 GND 0.00fF
C1585 VDD.n997 GND 0.00fF
C1586 VDD.n998 GND 0.00fF
C1587 VDD.n999 GND 0.01fF
C1588 VDD.n1000 GND 0.00fF
C1589 VDD.n1001 GND 0.01fF
C1590 VDD.n1002 GND 0.00fF
C1591 VDD.n1003 GND 0.00fF
C1592 VDD.n1004 GND 0.00fF
C1593 VDD.n1005 GND 0.00fF
C1594 VDD.n1006 GND 0.01fF
C1595 VDD.n1007 GND 0.00fF
C1596 VDD.n1008 GND 0.01fF
C1597 VDD.n1009 GND 0.00fF
C1598 VDD.n1010 GND 0.00fF
C1599 VDD.t35 GND 0.04fF $ **FLOATING
C1600 VDD.n1011 GND 0.07fF
C1601 VDD.n1012 GND 0.01fF
C1602 VDD.n1013 GND 0.01fF
C1603 VDD.n1014 GND 0.00fF
C1604 VDD.n1015 GND 0.00fF
C1605 VDD.n1016 GND 0.00fF
C1606 VDD.n1017 GND 0.01fF
C1607 VDD.n1018 GND 0.01fF
C1608 VDD.n1019 GND 0.00fF
C1609 VDD.n1020 GND 0.00fF
C1610 VDD.n1021 GND 0.00fF
C1611 VDD.n1022 GND 0.01fF
C1612 VDD.n1023 GND 0.00fF
C1613 VDD.n1024 GND 0.00fF
C1614 VDD.n1025 GND 0.01fF
C1615 VDD.n1026 GND 0.00fF
C1616 VDD.n1027 GND 0.00fF
C1617 VDD.n1028 GND 0.00fF
C1618 VDD.n1029 GND 0.01fF
C1619 VDD.n1030 GND 0.00fF
C1620 VDD.n1031 GND 0.00fF
C1621 VDD.n1032 GND 0.01fF
C1622 VDD.n1033 GND 0.00fF
C1623 VDD.n1034 GND 0.00fF
C1624 VDD.n1035 GND 0.00fF
C1625 VDD.n1036 GND 0.01fF
C1626 VDD.n1037 GND 0.00fF
C1627 VDD.n1038 GND 0.00fF
C1628 VDD.n1039 GND 0.01fF
C1629 VDD.n1040 GND 0.00fF
C1630 VDD.n1041 GND 0.00fF
C1631 VDD.n1042 GND 0.00fF
C1632 VDD.n1043 GND 0.01fF
C1633 VDD.n1044 GND 0.00fF
C1634 VDD.n1045 GND 0.00fF
C1635 VDD.n1046 GND 0.01fF
C1636 VDD.n1047 GND 0.00fF
C1637 VDD.n1048 GND 0.00fF
C1638 VDD.n1049 GND 0.00fF
C1639 VDD.n1050 GND 0.00fF
C1640 VDD.n1051 GND 0.00fF
C1641 VDD.n1052 GND 0.00fF
C1642 VDD.n1053 GND 0.00fF
C1643 VDD.n1054 GND 0.00fF
C1644 VDD.n1055 GND 0.00fF
C1645 VDD.n1056 GND 0.00fF
C1646 VDD.n1057 GND 0.00fF
C1647 VDD.n1058 GND 0.00fF
C1648 VDD.n1059 GND 0.00fF
C1649 VDD.n1060 GND 0.00fF
C1650 VDD.n1061 GND 0.00fF
C1651 VDD.n1062 GND 0.00fF
C1652 VDD.n1063 GND 0.00fF
C1653 VDD.n1064 GND 0.00fF
C1654 VDD.n1065 GND 0.00fF
C1655 VDD.n1066 GND 0.00fF
C1656 VDD.n1067 GND 0.00fF
C1657 VDD.n1068 GND 0.00fF
C1658 VDD.n1069 GND 0.00fF
C1659 VDD.n1070 GND 0.00fF
C1660 VDD.n1071 GND 0.00fF
C1661 VDD.n1072 GND 0.00fF
C1662 VDD.n1073 GND 0.00fF
C1663 VDD.n1074 GND 0.00fF
C1664 VDD.n1075 GND 0.00fF
C1665 VDD.n1076 GND 0.00fF
C1666 VDD.n1077 GND 0.00fF
C1667 VDD.n1078 GND 0.00fF
C1668 VDD.n1079 GND 0.00fF
C1669 VDD.t36 GND 0.04fF $ **FLOATING
C1670 VDD.n1080 GND 0.11fF
C1671 VDD.n1081 GND 0.01fF
C1672 VDD.n1082 GND 0.00fF
C1673 VDD.n1083 GND 0.01fF
C1674 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/BULK GND 0.01fF
C1675 VDD.n1084 GND 0.01fF
C1676 VDD.n1085 GND 0.01fF
C1677 VDD.n1086 GND 0.00fF
C1678 VDD.n1088 GND 0.00fF
C1679 VDD.n1089 GND 0.00fF
C1680 VDD.n1090 GND 0.00fF
C1681 VDD.n1091 GND 0.00fF
C1682 VDD.n1092 GND 0.00fF
C1683 VDD.n1093 GND 0.01fF
C1684 VDD.n1094 GND 0.01fF
C1685 VDD.n1095 GND 0.00fF
C1686 VDD.n1097 GND 0.01fF
C1687 VDD.n1099 GND 0.00fF
C1688 VDD.n1100 GND 0.00fF
C1689 VDD.n1101 GND 0.00fF
C1690 VDD.n1102 GND 0.00fF
C1691 VDD.n1103 GND 0.00fF
C1692 VDD.n1104 GND 0.00fF
C1693 VDD.n1105 GND 0.01fF
C1694 VDD.n1106 GND 0.01fF
C1695 VDD.n1108 GND 0.00fF
C1696 VDD.n1109 GND 0.00fF
C1697 VDD.n1110 GND 0.00fF
C1698 VDD.n1111 GND 0.01fF
C1699 VDD.n1112 GND 0.00fF
C1700 VDD.n1113 GND 0.00fF
C1701 VDD.n1114 GND 0.02fF
C1702 VDD.n1119 GND 0.01fF
C1703 VDD.n1120 GND 0.02fF
C1704 VDD.n1122 GND 0.01fF
C1705 VDD.n1123 GND 0.02fF
C1706 VDD.n1125 GND 0.01fF
C1707 VDD.n1126 GND 0.03fF
C1708 VDD.n1127 GND 0.01fF
C1709 VDD.n1128 GND 0.02fF
C1710 VDD.n1130 GND 0.01fF
C1711 VDD.n1132 GND 0.00fF
C1712 VDD.n1133 GND 0.00fF
C1713 VDD.n1134 GND 0.00fF
C1714 VDD.n1135 GND 0.00fF
C1715 VDD.n1136 GND 0.00fF
C1716 VDD.n1137 GND 0.00fF
C1717 VDD.n1138 GND 0.01fF
C1718 VDD.n1139 GND 0.01fF
C1719 VDD.n1141 GND 0.00fF
C1720 VDD.n1142 GND 0.00fF
C1721 VDD.n1143 GND 0.00fF
C1722 VDD.n1144 GND 0.00fF
C1723 VDD.n1145 GND 0.00fF
C1724 VDD.n1146 GND 0.00fF
C1725 VDD.n1147 GND 0.01fF
C1726 VDD.n1148 GND 0.00fF
C1727 VDD.n1149 GND 0.00fF
C1728 VDD.n1150 GND 0.00fF
C1729 VDD.n1151 GND 0.00fF
C1730 VDD.n1152 GND 0.00fF
C1731 VDD.n1153 GND 0.01fF
C1732 VDD.n1154 GND 0.01fF
C1733 VDD.n1155 GND 0.00fF
C1734 VDD.n1157 GND 0.00fF
C1735 VDD.n1158 GND 0.00fF
C1736 VDD.n1159 GND 0.00fF
C1737 VDD.n1160 GND 0.00fF
C1738 VDD.n1161 GND 0.00fF
C1739 VDD.n1162 GND 0.01fF
C1740 VDD.n1163 GND 0.01fF
C1741 VDD.n1164 GND 0.00fF
C1742 VDD.n1166 GND 0.35fF
C1743 VDD.n1167 GND 0.02fF
C1744 VDD.n1168 GND 0.01fF
C1745 VDD.n1169 GND 0.00fF
C1746 VDD.n1170 GND 0.00fF
C1747 VDD.n1171 GND 0.00fF
C1748 VDD.n1172 GND 0.00fF
C1749 VDD.n1173 GND 0.01fF
C1750 VDD.n1174 GND 0.00fF
C1751 VDD.n1175 GND 0.00fF
C1752 VDD.n1176 GND 0.01fF
C1753 VDD.n1177 GND 0.01fF
C1754 VDD.n1178 GND 0.00fF
C1755 VDD.n1179 GND 0.01fF
C1756 VDD.n1180 GND 0.01fF
C1757 VDD.n1181 GND 0.00fF
C1758 VDD.n1182 GND 0.01fF
C1759 VDD.n1183 GND 0.01fF
C1760 VDD.n1184 GND 0.00fF
C1761 VDD.n1185 GND 0.01fF
C1762 VDD.n1186 GND 0.01fF
C1763 VDD.n1187 GND 0.00fF
C1764 VDD.n1188 GND 0.01fF
C1765 VDD.n1189 GND 0.01fF
C1766 VDD.n1190 GND 0.00fF
C1767 VDD.n1191 GND 0.01fF
C1768 VDD.n1192 GND 0.01fF
C1769 VDD.n1193 GND 0.00fF
C1770 VDD.n1194 GND 0.01fF
C1771 VDD.n1195 GND 0.01fF
C1772 VDD.n1196 GND 0.00fF
C1773 VDD.n1197 GND 0.01fF
C1774 VDD.t20 GND 0.04fF $ **FLOATING
C1775 VDD.n1198 GND 0.11fF
C1776 VDD.n1199 GND 0.01fF
C1777 VDD.n1200 GND 0.00fF
C1778 VDD.n1201 GND 0.00fF
C1779 VDD.n1202 GND 0.00fF
C1780 VDD.n1203 GND 0.00fF
C1781 VDD.n1204 GND 0.00fF
C1782 VDD.n1205 GND 0.00fF
C1783 VDD.n1206 GND 0.00fF
C1784 VDD.n1207 GND 0.00fF
C1785 VDD.n1208 GND 0.00fF
C1786 VDD.n1209 GND 0.00fF
C1787 VDD.n1210 GND 0.00fF
C1788 VDD.n1211 GND 0.00fF
C1789 VDD.n1212 GND 0.00fF
C1790 VDD.n1213 GND 0.00fF
C1791 VDD.n1214 GND 0.00fF
C1792 VDD.n1215 GND 0.00fF
C1793 VDD.n1216 GND 0.00fF
C1794 VDD.n1217 GND 0.00fF
C1795 VDD.n1218 GND 0.00fF
C1796 VDD.n1219 GND 0.00fF
C1797 VDD.n1220 GND 0.00fF
C1798 VDD.n1221 GND 0.00fF
C1799 VDD.n1222 GND 0.00fF
C1800 VDD.n1223 GND 0.00fF
C1801 VDD.n1224 GND 0.00fF
C1802 VDD.n1225 GND 0.00fF
C1803 VDD.n1226 GND 0.00fF
C1804 VDD.n1227 GND 0.00fF
C1805 VDD.n1228 GND 0.00fF
C1806 VDD.n1229 GND 0.00fF
C1807 VDD.n1230 GND 0.00fF
C1808 VDD.n1231 GND 0.00fF
C1809 VDD.n1232 GND 0.00fF
C1810 VDD.n1233 GND 0.00fF
C1811 VDD.n1234 GND 0.00fF
C1812 VDD.n1235 GND 0.00fF
C1813 VDD.n1236 GND 0.00fF
C1814 VDD.n1237 GND 0.00fF
C1815 VDD.n1238 GND 0.00fF
C1816 VDD.n1239 GND 0.01fF
C1817 VDD.n1240 GND 0.00fF
C1818 VDD.n1241 GND 0.01fF
C1819 VDD.n1242 GND 0.00fF
C1820 VDD.n1243 GND 0.00fF
C1821 VDD.n1244 GND 0.00fF
C1822 VDD.n1245 GND 0.00fF
C1823 VDD.n1246 GND 0.01fF
C1824 VDD.n1247 GND 0.00fF
C1825 VDD.n1248 GND 0.01fF
C1826 VDD.n1249 GND 0.00fF
C1827 VDD.n1250 GND 0.00fF
C1828 VDD.n1251 GND 0.00fF
C1829 VDD.n1252 GND 0.00fF
C1830 VDD.n1253 GND 0.01fF
C1831 VDD.n1254 GND 0.00fF
C1832 VDD.n1255 GND 0.01fF
C1833 VDD.n1256 GND 0.00fF
C1834 VDD.n1257 GND 0.00fF
C1835 VDD.n1258 GND 0.00fF
C1836 VDD.n1259 GND 0.00fF
C1837 VDD.n1260 GND 0.01fF
C1838 VDD.n1261 GND 0.00fF
C1839 VDD.n1262 GND 0.01fF
C1840 VDD.n1263 GND 0.00fF
C1841 VDD.n1264 GND 0.00fF
C1842 VDD.n1265 GND 0.01fF
C1843 VDD.n1266 GND 0.01fF
C1844 VDD.n1267 GND 0.04fF
C1845 VDD.n1268 GND 0.01fF
C1846 VDD.n1269 GND 0.01fF
C1847 VDD.n1270 GND 0.01fF
C1848 VDD.n1271 GND 0.00fF
C1849 VDD.n1272 GND 0.00fF
C1850 VDD.n1273 GND 0.01fF
C1851 VDD.n1274 GND 0.00fF
C1852 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/GATE GND 0.04fF
C1853 VDD.n1275 GND 0.04fF
C1854 VDD.n1276 GND 0.02fF
C1855 VDD.n1277 GND 0.01fF
C1856 VDD.n1278 GND 0.02fF
C1857 VDD.n1279 GND 0.01fF
C1858 VDD.n1280 GND 0.07fF
C1859 VDD.n1281 GND 0.11fF
C1860 VDD.n1282 GND 0.01fF
C1861 VDD.n1283 GND 0.00fF
C1862 VDD.n1284 GND 0.02fF
C1863 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/SOURCE GND 0.01fF
C1864 VDD.n1285 GND 0.02fF
C1865 VDD.n1286 GND 0.01fF
C1866 VDD.n1287 GND 0.03fF
C1867 VDD.n1288 GND 0.03fF
C1868 VDD.n1289 GND 0.01fF
C1869 VDD.n1290 GND 0.02fF
C1870 VDD.n1291 GND 0.02fF
C1871 VDD.n1292 GND 0.01fF
C1872 VDD.n1293 GND 0.01fF
C1873 VDD.n1294 GND 0.02fF
C1874 VDD.n1295 GND 0.02fF
C1875 VDD.n1296 GND 0.01fF
C1876 VDD.n1297 GND 0.01fF
C1877 VDD.n1298 GND 0.00fF
C1878 VDD.n1299 GND 0.00fF
C1879 VDD.n1300 GND 0.00fF
C1880 VDD.n1301 GND 0.00fF
C1881 VDD.n1302 GND 0.00fF
C1882 VDD.n1303 GND 0.00fF
C1883 VDD.n1304 GND 0.00fF
C1884 VDD.n1305 GND 0.00fF
C1885 VDD.n1306 GND 0.00fF
C1886 VDD.n1307 GND 0.00fF
C1887 VDD.n1308 GND 0.00fF
C1888 VDD.n1309 GND 0.00fF
C1889 VDD.n1310 GND 0.00fF
C1890 VDD.n1311 GND 0.00fF
C1891 VDD.n1312 GND 0.00fF
C1892 VDD.n1313 GND 0.00fF
C1893 VDD.n1314 GND 0.00fF
C1894 VDD.n1315 GND 0.00fF
C1895 VDD.n1316 GND 0.00fF
C1896 VDD.n1317 GND 0.00fF
C1897 VDD.n1318 GND 0.00fF
C1898 VDD.n1319 GND 0.00fF
C1899 VDD.n1320 GND 0.00fF
C1900 VDD.n1321 GND 0.00fF
C1901 VDD.n1322 GND 0.00fF
C1902 VDD.n1323 GND 0.00fF
C1903 VDD.n1324 GND 0.00fF
C1904 VDD.n1325 GND 0.00fF
C1905 VDD.n1326 GND 0.00fF
C1906 VDD.n1327 GND 0.00fF
C1907 VDD.n1328 GND 0.00fF
C1908 VDD.n1329 GND 0.00fF
C1909 VDD.n1330 GND 0.00fF
C1910 VDD.n1331 GND 0.00fF
C1911 VDD.n1332 GND 0.00fF
C1912 VDD.n1333 GND 0.00fF
C1913 VDD.n1334 GND 0.00fF
C1914 VDD.n1335 GND 0.00fF
C1915 VDD.n1336 GND 0.01fF
C1916 VDD.n1337 GND 0.00fF
C1917 VDD.n1338 GND 0.01fF
C1918 VDD.n1339 GND 0.00fF
C1919 VDD.n1340 GND 0.00fF
C1920 VDD.n1341 GND 0.00fF
C1921 VDD.n1342 GND 0.00fF
C1922 VDD.n1343 GND 0.01fF
C1923 VDD.n1344 GND 0.00fF
C1924 VDD.n1345 GND 0.01fF
C1925 VDD.n1346 GND 0.00fF
C1926 VDD.n1347 GND 0.00fF
C1927 VDD.n1348 GND 0.00fF
C1928 VDD.n1349 GND 0.00fF
C1929 VDD.n1350 GND 0.01fF
C1930 VDD.n1351 GND 0.00fF
C1931 VDD.n1352 GND 0.01fF
C1932 VDD.n1353 GND 0.00fF
C1933 VDD.n1354 GND 0.00fF
C1934 VDD.n1355 GND 0.00fF
C1935 VDD.n1356 GND 0.00fF
C1936 VDD.n1357 GND 0.01fF
C1937 VDD.n1358 GND 0.00fF
C1938 VDD.n1359 GND 0.01fF
C1939 VDD.n1360 GND 0.00fF
C1940 VDD.n1361 GND 0.00fF
C1941 VDD.n1362 GND 0.01fF
C1942 VDD.n1363 GND 0.01fF
C1943 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/BULK GND 0.01fF
C1944 VDD.n1364 GND 0.01fF
C1945 VDD.n1365 GND 0.00fF
C1946 VDD.n1366 GND 0.00fF
C1947 VDD.n1367 GND 0.00fF
C1948 VDD.n1368 GND 0.00fF
C1949 VDD.n1369 GND 0.00fF
C1950 VDD.n1370 GND 0.01fF
C1951 VDD.n1371 GND 0.00fF
C1952 VDD.n1373 GND 0.01fF
C1953 VDD.n1374 GND 0.00fF
C1954 VDD.n1375 GND 0.01fF
C1955 VDD.n1376 GND 0.00fF
C1956 VDD.n1377 GND 0.01fF
C1957 VDD.n1378 GND 0.00fF
C1958 VDD.n1379 GND 0.00fF
C1959 VDD.n1380 GND 0.00fF
C1960 VDD.n1381 GND 0.00fF
C1961 VDD.n1382 GND 0.01fF
C1962 VDD.n1383 GND 0.00fF
C1963 VDD.n1385 GND 0.01fF
C1964 VDD.n1386 GND 0.00fF
C1965 VDD.n1387 GND 0.01fF
C1966 VDD.n1388 GND 0.00fF
C1967 VDD.n1389 GND 0.01fF
C1968 VDD.n1390 GND 0.00fF
C1969 VDD.n1391 GND 0.00fF
C1970 VDD.n1392 GND 0.00fF
C1971 VDD.n1393 GND 0.00fF
C1972 VDD.n1394 GND 0.01fF
C1973 VDD.n1395 GND 0.00fF
C1974 VDD.n1397 GND 0.01fF
C1975 VDD.n1398 GND 0.00fF
C1976 VDD.n1399 GND 0.01fF
C1977 VDD.n1400 GND 0.00fF
C1978 VDD.n1401 GND 0.01fF
C1979 VDD.n1402 GND 0.00fF
C1980 VDD.n1403 GND 0.00fF
C1981 VDD.n1404 GND 0.00fF
C1982 VDD.n1405 GND 0.00fF
C1983 VDD.n1406 GND 0.01fF
C1984 VDD.n1407 GND 0.00fF
C1985 VDD.n1409 GND 0.01fF
C1986 VDD.n1410 GND 0.00fF
C1987 VDD.n1411 GND 0.01fF
C1988 VDD.n1412 GND 0.00fF
C1989 VDD.n1413 GND 0.00fF
C1990 VDD.n1414 GND 0.01fF
C1991 VDD.n1416 GND 0.00fF
C1992 VDD.n1417 GND 0.01fF
C1993 VDD.n1418 GND 0.00fF
C1994 VDD.n1419 GND 0.01fF
C1995 VDD.n1420 GND 0.00fF
C1996 VDD.n1421 GND 0.00fF
C1997 VDD.n1422 GND 0.00fF
C1998 VDD.n1423 GND 0.01fF
C1999 VDD.n1424 GND 0.00fF
C2000 VDD.n1425 GND 0.00fF
C2001 VDD.n1426 GND 0.01fF
C2002 VDD.n1428 GND 0.00fF
C2003 VDD.n1429 GND 0.01fF
C2004 VDD.n1430 GND 0.00fF
C2005 VDD.n1431 GND 0.01fF
C2006 VDD.n1432 GND 0.00fF
C2007 VDD.n1433 GND 0.00fF
C2008 VDD.n1434 GND 0.00fF
C2009 VDD.n1435 GND 0.01fF
C2010 VDD.n1436 GND 0.00fF
C2011 VDD.n1437 GND 0.00fF
C2012 VDD.n1438 GND 0.01fF
C2013 VDD.n1440 GND 0.00fF
C2014 VDD.n1441 GND 0.01fF
C2015 VDD.n1442 GND 0.00fF
C2016 VDD.n1443 GND 0.01fF
C2017 VDD.n1444 GND 0.00fF
C2018 VDD.n1445 GND 0.00fF
C2019 VDD.n1446 GND 0.00fF
C2020 VDD.n1447 GND 0.01fF
C2021 VDD.n1448 GND 0.00fF
C2022 VDD.n1449 GND 0.00fF
C2023 VDD.n1450 GND 0.01fF
C2024 VDD.n1452 GND 0.00fF
C2025 VDD.n1453 GND 0.01fF
C2026 VDD.n1454 GND 0.00fF
C2027 VDD.n1455 GND 0.01fF
C2028 VDD.n1456 GND 0.00fF
C2029 VDD.n1457 GND 0.00fF
C2030 VDD.n1458 GND 0.01fF
C2031 VDD.n1459 GND 0.01fF
C2032 VDD.n1460 GND 0.03fF
C2033 VDD.n1461 GND 0.02fF
C2034 VDD.n1462 GND 0.03fF
C2035 VDD.n1463 GND 0.03fF
C2036 VDD.n1464 GND 0.02fF
C2037 VDD.n1465 GND 0.05fF
C2038 VDD.n1466 GND 0.04fF
C2039 VDD.n1467 GND 0.02fF
C2040 VDD.n1468 GND 0.01fF
C2041 VDD.n1469 GND 0.00fF
C2042 VDD.n1470 GND 0.00fF
C2043 VDD.n1471 GND 0.00fF
C2044 VDD.n1472 GND 0.04fF
C2045 VDD.n1473 GND 0.01fF
C2046 VDD.n1474 GND 0.01fF
C2047 VDD.n1475 GND 0.02fF
C2048 VDD.n1476 GND 0.02fF
C2049 VDD.n1477 GND 0.01fF
C2050 VDD.n1478 GND 0.02fF
C2051 VDD.n1479 GND 0.01fF
C2052 VDD.n1480 GND 0.01fF
C2053 VDD.n1481 GND 0.03fF
C2054 VDD.n1482 GND 0.04fF
C2055 VDD.n1483 GND 0.01fF
C2056 VDD.n1484 GND 0.01fF
C2057 VDD.n1485 GND 0.02fF
C2058 VDD.n1486 GND 0.00fF
C2059 VDD.n1487 GND 0.00fF
C2060 VDD.n1488 GND 0.02fF
C2061 VDD.n1489 GND 0.01fF
C2062 VDD.n1490 GND 0.00fF
C2063 VDD.n1491 GND 0.02fF
C2064 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_7/GATE GND 0.04fF
C2065 VDD.n1492 GND 0.02fF
C2066 VDD.n1493 GND 0.01fF
C2067 VDD.n1494 GND 0.03fF
C2068 VDD.n1495 GND 0.02fF
C2069 VDD.n1496 GND 0.01fF
C2070 VDD.n1497 GND 0.02fF
C2071 VDD.n1498 GND 0.02fF
C2072 VDD.n1499 GND 0.01fF
C2073 VDD.n1500 GND 0.02fF
C2074 VDD.n1501 GND 0.02fF
C2075 VDD.n1502 GND 0.01fF
C2076 VDD.n1503 GND 0.02fF
C2077 VDD.n1504 GND 0.01fF
C2078 VDD.n1505 GND 0.02fF
C2079 VDD.n1506 GND 0.02fF
C2080 VDD.n1507 GND 0.01fF
C2081 VDD.n1508 GND 0.02fF
C2082 VDD.n1509 GND 0.03fF
C2083 VDD.n1510 GND 0.01fF
C2084 VDD.n1511 GND 0.01fF
C2085 VDD.n1512 GND 0.01fF
C2086 VDD.n1513 GND 0.00fF
C2087 VDD.n1514 GND 0.00fF
C2088 VDD.n1515 GND 0.00fF
C2089 VDD.n1516 GND 0.00fF
C2090 VDD.n1517 GND 0.01fF
C2091 VDD.n1519 GND 0.00fF
C2092 VDD.n1520 GND 0.01fF
C2093 VDD.n1521 GND 0.00fF
C2094 VDD.n1522 GND 0.01fF
C2095 VDD.n1523 GND 0.00fF
C2096 VDD.n1524 GND 0.01fF
C2097 VDD.n1525 GND 0.00fF
C2098 VDD.n1526 GND 0.00fF
C2099 VDD.n1527 GND 0.00fF
C2100 VDD.n1528 GND 0.00fF
C2101 VDD.n1529 GND 0.01fF
C2102 VDD.n1530 GND 0.00fF
C2103 VDD.n1532 GND 0.01fF
C2104 VDD.n1533 GND 0.00fF
C2105 VDD.n1534 GND 0.01fF
C2106 VDD.n1535 GND 0.00fF
C2107 VDD.n1536 GND 0.01fF
C2108 VDD.n1537 GND 0.00fF
C2109 VDD.n1538 GND 0.00fF
C2110 VDD.n1539 GND 0.00fF
C2111 VDD.n1540 GND 0.00fF
C2112 VDD.n1541 GND 0.01fF
C2113 VDD.n1543 GND 0.00fF
C2114 VDD.n1544 GND 0.01fF
C2115 VDD.n1545 GND 0.00fF
C2116 VDD.n1546 GND 0.01fF
C2117 VDD.n1547 GND 0.00fF
C2118 VDD.n1548 GND 0.01fF
C2119 VDD.n1549 GND 0.00fF
C2120 VDD.n1550 GND 0.00fF
C2121 VDD.n1551 GND 0.00fF
C2122 VDD.n1552 GND 0.00fF
C2123 VDD.n1554 GND 0.01fF
C2124 VDD.n1555 GND 0.00fF
C2125 VDD.n1557 GND 0.01fF
C2126 VDD.n1558 GND 0.00fF
C2127 VDD.n1559 GND 0.01fF
C2128 VDD.n1560 GND 0.00fF
C2129 VDD.n1561 GND 0.00fF
C2130 VDD.n1562 GND 0.01fF
C2131 VDD.n1563 GND 0.00fF
C2132 VDD.n1565 GND 0.01fF
C2133 VDD.n1566 GND 0.00fF
C2134 VDD.n1567 GND 0.01fF
C2135 VDD.n1568 GND 0.00fF
C2136 VDD.n1569 GND 0.00fF
C2137 VDD.n1570 GND 0.00fF
C2138 VDD.n1571 GND 0.01fF
C2139 VDD.n1572 GND 0.00fF
C2140 VDD.n1573 GND 0.00fF
C2141 VDD.n1574 GND 0.01fF
C2142 VDD.n1576 GND 0.00fF
C2143 VDD.n1577 GND 0.01fF
C2144 VDD.n1578 GND 0.00fF
C2145 VDD.n1579 GND 0.01fF
C2146 VDD.n1580 GND 0.00fF
C2147 VDD.n1581 GND 0.00fF
C2148 VDD.n1582 GND 0.00fF
C2149 VDD.n1583 GND 0.01fF
C2150 VDD.n1584 GND 0.00fF
C2151 VDD.n1585 GND 0.00fF
C2152 VDD.n1586 GND 0.01fF
C2153 VDD.n1587 GND 0.00fF
C2154 VDD.n1589 GND 0.01fF
C2155 VDD.n1590 GND 0.00fF
C2156 VDD.n1591 GND 0.01fF
C2157 VDD.n1592 GND 0.00fF
C2158 VDD.n1593 GND 0.00fF
C2159 VDD.n1594 GND 0.00fF
C2160 VDD.n1595 GND 0.01fF
C2161 VDD.n1596 GND 0.00fF
C2162 VDD.n1597 GND 0.00fF
C2163 VDD.n1598 GND 0.01fF
C2164 VDD.n1600 GND 0.00fF
C2165 VDD.n1601 GND 0.01fF
C2166 VDD.n1602 GND 0.00fF
C2167 VDD.n1603 GND 0.01fF
C2168 VDD.n1604 GND 0.00fF
C2169 VDD.n1605 GND 0.00fF
C2170 VDD.n1606 GND 0.01fF
C2171 VDD.n1607 GND 0.00fF
C2172 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/BULK GND 0.01fF
C2173 VDD.n1608 GND 0.01fF
C2174 VDD.n1609 GND 0.02fF
C2175 VDD.n1610 GND 0.00fF
C2176 VDD.n1611 GND 0.01fF
C2177 VDD.n1612 GND 0.00fF
C2178 VDD.n1613 GND 0.00fF
C2179 VDD.t34 GND 0.04fF $ **FLOATING
C2180 VDD.n1614 GND 0.04fF
C2181 VDD.n1615 GND 0.01fF
C2182 VDD.n1616 GND 0.01fF
C2183 VDD.n1617 GND 0.01fF
C2184 VDD.n1618 GND 0.01fF
C2185 VDD.n1619 GND 0.01fF
C2186 VDD.n1620 GND 0.03fF
C2187 VDD.t21 GND 0.04fF $ **FLOATING
C2188 VDD.n1621 GND 0.04fF
C2189 VDD.n1622 GND 0.01fF
C2190 VDD.n1623 GND 0.01fF
C2191 VDD.n1624 GND 0.01fF
C2192 VDD.n1625 GND 0.00fF
C2193 VDD.n1626 GND 0.00fF
C2194 VDD.n1627 GND 0.01fF
C2195 VDD.n1628 GND 0.02fF
C2196 VDD.n1629 GND 0.03fF
C2197 VDD.n1631 GND 0.02fF
C2198 VDD.n1632 GND 0.01fF
C2199 VDD.n1633 GND 0.01fF
C2200 VDD.n1635 GND 0.02fF
C2201 VDD.n1636 GND 0.01fF
C2202 VDD.n1637 GND 0.02fF
C2203 VDD.n1638 GND 0.07fF
C2204 VDD.n1639 GND 0.11fF
C2205 VDD.n1640 GND 0.01fF
C2206 VDD.n1641 GND 0.00fF
C2207 VDD.n1642 GND 0.02fF
C2208 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/SOURCE GND 0.01fF
C2209 VDD.n1643 GND 0.02fF
C2210 VDD.n1644 GND 0.01fF
C2211 VDD.n1645 GND 0.03fF
C2212 VDD.n1646 GND 0.03fF
C2213 VDD.n1647 GND 0.01fF
C2214 VDD.n1648 GND 0.02fF
C2215 VDD.n1649 GND 0.02fF
C2216 VDD.n1650 GND 0.01fF
C2217 VDD.n1651 GND 0.01fF
C2218 VDD.n1652 GND 0.02fF
C2219 VDD.n1653 GND 0.02fF
C2220 VDD.n1654 GND 0.01fF
C2221 VDD.n1655 GND 0.01fF
C2222 VDD.n1656 GND 0.00fF
C2223 VDD.n1657 GND 0.00fF
C2224 VDD.n1658 GND 0.00fF
C2225 VDD.n1659 GND 0.00fF
C2226 VDD.n1660 GND 0.00fF
C2227 VDD.n1661 GND 0.00fF
C2228 VDD.n1662 GND 0.00fF
C2229 VDD.n1663 GND 0.00fF
C2230 VDD.n1664 GND 0.00fF
C2231 VDD.n1665 GND 0.00fF
C2232 VDD.n1666 GND 0.00fF
C2233 VDD.n1667 GND 0.00fF
C2234 VDD.n1668 GND 0.00fF
C2235 VDD.n1669 GND 0.00fF
C2236 VDD.n1670 GND 0.00fF
C2237 VDD.n1671 GND 0.00fF
C2238 VDD.n1672 GND 0.00fF
C2239 VDD.n1673 GND 0.00fF
C2240 VDD.n1674 GND 0.00fF
C2241 VDD.n1675 GND 0.00fF
C2242 VDD.n1676 GND 0.00fF
C2243 VDD.n1677 GND 0.00fF
C2244 VDD.n1678 GND 0.00fF
C2245 VDD.n1679 GND 0.00fF
C2246 VDD.n1680 GND 0.00fF
C2247 VDD.n1681 GND 0.00fF
C2248 VDD.n1682 GND 0.00fF
C2249 VDD.n1683 GND 0.00fF
C2250 VDD.n1684 GND 0.00fF
C2251 VDD.n1685 GND 0.00fF
C2252 VDD.n1686 GND 0.00fF
C2253 VDD.n1687 GND 0.00fF
C2254 VDD.n1688 GND 0.00fF
C2255 VDD.n1689 GND 0.00fF
C2256 VDD.n1690 GND 0.00fF
C2257 VDD.n1691 GND 0.00fF
C2258 VDD.n1692 GND 0.00fF
C2259 VDD.n1693 GND 0.00fF
C2260 VDD.n1694 GND 0.01fF
C2261 VDD.n1695 GND 0.00fF
C2262 VDD.n1696 GND 0.01fF
C2263 VDD.n1697 GND 0.00fF
C2264 VDD.n1698 GND 0.00fF
C2265 VDD.n1699 GND 0.00fF
C2266 VDD.n1700 GND 0.00fF
C2267 VDD.n1701 GND 0.01fF
C2268 VDD.n1702 GND 0.00fF
C2269 VDD.n1703 GND 0.01fF
C2270 VDD.n1704 GND 0.00fF
C2271 VDD.n1705 GND 0.00fF
C2272 VDD.n1706 GND 0.00fF
C2273 VDD.n1707 GND 0.00fF
C2274 VDD.n1708 GND 0.01fF
C2275 VDD.n1709 GND 0.00fF
C2276 VDD.n1710 GND 0.01fF
C2277 VDD.n1711 GND 0.00fF
C2278 VDD.n1712 GND 0.00fF
C2279 VDD.n1713 GND 0.00fF
C2280 VDD.n1714 GND 0.00fF
C2281 VDD.n1715 GND 0.01fF
C2282 VDD.n1716 GND 0.00fF
C2283 VDD.n1717 GND 0.01fF
C2284 VDD.n1718 GND 0.00fF
C2285 VDD.n1719 GND 0.00fF
C2286 VDD.n1720 GND 0.01fF
C2287 VDD.n1721 GND 0.01fF
C2288 VDD.n1722 GND 0.04fF
C2289 VDD.n1723 GND 0.01fF
C2290 VDD.n1724 GND 0.01fF
C2291 VDD.n1725 GND 0.01fF
C2292 VDD.n1726 GND 0.00fF
C2293 VDD.n1727 GND 0.00fF
C2294 VDD.n1728 GND 0.01fF
C2295 VDD.n1729 GND 0.02fF
C2296 VDD.n1730 GND 0.03fF
C2297 VDD.n1731 GND 0.01fF
C2298 VDD.n1732 GND 0.04fF
C2299 VDD.n1733 GND 0.01fF
C2300 VDD.n1734 GND 0.01fF
C2301 VDD.n1735 GND 0.00fF
C2302 VDD.n1736 GND 0.00fF
C2303 VDD.n1737 GND 0.00fF
C2304 VDD.n1738 GND 0.00fF
C2305 VDD.n1739 GND 0.01fF
C2306 VDD.n1741 GND 0.00fF
C2307 VDD.n1742 GND 0.02fF
C2308 VDD.n1743 GND 0.00fF
C2309 VDD.n1744 GND 0.01fF
C2310 VDD.n1745 GND 0.00fF
C2311 VDD.n1746 GND 0.01fF
C2312 VDD.n1747 GND 0.00fF
C2313 VDD.n1748 GND 0.00fF
C2314 VDD.n1749 GND 0.00fF
C2315 VDD.n1750 GND 0.00fF
C2316 VDD.n1751 GND 0.01fF
C2317 VDD.n1753 GND 0.00fF
C2318 VDD.n1754 GND 0.01fF
C2319 VDD.n1755 GND 0.00fF
C2320 VDD.n1756 GND 0.01fF
C2321 VDD.n1757 GND 0.00fF
C2322 VDD.n1758 GND 0.01fF
C2323 VDD.n1759 GND 0.00fF
C2324 VDD.n1760 GND 0.00fF
C2325 VDD.n1761 GND 0.00fF
C2326 VDD.n1762 GND 0.00fF
C2327 VDD.n1763 GND 0.01fF
C2328 VDD.n1765 GND 0.00fF
C2329 VDD.n1766 GND 0.01fF
C2330 VDD.n1767 GND 0.00fF
C2331 VDD.n1768 GND 0.01fF
C2332 VDD.n1769 GND 0.00fF
C2333 VDD.n1770 GND 0.01fF
C2334 VDD.n1771 GND 0.00fF
C2335 VDD.n1772 GND 0.00fF
C2336 VDD.n1773 GND 0.00fF
C2337 VDD.n1774 GND 0.00fF
C2338 VDD.n1775 GND 0.01fF
C2339 VDD.n1777 GND 0.00fF
C2340 VDD.n1778 GND 0.01fF
C2341 VDD.n1779 GND 0.00fF
C2342 VDD.n1780 GND 0.01fF
C2343 VDD.n1781 GND 0.00fF
C2344 VDD.n1782 GND 0.00fF
C2345 VDD.n1783 GND 0.01fF
C2346 VDD.n1784 GND 0.00fF
C2347 VDD.n1786 GND 0.01fF
C2348 VDD.n1787 GND 0.00fF
C2349 VDD.n1788 GND 0.01fF
C2350 VDD.n1789 GND 0.00fF
C2351 VDD.n1790 GND 0.00fF
C2352 VDD.n1791 GND 0.00fF
C2353 VDD.n1792 GND 0.01fF
C2354 VDD.n1793 GND 0.00fF
C2355 VDD.n1794 GND 0.00fF
C2356 VDD.n1795 GND 0.01fF
C2357 VDD.n1796 GND 0.00fF
C2358 VDD.n1798 GND 0.01fF
C2359 VDD.n1799 GND 0.00fF
C2360 VDD.n1800 GND 0.01fF
C2361 VDD.n1801 GND 0.00fF
C2362 VDD.n1802 GND 0.00fF
C2363 VDD.n1803 GND 0.00fF
C2364 VDD.n1804 GND 0.01fF
C2365 VDD.n1805 GND 0.00fF
C2366 VDD.n1806 GND 0.00fF
C2367 VDD.n1807 GND 0.01fF
C2368 VDD.n1808 GND 0.00fF
C2369 VDD.n1810 GND 0.01fF
C2370 VDD.n1811 GND 0.00fF
C2371 VDD.n1812 GND 0.01fF
C2372 VDD.n1813 GND 0.00fF
C2373 VDD.n1814 GND 0.00fF
C2374 VDD.n1815 GND 0.00fF
C2375 VDD.n1816 GND 0.01fF
C2376 VDD.n1817 GND 0.00fF
C2377 VDD.n1818 GND 0.00fF
C2378 VDD.n1819 GND 0.01fF
C2379 VDD.n1821 GND 0.00fF
C2380 VDD.n1822 GND 0.01fF
C2381 VDD.n1823 GND 0.00fF
C2382 VDD.n1824 GND 0.01fF
C2383 VDD.n1825 GND 0.00fF
C2384 VDD.n1826 GND 0.00fF
C2385 VDD.n1827 GND 0.01fF
C2386 VDD.n1828 GND 0.00fF
C2387 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_0/BULK GND 0.01fF
C2388 VDD.n1831 GND 0.72fF
C2389 VDD.n1833 GND 0.03fF
C2390 VDD.n1834 GND 0.02fF
C2391 VDD.n1835 GND 0.03fF
C2392 VDD.n1836 GND 0.50fF
C2393 VDD.n1837 GND 0.03fF
C2394 VDD.n1838 GND 0.02fF
C2395 VDD.n1839 GND 0.05fF
C2396 VDD.n1840 GND 0.04fF
C2397 VDD.t13 GND 0.35fF $ **FLOATING
C2398 VDD.n1841 GND 0.53fF
C2399 VDD.n1842 GND 0.02fF
C2400 VDD.n1843 GND 0.01fF
C2401 VDD.n1844 GND 0.00fF
C2402 VDD.n1845 GND 0.00fF
C2403 VDD.n1846 GND 0.00fF
C2404 VDD.t12 GND 0.04fF $ **FLOATING
C2405 VDD.n1847 GND 0.04fF
C2406 VDD.n1848 GND 0.01fF
C2407 VDD.n1849 GND 0.01fF
C2408 VDD.n1850 GND 0.01fF
C2409 VDD.n1851 GND 0.03fF
C2410 VDD.n1852 GND 0.38fF
C2411 VDD.n1853 GND 0.02fF
C2412 VDD.n1854 GND 0.01fF
C2413 VDD.n1855 GND 0.02fF
C2414 VDD.n1856 GND 0.01fF
C2415 VDD.n1857 GND 0.01fF
C2416 VDD.n1858 GND 0.03fF
C2417 VDD.t17 GND 0.04fF $ **FLOATING
C2418 VDD.n1859 GND 0.04fF
C2419 VDD.n1860 GND 0.01fF
C2420 VDD.n1861 GND 0.01fF
C2421 VDD.n1862 GND 0.02fF
C2422 VDD.n1863 GND 0.00fF
C2423 VDD.n1864 GND 0.00fF
C2424 VDD.t18 GND 0.35fF $ **FLOATING
C2425 VDD.n1865 GND 0.50fF
C2426 VDD.n1866 GND 0.02fF
C2427 VDD.n1867 GND 0.01fF
C2428 VDD.n1868 GND 0.00fF
C2429 VDD.n1869 GND 0.02fF
C2430 VDD.n1870 GND 0.53fF
C2431 VDD.n1871 GND 0.02fF
C2432 VDD.n1872 GND 0.01fF
C2433 VDD.n1873 GND 0.03fF
C2434 VDD.n1874 GND 0.03fF
C2435 VDD.n1875 GND 0.01fF
C2436 VDD.n1876 GND 0.02fF
C2437 VDD.n1877 GND 0.53fF
C2438 VDD.n1878 GND 0.02fF
C2439 VDD.n1879 GND 0.01fF
C2440 VDD.n1880 GND 0.02fF
C2441 VDD.t50 GND 0.35fF $ **FLOATING
C2442 VDD.n1881 GND 0.50fF
C2443 VDD.n1882 GND 0.02fF
C2444 VDD.n1883 GND 0.01fF
C2445 VDD.n1884 GND 0.02fF
C2446 VDD.n1885 GND 0.38fF
C2447 VDD.n1886 GND 0.02fF
C2448 VDD.n1887 GND 0.01fF
C2449 VDD.n1888 GND 0.02fF
C2450 VDD.t59 GND 0.35fF $ **FLOATING
C2451 VDD.n1889 GND 0.53fF
C2452 VDD.n1890 GND 0.02fF
C2453 VDD.n1891 GND 0.01fF
C2454 VDD.n1892 GND 0.02fF
C2455 VDD.n1893 GND 0.01fF
C2456 VDD.n1894 GND 0.02fF
C2457 VDD.n1895 GND 0.50fF
C2458 VDD.n1896 GND 0.01fF
C2459 VDD.n1897 GND 0.01fF
C2460 VDD.n1898 GND 0.01fF
C2461 VDD.n1903 GND 0.35fF
C2462 VDD.n1904 GND 0.02fF
C2463 VDD.n1905 GND 0.01fF
C2464 VDD.n1906 GND 0.01fF
C2465 VDD.t25 GND 0.04fF $ **FLOATING
C2466 VDD.n1907 GND 0.04fF
C2467 VDD.n1908 GND 0.02fF
C2468 VDD.t26 GND 0.35fF $ **FLOATING
C2469 VDD.n1909 GND 0.45fF
C2470 VDD.n1910 GND 0.02fF
C2471 VDD.n1911 GND 0.01fF
C2472 VDD.n1912 GND 0.03fF
C2473 VDD.n1913 GND 0.01fF
C2474 VDD.n1914 GND 0.00fF
C2475 VDD.n1915 GND 0.00fF
C2476 VDD.n1916 GND 0.01fF
C2477 VDD.n1917 GND 0.01fF
C2478 VDD.n1918 GND 0.00fF
C2479 VDD.n1919 GND 0.00fF
C2480 VDD.n1920 GND 0.00fF
C2481 VDD.n1921 GND 0.00fF
C2482 VDD.n1922 GND 0.01fF
C2483 VDD.n1923 GND 0.00fF
C2484 VDD.n1924 GND 0.01fF
C2485 VDD.n1925 GND 0.00fF
C2486 VDD.n1926 GND 0.01fF
C2487 VDD.n1927 GND 0.00fF
C2488 VDD.n1928 GND 0.01fF
C2489 VDD.n1929 GND 0.00fF
C2490 VDD.n1930 GND 0.00fF
C2491 VDD.n1931 GND 0.00fF
C2492 VDD.n1932 GND 0.00fF
C2493 VDD.n1933 GND 0.01fF
C2494 VDD.n1935 GND 0.00fF
C2495 VDD.n1936 GND 0.01fF
C2496 VDD.n1937 GND 0.00fF
C2497 VDD.n1938 GND 0.01fF
C2498 VDD.n1939 GND 0.00fF
C2499 VDD.n1940 GND 0.01fF
C2500 VDD.n1941 GND 0.00fF
C2501 VDD.n1942 GND 0.00fF
C2502 VDD.n1943 GND 0.00fF
C2503 VDD.n1944 GND 0.00fF
C2504 VDD.n1945 GND 0.01fF
C2505 VDD.n1947 GND 0.00fF
C2506 VDD.n1948 GND 0.01fF
C2507 VDD.n1949 GND 0.00fF
C2508 VDD.n1950 GND 0.01fF
C2509 VDD.n1951 GND 0.00fF
C2510 VDD.n1952 GND 0.01fF
C2511 VDD.n1953 GND 0.00fF
C2512 VDD.n1954 GND 0.00fF
C2513 VDD.n1955 GND 0.00fF
C2514 VDD.n1956 GND 0.00fF
C2515 VDD.n1957 GND 0.01fF
C2516 VDD.n1959 GND 0.00fF
C2517 VDD.n1960 GND 0.01fF
C2518 VDD.n1961 GND 0.00fF
C2519 VDD.n1962 GND 0.01fF
C2520 VDD.n1963 GND 0.00fF
C2521 VDD.n1964 GND 0.00fF
C2522 VDD.n1965 GND 0.01fF
C2523 VDD.n1966 GND 0.00fF
C2524 VDD.n1968 GND 0.01fF
C2525 VDD.n1969 GND 0.00fF
C2526 VDD.n1970 GND 0.01fF
C2527 VDD.n1971 GND 0.00fF
C2528 VDD.n1972 GND 0.00fF
C2529 VDD.n1973 GND 0.00fF
C2530 VDD.n1974 GND 0.01fF
C2531 VDD.n1975 GND 0.00fF
C2532 VDD.n1976 GND 0.00fF
C2533 VDD.n1977 GND 0.01fF
C2534 VDD.n1978 GND 0.00fF
C2535 VDD.n1980 GND 0.01fF
C2536 VDD.n1981 GND 0.00fF
C2537 VDD.n1982 GND 0.01fF
C2538 VDD.n1983 GND 0.00fF
C2539 VDD.n1984 GND 0.00fF
C2540 VDD.n1985 GND 0.00fF
C2541 VDD.n1986 GND 0.01fF
C2542 VDD.n1987 GND 0.00fF
C2543 VDD.n1988 GND 0.00fF
C2544 VDD.n1989 GND 0.01fF
C2545 VDD.n1990 GND 0.00fF
C2546 VDD.n1992 GND 0.01fF
C2547 VDD.n1993 GND 0.00fF
C2548 VDD.n1994 GND 0.01fF
C2549 VDD.n1995 GND 0.00fF
C2550 VDD.n1996 GND 0.00fF
C2551 VDD.n1997 GND 0.00fF
C2552 VDD.n1998 GND 0.01fF
C2553 VDD.n1999 GND 0.00fF
C2554 VDD.n2000 GND 0.00fF
C2555 VDD.n2001 GND 0.01fF
C2556 VDD.n2002 GND 0.00fF
C2557 VDD.n2004 GND 0.01fF
C2558 VDD.n2005 GND 0.00fF
C2559 VDD.n2006 GND 0.01fF
C2560 VDD.n2007 GND 0.00fF
C2561 VDD.n2008 GND 0.00fF
C2562 VDD.n2009 GND 0.01fF
C2563 VDD.n2010 GND 0.00fF
C2564 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/BULK GND 0.01fF
C2565 VDD.n2011 GND 0.02fF
C2566 VDD.n2012 GND 0.01fF
C2567 VDD.n2013 GND 0.02fF
C2568 VDD.n2014 GND 0.02fF
C2569 VDD.n2015 GND 0.01fF
C2570 VDD.n2016 GND 0.02fF
C2571 VDD.n2018 GND 0.02fF
C2572 VDD.n2019 GND 0.01fF
C2573 VDD.n2020 GND 0.02fF
C2574 VDD.n2021 GND 0.03fF
C2575 VDD.n2022 GND 0.01fF
C2576 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_3/BULK GND 0.01fF
C2577 VDD.n2023 GND 0.01fF
C2578 VDD.n2024 GND 0.00fF
C2579 VDD.n2025 GND 0.00fF
C2580 VDD.n2026 GND 0.00fF
C2581 VDD.n2027 GND 0.00fF
C2582 VDD.n2028 GND 0.00fF
C2583 VDD.n2029 GND 0.01fF
C2584 VDD.n2030 GND 0.00fF
C2585 VDD.n2032 GND 0.01fF
C2586 VDD.n2033 GND 0.00fF
C2587 VDD.n2034 GND 0.01fF
C2588 VDD.n2035 GND 0.00fF
C2589 VDD.n2036 GND 0.01fF
C2590 VDD.n2037 GND 0.00fF
C2591 VDD.n2038 GND 0.00fF
C2592 VDD.n2039 GND 0.00fF
C2593 VDD.n2040 GND 0.00fF
C2594 VDD.n2041 GND 0.01fF
C2595 VDD.n2042 GND 0.00fF
C2596 VDD.n2044 GND 0.01fF
C2597 VDD.n2045 GND 0.00fF
C2598 VDD.n2046 GND 0.01fF
C2599 VDD.n2047 GND 0.00fF
C2600 VDD.n2048 GND 0.01fF
C2601 VDD.n2049 GND 0.00fF
C2602 VDD.n2050 GND 0.00fF
C2603 VDD.n2051 GND 0.00fF
C2604 VDD.n2052 GND 0.00fF
C2605 VDD.n2053 GND 0.01fF
C2606 VDD.n2054 GND 0.00fF
C2607 VDD.n2056 GND 0.01fF
C2608 VDD.n2057 GND 0.00fF
C2609 VDD.n2058 GND 0.01fF
C2610 VDD.n2059 GND 0.00fF
C2611 VDD.n2060 GND 0.01fF
C2612 VDD.n2061 GND 0.00fF
C2613 VDD.n2062 GND 0.00fF
C2614 VDD.n2063 GND 0.00fF
C2615 VDD.n2064 GND 0.00fF
C2616 VDD.n2065 GND 0.01fF
C2617 VDD.n2066 GND 0.00fF
C2618 VDD.n2068 GND 0.01fF
C2619 VDD.n2069 GND 0.00fF
C2620 VDD.n2070 GND 0.01fF
C2621 VDD.n2071 GND 0.00fF
C2622 VDD.n2072 GND 0.00fF
C2623 VDD.n2073 GND 0.01fF
C2624 VDD.n2075 GND 0.00fF
C2625 VDD.n2076 GND 0.01fF
C2626 VDD.n2077 GND 0.00fF
C2627 VDD.n2078 GND 0.01fF
C2628 VDD.n2079 GND 0.00fF
C2629 VDD.n2080 GND 0.00fF
C2630 VDD.n2081 GND 0.00fF
C2631 VDD.n2082 GND 0.01fF
C2632 VDD.n2083 GND 0.00fF
C2633 VDD.n2084 GND 0.00fF
C2634 VDD.n2085 GND 0.01fF
C2635 VDD.n2087 GND 0.00fF
C2636 VDD.n2088 GND 0.01fF
C2637 VDD.n2089 GND 0.00fF
C2638 VDD.n2090 GND 0.01fF
C2639 VDD.n2091 GND 0.00fF
C2640 VDD.n2092 GND 0.00fF
C2641 VDD.n2093 GND 0.00fF
C2642 VDD.n2094 GND 0.01fF
C2643 VDD.n2095 GND 0.00fF
C2644 VDD.n2096 GND 0.00fF
C2645 VDD.n2097 GND 0.01fF
C2646 VDD.n2099 GND 0.00fF
C2647 VDD.n2100 GND 0.01fF
C2648 VDD.n2101 GND 0.00fF
C2649 VDD.n2102 GND 0.01fF
C2650 VDD.n2103 GND 0.00fF
C2651 VDD.n2104 GND 0.00fF
C2652 VDD.n2105 GND 0.00fF
C2653 VDD.n2106 GND 0.01fF
C2654 VDD.n2107 GND 0.00fF
C2655 VDD.n2108 GND 0.00fF
C2656 VDD.n2109 GND 0.01fF
C2657 VDD.n2111 GND 0.00fF
C2658 VDD.n2112 GND 0.02fF
C2659 VDD.n2113 GND 0.00fF
C2660 VDD.n2114 GND 0.01fF
C2661 VDD.n2115 GND 0.00fF
C2662 VDD.n2116 GND 0.00fF
C2663 VDD.n2117 GND 0.01fF
C2664 VDD.n2118 GND 0.01fF
C2665 VDD.n2119 GND 0.04fF
C2666 VDD.n2120 GND 0.02fF
C2667 VDD.n2121 GND 0.04fF
C2668 VDD.n2122 GND 0.01fF
C2669 VDD.n2123 GND 0.01fF
C2670 VDD.n2124 GND 0.01fF
C2671 VDD.n2125 GND 0.00fF
C2672 VDD.n2126 GND 0.00fF
C2673 VDD.n2127 GND 0.01fF
C2674 VDD.n2128 GND 0.01fF
C2675 VDD.n2129 GND 0.01fF
C2676 VDD.n2130 GND 0.00fF
C2677 VDD.n2131 GND 0.00fF
C2678 VDD.n2132 GND 0.00fF
C2679 VDD.n2133 GND 0.01fF
C2680 VDD.n2134 GND 0.00fF
C2681 VDD.n2135 GND 0.00fF
C2682 VDD.n2136 GND 0.01fF
C2683 VDD.n2137 GND 0.00fF
C2684 VDD.n2138 GND 0.00fF
C2685 VDD.n2139 GND 0.00fF
C2686 VDD.n2140 GND 0.01fF
C2687 VDD.n2141 GND 0.00fF
C2688 VDD.n2142 GND 0.00fF
C2689 VDD.n2143 GND 0.01fF
C2690 VDD.n2144 GND 0.00fF
C2691 VDD.n2145 GND 0.00fF
C2692 VDD.n2146 GND 0.00fF
C2693 VDD.n2147 GND 0.01fF
C2694 VDD.n2148 GND 0.00fF
C2695 VDD.n2149 GND 0.00fF
C2696 VDD.n2150 GND 0.01fF
C2697 VDD.n2151 GND 0.00fF
C2698 VDD.n2152 GND 0.00fF
C2699 VDD.n2153 GND 0.00fF
C2700 VDD.n2154 GND 0.01fF
C2701 VDD.n2155 GND 0.00fF
C2702 VDD.n2156 GND 0.00fF
C2703 VDD.n2157 GND 0.01fF
C2704 VDD.n2158 GND 0.00fF
C2705 VDD.n2159 GND 0.00fF
C2706 VDD.n2160 GND 0.00fF
C2707 VDD.n2161 GND 0.00fF
C2708 VDD.n2162 GND 0.00fF
C2709 VDD.n2163 GND 0.00fF
C2710 VDD.n2164 GND 0.00fF
C2711 VDD.n2165 GND 0.00fF
C2712 VDD.n2166 GND 0.00fF
C2713 VDD.n2167 GND 0.00fF
C2714 VDD.n2168 GND 0.00fF
C2715 VDD.n2169 GND 0.00fF
C2716 VDD.n2170 GND 0.00fF
C2717 VDD.n2171 GND 0.00fF
C2718 VDD.n2172 GND 0.00fF
C2719 VDD.n2173 GND 0.00fF
C2720 VDD.n2174 GND 0.00fF
C2721 VDD.n2175 GND 0.00fF
C2722 VDD.n2176 GND 0.00fF
C2723 VDD.n2177 GND 0.00fF
C2724 VDD.n2178 GND 0.00fF
C2725 VDD.n2179 GND 0.00fF
C2726 VDD.n2180 GND 0.00fF
C2727 VDD.n2181 GND 0.00fF
C2728 VDD.n2182 GND 0.00fF
C2729 VDD.n2183 GND 0.00fF
C2730 VDD.n2184 GND 0.00fF
C2731 VDD.n2185 GND 0.00fF
C2732 VDD.n2186 GND 0.00fF
C2733 VDD.n2187 GND 0.00fF
C2734 VDD.n2188 GND 0.00fF
C2735 VDD.n2189 GND 0.00fF
C2736 VDD.n2190 GND 0.00fF
C2737 VDD.n2191 GND 0.00fF
C2738 VDD.n2192 GND 0.11fF
C2739 VDD.n2193 GND 0.01fF
C2740 VDD.n2194 GND 0.00fF
C2741 VDD.n2195 GND 0.01fF
C2742 VDD.n2196 GND 0.03fF
C2743 VDD.n2197 GND 0.58fF
C2744 VDD.n2198 GND 0.02fF
C2745 VDD.n2199 GND 0.01fF
C2746 VDD.n2200 GND 0.04fF
C2747 VDD.n2201 GND 0.03fF
C2748 VDD.n2202 GND 0.02fF
C2749 VDD.n2203 GND 0.47fF
C2750 VDD.n2204 GND 0.01fF
C2751 VDD.n2205 GND 0.01fF
C2752 VDD.n2206 GND 0.01fF
C2753 VDD.n2207 GND 0.02fF
C2754 VDD.n2208 GND 0.55fF
C2755 VDD.n2209 GND 0.02fF
C2756 VDD.n2210 GND 0.01fF
C2757 VDD.n2211 GND 0.02fF
C2758 VDD.t43 GND 0.35fF $ **FLOATING
C2759 VDD.n2212 GND 0.38fF
C2760 VDD.n2213 GND 0.02fF
C2761 VDD.n2214 GND 0.01fF
C2762 VDD.n2215 GND 0.02fF
C2763 VDD.t53 GND 0.35fF $ **FLOATING
C2764 VDD.n2216 GND 0.47fF
C2765 VDD.n2217 GND 0.02fF
C2766 VDD.n2218 GND 0.01fF
C2767 VDD.n2219 GND 0.02fF
C2768 VDD.n2220 GND 0.55fF
C2769 VDD.n2221 GND 0.02fF
C2770 VDD.n2222 GND 0.01fF
C2771 VDD.n2223 GND 0.02fF
C2772 VDD.n2224 GND 0.02fF
C2773 VDD.n2225 GND 0.02fF
C2774 VDD.n2226 GND 0.01fF
C2775 VDD.n2227 GND 0.00fF
C2776 VDD.n2228 GND 0.00fF
C2777 VDD.n2229 GND 0.00fF
C2778 VDD.n2230 GND 0.00fF
C2779 VDD.n2231 GND 0.01fF
C2780 VDD.n2232 GND 0.00fF
C2781 VDD.n2233 GND 0.00fF
C2782 VDD.n2234 GND 0.01fF
C2783 VDD.n2235 GND 0.01fF
C2784 VDD.n2236 GND 0.00fF
C2785 VDD.n2237 GND 0.01fF
C2786 VDD.n2238 GND 0.01fF
C2787 VDD.n2239 GND 0.00fF
C2788 VDD.n2240 GND 0.01fF
C2789 VDD.n2241 GND 0.01fF
C2790 VDD.n2242 GND 0.00fF
C2791 VDD.n2243 GND 0.01fF
C2792 VDD.n2244 GND 0.01fF
C2793 VDD.n2245 GND 0.00fF
C2794 VDD.n2246 GND 0.01fF
C2795 VDD.n2247 GND 0.01fF
C2796 VDD.n2248 GND 0.00fF
C2797 VDD.n2249 GND 0.01fF
C2798 VDD.n2250 GND 0.01fF
C2799 VDD.n2251 GND 0.00fF
C2800 VDD.n2252 GND 0.01fF
C2801 VDD.n2253 GND 0.01fF
C2802 VDD.n2254 GND 0.00fF
C2803 VDD.n2255 GND 0.01fF
C2804 VDD.n2256 GND 0.02fF
C2805 VDD.n2257 GND 0.02fF
C2806 VDD.n2258 GND 0.02fF
C2807 VDD.n2259 GND 0.02fF
C2808 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/BULK GND 0.01fF
C2809 VDD.n2260 GND 0.01fF
C2810 VDD.n2261 GND 0.00fF
C2811 VDD.n2262 GND 0.00fF
C2812 VDD.n2263 GND 0.00fF
C2813 VDD.n2264 GND 0.00fF
C2814 VDD.n2265 GND 0.00fF
C2815 VDD.n2266 GND 0.01fF
C2816 VDD.n2267 GND 0.00fF
C2817 VDD.n2269 GND 0.01fF
C2818 VDD.n2270 GND 0.00fF
C2819 VDD.n2271 GND 0.01fF
C2820 VDD.n2272 GND 0.00fF
C2821 VDD.n2273 GND 0.01fF
C2822 VDD.n2274 GND 0.00fF
C2823 VDD.n2275 GND 0.00fF
C2824 VDD.n2276 GND 0.00fF
C2825 VDD.n2277 GND 0.00fF
C2826 VDD.n2278 GND 0.01fF
C2827 VDD.n2279 GND 0.00fF
C2828 VDD.n2281 GND 0.01fF
C2829 VDD.n2282 GND 0.00fF
C2830 VDD.n2283 GND 0.01fF
C2831 VDD.n2284 GND 0.00fF
C2832 VDD.n2285 GND 0.01fF
C2833 VDD.n2286 GND 0.00fF
C2834 VDD.n2287 GND 0.00fF
C2835 VDD.n2288 GND 0.00fF
C2836 VDD.n2289 GND 0.00fF
C2837 VDD.n2290 GND 0.01fF
C2838 VDD.n2291 GND 0.00fF
C2839 VDD.n2293 GND 0.01fF
C2840 VDD.n2294 GND 0.00fF
C2841 VDD.n2295 GND 0.01fF
C2842 VDD.n2296 GND 0.00fF
C2843 VDD.n2297 GND 0.01fF
C2844 VDD.n2298 GND 0.00fF
C2845 VDD.n2299 GND 0.00fF
C2846 VDD.n2300 GND 0.00fF
C2847 VDD.n2301 GND 0.00fF
C2848 VDD.n2302 GND 0.01fF
C2849 VDD.n2303 GND 0.00fF
C2850 VDD.n2305 GND 0.01fF
C2851 VDD.n2306 GND 0.00fF
C2852 VDD.n2307 GND 0.01fF
C2853 VDD.n2308 GND 0.00fF
C2854 VDD.n2309 GND 0.00fF
C2855 VDD.n2310 GND 0.01fF
C2856 VDD.n2312 GND 0.00fF
C2857 VDD.n2313 GND 0.01fF
C2858 VDD.n2314 GND 0.00fF
C2859 VDD.n2315 GND 0.01fF
C2860 VDD.n2316 GND 0.00fF
C2861 VDD.n2317 GND 0.00fF
C2862 VDD.n2318 GND 0.00fF
C2863 VDD.n2319 GND 0.01fF
C2864 VDD.n2320 GND 0.00fF
C2865 VDD.n2321 GND 0.00fF
C2866 VDD.n2322 GND 0.01fF
C2867 VDD.n2324 GND 0.00fF
C2868 VDD.n2325 GND 0.01fF
C2869 VDD.n2326 GND 0.00fF
C2870 VDD.n2327 GND 0.01fF
C2871 VDD.n2328 GND 0.00fF
C2872 VDD.n2329 GND 0.00fF
C2873 VDD.n2330 GND 0.00fF
C2874 VDD.n2331 GND 0.01fF
C2875 VDD.n2332 GND 0.00fF
C2876 VDD.n2333 GND 0.00fF
C2877 VDD.n2334 GND 0.01fF
C2878 VDD.n2336 GND 0.00fF
C2879 VDD.n2337 GND 0.01fF
C2880 VDD.n2338 GND 0.00fF
C2881 VDD.n2339 GND 0.01fF
C2882 VDD.n2340 GND 0.00fF
C2883 VDD.n2341 GND 0.00fF
C2884 VDD.n2342 GND 0.00fF
C2885 VDD.n2343 GND 0.01fF
C2886 VDD.n2344 GND 0.00fF
C2887 VDD.n2345 GND 0.00fF
C2888 VDD.n2346 GND 0.01fF
C2889 VDD.n2347 GND 0.00fF
C2890 VDD.n2348 GND 0.01fF
C2891 VDD.n2349 GND 0.00fF
C2892 VDD.n2350 GND 0.01fF
C2893 VDD.n2351 GND 0.00fF
C2894 VDD.n2352 GND 0.00fF
C2895 VDD.n2353 GND 0.01fF
C2896 VDD.n2354 GND 0.01fF
C2897 VDD.n2355 GND 0.02fF
C2898 VDD.n2356 GND 0.01fF
C2899 VDD.n2357 GND 0.02fF
C2900 VDD.n2358 GND 0.02fF
C2901 VDD.n2359 GND 0.02fF
C2902 VDD.n2360 GND 0.01fF
C2903 VDD.n2361 GND 0.02fF
C2904 VDD.n2362 GND 0.02fF
C2905 VDD.n2363 GND 0.01fF
C2906 VDD.n2364 GND 0.02fF
C2907 VDD.n2365 GND 0.02fF
C2908 VDD.n2366 GND 0.01fF
C2909 VDD.n2367 GND 0.02fF
C2910 VDD.n2368 GND 0.02fF
C2911 VDD.n2369 GND 0.01fF
C2912 VDD.n2370 GND 0.02fF
C2913 VDD.n2371 GND 0.01fF
C2914 VDD.n2372 GND 0.02fF
C2915 VDD.n2373 GND 0.01fF
C2916 VDD.n2374 GND 0.01fF
C2917 VDD.n2375 GND 0.01fF
C2918 VDD.n2376 GND 0.02fF
C2919 VDD.n2377 GND 0.02fF
C2920 VDD.n2378 GND 0.01fF
C2921 VDD.n2379 GND 0.02fF
C2922 VDD.n2380 GND 0.02fF
C2923 VDD.n2381 GND 0.01fF
C2924 VDD.n2382 GND 0.02fF
C2925 VDD.n2383 GND 0.02fF
C2926 VDD.n2384 GND 0.01fF
C2927 VDD.n2385 GND 0.02fF
C2928 VDD.n2386 GND 0.02fF
C2929 VDD.n2387 GND 0.01fF
C2930 VDD.n2388 GND 0.02fF
C2931 VDD.n2389 GND 0.01fF
C2932 VDD.n2390 GND 0.02fF
C2933 VDD.n2391 GND 0.01fF
C2934 VDD.n2392 GND 0.01fF
C2935 VDD.n2393 GND 0.01fF
C2936 VDD.n2394 GND 0.02fF
C2937 VDD.n2395 GND 0.02fF
C2938 VDD.n2396 GND 0.01fF
C2939 VDD.n2397 GND 0.02fF
C2940 VDD.n2398 GND 0.02fF
C2941 VDD.n2399 GND 0.01fF
C2942 VDD.n2400 GND 0.02fF
C2943 VDD.n2401 GND 0.02fF
C2944 VDD.n2402 GND 0.01fF
C2945 VDD.n2403 GND 0.02fF
C2946 VDD.n2404 GND 0.02fF
C2947 VDD.n2405 GND 0.01fF
C2948 VDD.n2406 GND 0.02fF
C2949 VDD.n2407 GND 0.01fF
C2950 VDD.n2408 GND 0.02fF
C2951 VDD.n2409 GND 0.01fF
C2952 VDD.n2410 GND 0.01fF
C2953 VDD.n2411 GND 0.01fF
C2954 VDD.n2412 GND 0.02fF
C2955 VDD.n2413 GND 0.01fF
C2956 VDD.n2414 GND 0.01fF
C2957 VDD.n2415 GND 0.01fF
C2958 VDD.n2416 GND 0.01fF
C2959 VDD.t5 GND 0.04fF $ **FLOATING
C2960 VDD.n2417 GND 0.04fF
C2961 VDD.n2418 GND 0.02fF
C2962 VDD.n2419 GND 0.02fF
C2963 VDD.n2420 GND 0.02fF
C2964 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/GATE GND 0.02fF
C2965 VDD.n2421 GND 0.01fF
C2966 VDD.n2422 GND 0.00fF
C2967 VDD.n2423 GND 0.00fF
C2968 VDD.n2424 GND 0.00fF
C2969 VDD.n2425 GND 0.01fF
C2970 VDD.n2426 GND 0.01fF
C2971 VDD.n2427 GND 0.00fF
C2972 VDD.n2428 GND 0.00fF
C2973 VDD.n2429 GND 0.00fF
C2974 VDD.n2430 GND 0.01fF
C2975 VDD.n2431 GND 0.00fF
C2976 VDD.n2432 GND 0.00fF
C2977 VDD.n2433 GND 0.01fF
C2978 VDD.n2434 GND 0.00fF
C2979 VDD.n2435 GND 0.00fF
C2980 VDD.n2436 GND 0.00fF
C2981 VDD.n2437 GND 0.01fF
C2982 VDD.n2438 GND 0.00fF
C2983 VDD.n2439 GND 0.00fF
C2984 VDD.n2440 GND 0.01fF
C2985 VDD.n2441 GND 0.00fF
C2986 VDD.n2442 GND 0.00fF
C2987 VDD.n2443 GND 0.00fF
C2988 VDD.n2444 GND 0.01fF
C2989 VDD.n2445 GND 0.00fF
C2990 VDD.n2446 GND 0.00fF
C2991 VDD.n2447 GND 0.01fF
C2992 VDD.n2448 GND 0.00fF
C2993 VDD.n2449 GND 0.00fF
C2994 VDD.n2450 GND 0.00fF
C2995 VDD.n2451 GND 0.01fF
C2996 VDD.n2452 GND 0.00fF
C2997 VDD.n2453 GND 0.00fF
C2998 VDD.n2454 GND 0.01fF
C2999 VDD.n2455 GND 0.00fF
C3000 VDD.n2456 GND 0.00fF
C3001 VDD.n2457 GND 0.00fF
C3002 VDD.n2458 GND 0.00fF
C3003 VDD.n2459 GND 0.00fF
C3004 VDD.n2460 GND 0.00fF
C3005 VDD.n2461 GND 0.00fF
C3006 VDD.n2462 GND 0.00fF
C3007 VDD.n2463 GND 0.00fF
C3008 VDD.n2464 GND 0.00fF
C3009 VDD.n2465 GND 0.00fF
C3010 VDD.n2466 GND 0.00fF
C3011 VDD.n2467 GND 0.00fF
C3012 VDD.n2468 GND 0.00fF
C3013 VDD.n2469 GND 0.00fF
C3014 VDD.n2470 GND 0.00fF
C3015 VDD.n2471 GND 0.00fF
C3016 VDD.n2472 GND 0.00fF
C3017 VDD.n2473 GND 0.00fF
C3018 VDD.n2474 GND 0.00fF
C3019 VDD.n2475 GND 0.00fF
C3020 VDD.n2476 GND 0.00fF
C3021 VDD.n2477 GND 0.00fF
C3022 VDD.n2478 GND 0.00fF
C3023 VDD.n2479 GND 0.00fF
C3024 VDD.n2480 GND 0.00fF
C3025 VDD.n2481 GND 0.00fF
C3026 VDD.n2482 GND 0.00fF
C3027 VDD.n2483 GND 0.00fF
C3028 VDD.n2484 GND 0.00fF
C3029 VDD.n2485 GND 0.00fF
C3030 VDD.n2486 GND 0.00fF
C3031 VDD.n2487 GND 0.00fF
C3032 VDD.t8 GND 0.04fF $ **FLOATING
C3033 VDD.n2488 GND 0.11fF
C3034 VDD.n2489 GND 0.01fF
C3035 VDD.n2490 GND 0.00fF
C3036 VDD.n2491 GND 0.01fF
C3037 VDD.n2492 GND 0.00fF
C3038 VDD.n2493 GND 0.00fF
C3039 VDD.n2494 GND 0.00fF
C3040 VDD.n2495 GND 0.01fF
C3041 VDD.n2496 GND 0.01fF
C3042 VDD.n2497 GND 0.00fF
C3043 VDD.n2498 GND 0.00fF
C3044 VDD.n2499 GND 0.00fF
C3045 VDD.n2500 GND 0.00fF
C3046 VDD.n2501 GND 0.00fF
C3047 VDD.n2502 GND 0.00fF
C3048 VDD.n2503 GND 0.00fF
C3049 VDD.n2504 GND 0.00fF
C3050 VDD.n2505 GND 0.00fF
C3051 VDD.n2506 GND 0.00fF
C3052 VDD.n2507 GND 0.00fF
C3053 VDD.n2508 GND 0.00fF
C3054 VDD.n2509 GND 0.00fF
C3055 VDD.n2510 GND 0.00fF
C3056 VDD.n2511 GND 0.00fF
C3057 VDD.n2512 GND 0.00fF
C3058 VDD.n2513 GND 0.00fF
C3059 VDD.n2514 GND 0.00fF
C3060 VDD.n2515 GND 0.00fF
C3061 VDD.n2516 GND 0.00fF
C3062 VDD.n2517 GND 0.00fF
C3063 VDD.n2518 GND 0.00fF
C3064 VDD.n2519 GND 0.00fF
C3065 VDD.n2520 GND 0.00fF
C3066 VDD.n2521 GND 0.00fF
C3067 VDD.n2522 GND 0.00fF
C3068 VDD.n2523 GND 0.00fF
C3069 VDD.n2524 GND 0.00fF
C3070 VDD.n2525 GND 0.00fF
C3071 VDD.n2526 GND 0.00fF
C3072 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/DRAIN GND 0.00fF
C3073 VDD.n2527 GND 0.01fF
C3074 VDD.n2528 GND 0.01fF
C3075 VDD.n2529 GND 0.01fF
C3076 VDD.n2530 GND 0.02fF
C3077 VDD.n2531 GND 0.02fF
C3078 VDD.n2532 GND 0.01fF
C3079 VDD.n2533 GND 0.01fF
C3080 VDD.n2534 GND 0.02fF
C3081 VDD.n2535 GND 0.02fF
C3082 VDD.n2536 GND 0.01fF
C3083 VDD.n2537 GND 0.03fF
C3084 VDD.n2538 GND 0.03fF
C3085 VDD.n2539 GND 0.04fF
C3086 VDD.n2540 GND 0.00fF
C3087 VDD.n2541 GND 0.00fF
C3088 VDD.n2542 GND 0.00fF
C3089 VDD.n2543 GND 0.00fF
C3090 VDD.n2544 GND 0.00fF
C3091 VDD.n2545 GND 0.00fF
C3092 VDD.n2546 GND 0.01fF
C3093 VDD.n2547 GND 0.00fF
C3094 VDD.n2548 GND 0.01fF
C3095 VDD.n2549 GND 0.00fF
C3096 VDD.n2550 GND 0.00fF
C3097 VDD.n2551 GND 0.00fF
C3098 VDD.n2552 GND 0.00fF
C3099 VDD.n2553 GND 0.01fF
C3100 VDD.n2554 GND 0.00fF
C3101 VDD.n2555 GND 0.01fF
C3102 VDD.n2556 GND 0.00fF
C3103 VDD.n2557 GND 0.00fF
C3104 VDD.n2558 GND 0.00fF
C3105 VDD.n2559 GND 0.00fF
C3106 VDD.n2560 GND 0.01fF
C3107 VDD.n2561 GND 0.00fF
C3108 VDD.n2562 GND 0.01fF
C3109 VDD.n2563 GND 0.00fF
C3110 VDD.n2564 GND 0.00fF
C3111 VDD.n2565 GND 0.00fF
C3112 VDD.n2566 GND 0.00fF
C3113 VDD.n2567 GND 0.01fF
C3114 VDD.n2568 GND 0.00fF
C3115 VDD.n2569 GND 0.01fF
C3116 VDD.n2570 GND 0.00fF
C3117 VDD.n2571 GND 0.00fF
C3118 VDD.t7 GND 0.04fF $ **FLOATING
C3119 VDD.n2572 GND 0.07fF
C3120 VDD.n2573 GND 0.01fF
C3121 VDD.n2574 GND 0.01fF
C3122 VDD.n2575 GND 0.00fF
C3123 VDD.n2576 GND 0.00fF
C3124 VDD.n2577 GND 0.00fF
C3125 VDD.n2578 GND 0.00fF
C3126 VDD.n2579 GND 0.00fF
C3127 VDD.n2580 GND 0.00fF
C3128 VDD.n2581 GND 0.00fF
C3129 VDD.n2582 GND 0.01fF
C3130 VDD.n2583 GND 0.00fF
C3131 VDD.n2584 GND 0.00fF
C3132 VDD.n2585 GND 0.01fF
C3133 VDD.n2586 GND 0.00fF
C3134 VDD.n2587 GND 0.00fF
C3135 VDD.n2588 GND 0.00fF
C3136 VDD.n2589 GND 0.01fF
C3137 VDD.n2590 GND 0.00fF
C3138 VDD.n2591 GND 0.00fF
C3139 VDD.n2592 GND 0.01fF
C3140 VDD.n2593 GND 0.00fF
C3141 VDD.n2594 GND 0.00fF
C3142 VDD.n2595 GND 0.00fF
C3143 VDD.n2596 GND 0.01fF
C3144 VDD.n2597 GND 0.00fF
C3145 VDD.n2598 GND 0.00fF
C3146 VDD.n2599 GND 0.01fF
C3147 VDD.n2600 GND 0.00fF
C3148 VDD.n2601 GND 0.00fF
C3149 VDD.n2602 GND 0.00fF
C3150 VDD.n2603 GND 0.01fF
C3151 VDD.n2604 GND 0.00fF
C3152 VDD.n2605 GND 0.00fF
C3153 VDD.n2606 GND 0.01fF
C3154 VDD.n2607 GND 0.00fF
C3155 VDD.n2608 GND 0.00fF
C3156 VDD.n2609 GND 0.00fF
C3157 VDD.n2610 GND 0.00fF
C3158 VDD.n2611 GND 0.00fF
C3159 VDD.n2612 GND 0.00fF
C3160 VDD.n2613 GND 0.00fF
C3161 VDD.n2614 GND 0.00fF
C3162 VDD.n2615 GND 0.00fF
C3163 VDD.n2616 GND 0.00fF
C3164 VDD.n2617 GND 0.00fF
C3165 VDD.n2618 GND 0.00fF
C3166 VDD.n2619 GND 0.00fF
C3167 VDD.n2620 GND 0.00fF
C3168 VDD.n2621 GND 0.00fF
C3169 VDD.n2622 GND 0.00fF
C3170 VDD.n2623 GND 0.00fF
C3171 VDD.n2624 GND 0.00fF
C3172 VDD.n2625 GND 0.00fF
C3173 VDD.n2626 GND 0.00fF
C3174 VDD.n2627 GND 0.00fF
C3175 VDD.n2628 GND 0.00fF
C3176 VDD.n2629 GND 0.00fF
C3177 VDD.n2630 GND 0.00fF
C3178 VDD.n2631 GND 0.00fF
C3179 VDD.n2632 GND 0.00fF
C3180 VDD.n2633 GND 0.00fF
C3181 VDD.n2634 GND 0.00fF
C3182 VDD.n2635 GND 0.00fF
C3183 VDD.n2636 GND 0.00fF
C3184 VDD.n2637 GND 0.00fF
C3185 VDD.n2638 GND 0.02fF
C3186 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/SOURCE GND 0.01fF
C3187 VDD.n2639 GND 0.02fF
C3188 VDD.n2640 GND 0.01fF
C3189 VDD.n2641 GND 0.03fF
C3190 VDD.n2642 GND 0.03fF
C3191 VDD.n2643 GND 0.01fF
C3192 VDD.n2644 GND 0.02fF
C3193 VDD.n2645 GND 0.02fF
C3194 VDD.n2646 GND 0.01fF
C3195 VDD.n2647 GND 0.01fF
C3196 VDD.n2648 GND 0.02fF
C3197 VDD.n2649 GND 0.02fF
C3198 VDD.n2650 GND 0.01fF
C3199 VDD.n2651 GND 0.01fF
C3200 VDD.n2652 GND 0.00fF
C3201 VDD.n2653 GND 0.07fF
C3202 VDD.n2654 GND 0.11fF
C3203 VDD.n2655 GND 0.01fF
C3204 VDD.n2656 GND 0.00fF
C3205 VDD.n2657 GND 0.01fF
C3206 VDD.n2658 GND 0.03fF
C3207 VDD.n2659 GND 0.01fF
C3208 VDD.n2660 GND 0.02fF
C3209 VDD.t46 GND 0.35fF $ **FLOATING
C3210 VDD.n2661 GND 0.39fF
C3211 VDD.n2662 GND 0.02fF
C3212 VDD.n2663 GND 0.01fF
C3213 VDD.n2664 GND 0.02fF
C3214 VDD.t55 GND 0.35fF $ **FLOATING
C3215 VDD.n2665 GND 0.38fF
C3216 VDD.n2666 GND 0.02fF
C3217 VDD.n2667 GND 0.01fF
C3218 VDD.n2668 GND 0.02fF
C3219 VDD.n2669 GND 0.63fF
C3220 VDD.n2670 GND 0.02fF
C3221 VDD.n2671 GND 0.01fF
C3222 VDD.n2672 GND 0.02fF
C3223 VDD.n2673 GND 0.01fF
C3224 VDD.n2674 GND 0.02fF
C3225 VDD.n2675 GND 0.39fF
C3226 VDD.n2676 GND 0.01fF
C3227 VDD.n2677 GND 0.01fF
C3228 VDD.n2678 GND 0.02fF
C3229 VDD.n2679 GND 0.00fF
C3230 VDD.n2680 GND 0.00fF
C3231 VDD.n2681 GND 0.04fF
C3232 VDD.n2682 GND 0.01fF
C3233 VDD.n2683 GND 0.01fF
C3234 VDD.n2684 GND 0.01fF
C3235 VDD.n2685 GND 0.00fF
C3236 VDD.n2686 GND 0.00fF
C3237 VDD.n2687 GND 0.01fF
C3238 VDD.n2688 GND 0.01fF
C3239 VDD.n2689 GND 0.01fF
C3240 VDD.n2690 GND 0.00fF
C3241 VDD.n2691 GND 0.00fF
C3242 VDD.n2692 GND 0.00fF
C3243 VDD.n2693 GND 0.01fF
C3244 VDD.n2694 GND 0.00fF
C3245 VDD.n2695 GND 0.00fF
C3246 VDD.n2696 GND 0.01fF
C3247 VDD.n2697 GND 0.00fF
C3248 VDD.n2698 GND 0.00fF
C3249 VDD.n2699 GND 0.00fF
C3250 VDD.n2700 GND 0.01fF
C3251 VDD.n2701 GND 0.00fF
C3252 VDD.n2702 GND 0.00fF
C3253 VDD.n2703 GND 0.01fF
C3254 VDD.n2704 GND 0.00fF
C3255 VDD.n2705 GND 0.00fF
C3256 VDD.n2706 GND 0.00fF
C3257 VDD.n2707 GND 0.01fF
C3258 VDD.n2708 GND 0.00fF
C3259 VDD.n2709 GND 0.00fF
C3260 VDD.n2710 GND 0.01fF
C3261 VDD.n2711 GND 0.00fF
C3262 VDD.n2712 GND 0.00fF
C3263 VDD.n2713 GND 0.00fF
C3264 VDD.n2714 GND 0.01fF
C3265 VDD.n2715 GND 0.00fF
C3266 VDD.n2716 GND 0.00fF
C3267 VDD.n2717 GND 0.01fF
C3268 VDD.n2718 GND 0.00fF
C3269 VDD.n2719 GND 0.00fF
C3270 VDD.n2720 GND 0.00fF
C3271 VDD.n2721 GND 0.00fF
C3272 VDD.n2722 GND 0.00fF
C3273 VDD.n2723 GND 0.00fF
C3274 VDD.n2724 GND 0.00fF
C3275 VDD.n2725 GND 0.00fF
C3276 VDD.n2726 GND 0.00fF
C3277 VDD.n2727 GND 0.00fF
C3278 VDD.n2728 GND 0.00fF
C3279 VDD.n2729 GND 0.00fF
C3280 VDD.n2730 GND 0.00fF
C3281 VDD.n2731 GND 0.00fF
C3282 VDD.n2732 GND 0.00fF
C3283 VDD.n2733 GND 0.00fF
C3284 VDD.n2734 GND 0.00fF
C3285 VDD.n2735 GND 0.00fF
C3286 VDD.n2736 GND 0.00fF
C3287 VDD.n2737 GND 0.00fF
C3288 VDD.n2738 GND 0.00fF
C3289 VDD.n2739 GND 0.00fF
C3290 VDD.n2740 GND 0.00fF
C3291 VDD.n2741 GND 0.00fF
C3292 VDD.n2742 GND 0.00fF
C3293 VDD.n2743 GND 0.00fF
C3294 VDD.n2744 GND 0.00fF
C3295 VDD.n2745 GND 0.00fF
C3296 VDD.n2746 GND 0.00fF
C3297 VDD.n2747 GND 0.00fF
C3298 VDD.n2748 GND 0.00fF
C3299 VDD.n2749 GND 0.00fF
C3300 VDD.n2750 GND 0.00fF
C3301 VDD.n2751 GND 0.00fF
C3302 VDD.n2752 GND 0.11fF
C3303 VDD.n2753 GND 0.01fF
C3304 VDD.n2754 GND 0.00fF
C3305 VDD.n2755 GND 0.01fF
C3306 VDD.n2756 GND 0.00fF
C3307 VDD.n2757 GND 0.00fF
C3308 VDD.n2758 GND 0.00fF
C3309 VDD.n2759 GND 0.01fF
C3310 VDD.n2760 GND 0.01fF
C3311 VDD.n2761 GND 0.03fF
C3312 VDD.n2762 GND 0.01fF
C3313 VDD.n2763 GND 0.01fF
C3314 VDD.n2764 GND 0.00fF
C3315 VDD.n2765 GND 0.00fF
C3316 VDD.n2766 GND 0.00fF
C3317 VDD.n2767 GND 0.00fF
C3318 VDD.n2768 GND 0.00fF
C3319 VDD.n2769 GND 0.00fF
C3320 VDD.n2770 GND 0.00fF
C3321 VDD.n2771 GND 0.00fF
C3322 VDD.n2772 GND 0.00fF
C3323 VDD.n2773 GND 0.00fF
C3324 VDD.n2774 GND 0.00fF
C3325 VDD.n2775 GND 0.00fF
C3326 VDD.n2776 GND 0.00fF
C3327 VDD.n2777 GND 0.00fF
C3328 VDD.n2778 GND 0.00fF
C3329 VDD.n2779 GND 0.00fF
C3330 VDD.n2780 GND 0.00fF
C3331 VDD.n2781 GND 0.00fF
C3332 VDD.n2782 GND 0.00fF
C3333 VDD.n2783 GND 0.00fF
C3334 VDD.n2784 GND 0.00fF
C3335 VDD.n2785 GND 0.00fF
C3336 VDD.n2786 GND 0.00fF
C3337 VDD.n2787 GND 0.00fF
C3338 VDD.n2788 GND 0.00fF
C3339 VDD.n2789 GND 0.00fF
C3340 VDD.n2790 GND 0.00fF
C3341 VDD.n2791 GND 0.00fF
C3342 VDD.n2792 GND 0.00fF
C3343 VDD.n2793 GND 0.00fF
C3344 VDD.n2794 GND 0.00fF
C3345 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/DRAIN GND 0.00fF
C3346 VDD.n2795 GND 0.01fF
C3347 VDD.n2796 GND 0.01fF
C3348 VDD.n2797 GND 0.01fF
C3349 VDD.n2798 GND 0.02fF
C3350 VDD.n2799 GND 0.02fF
C3351 VDD.n2800 GND 0.01fF
C3352 VDD.n2801 GND 0.01fF
C3353 VDD.n2802 GND 0.02fF
C3354 VDD.n2803 GND 0.02fF
C3355 VDD.n2804 GND 0.01fF
C3356 VDD.n2805 GND 0.03fF
C3357 VDD.n2806 GND 0.03fF
C3358 VDD.n2807 GND 0.04fF
C3359 VDD.n2808 GND 0.00fF
C3360 VDD.n2809 GND 0.00fF
C3361 VDD.n2810 GND 0.00fF
C3362 VDD.n2811 GND 0.00fF
C3363 VDD.n2812 GND 0.00fF
C3364 VDD.n2813 GND 0.01fF
C3365 VDD.n2814 GND 0.00fF
C3366 VDD.n2815 GND 0.01fF
C3367 VDD.n2816 GND 0.00fF
C3368 VDD.n2817 GND 0.00fF
C3369 VDD.n2818 GND 0.00fF
C3370 VDD.n2819 GND 0.00fF
C3371 VDD.n2820 GND 0.01fF
C3372 VDD.n2821 GND 0.00fF
C3373 VDD.n2822 GND 0.01fF
C3374 VDD.n2823 GND 0.00fF
C3375 VDD.n2824 GND 0.00fF
C3376 VDD.n2825 GND 0.00fF
C3377 VDD.n2826 GND 0.00fF
C3378 VDD.n2827 GND 0.01fF
C3379 VDD.n2828 GND 0.00fF
C3380 VDD.n2829 GND 0.01fF
C3381 VDD.n2830 GND 0.00fF
C3382 VDD.n2831 GND 0.00fF
C3383 VDD.n2832 GND 0.00fF
C3384 VDD.n2833 GND 0.00fF
C3385 VDD.n2834 GND 0.01fF
C3386 VDD.n2835 GND 0.00fF
C3387 VDD.n2836 GND 0.01fF
C3388 VDD.n2837 GND 0.00fF
C3389 VDD.n2838 GND 0.00fF
C3390 VDD.n2839 GND 0.07fF
C3391 VDD.t10 GND 0.04fF $ **FLOATING
C3392 VDD.n2840 GND 0.07fF
C3393 VDD.n2841 GND 0.01fF
C3394 VDD.n2842 GND 0.01fF
C3395 VDD.n2843 GND 0.01fF
C3396 VDD.n2844 GND 0.00fF
C3397 VDD.n2845 GND 0.01fF
C3398 VDD.n2846 GND 0.01fF
C3399 VDD.n2847 GND 0.02fF
C3400 VDD.n2848 GND 0.02fF
C3401 VDD.n2849 GND 0.02fF
C3402 VDD.n2850 GND 0.02fF
C3403 VDD.t6 GND 0.35fF $ **FLOATING
C3404 VDD.n2851 GND 0.38fF
C3405 VDD.n2852 GND 0.02fF
C3406 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/GATE GND 0.02fF
C3407 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_6/BULK GND 0.02fF
C3408 VDD.n2853 GND 0.00fF
C3409 VDD.n2854 GND 0.00fF
C3410 VDD.n2855 GND 0.00fF
C3411 VDD.n2856 GND 0.00fF
C3412 VDD.n2857 GND 0.02fF
C3413 VDD.t9 GND 0.04fF $ **FLOATING
C3414 VDD.n2858 GND 0.04fF
C3415 VDD.n2859 GND 0.02fF
C3416 VDD.n2860 GND 0.01fF
C3417 VDD.n2861 GND 0.02fF
C3418 VDD.n2862 GND 0.01fF
C3419 VDD.t11 GND 0.04fF $ **FLOATING
C3420 VDD.n2863 GND 0.11fF
C3421 VDD.n2864 GND 0.01fF
C3422 VDD.n2865 GND 0.00fF
C3423 VDD.n2866 GND 0.02fF
C3424 VDD.n2867 GND 0.02fF
C3425 VDD.n2868 GND 0.01fF
C3426 VDD.n2869 GND 0.03fF
C3427 VDD.n2870 GND 0.03fF
C3428 VDD.n2871 GND 0.01fF
C3429 VDD.n2872 GND 0.02fF
C3430 VDD.n2873 GND 0.02fF
C3431 VDD.n2874 GND 0.01fF
C3432 VDD.n2875 GND 0.01fF
C3433 VDD.n2876 GND 0.02fF
C3434 VDD.n2877 GND 0.02fF
C3435 VDD.n2878 GND 0.01fF
C3436 VDD.n2879 GND 0.01fF
C3437 VDD.n2880 GND 0.00fF
C3438 VDD.n2881 GND 0.00fF
C3439 VDD.n2882 GND 0.00fF
C3440 VDD.n2883 GND 0.00fF
C3441 VDD.n2884 GND 0.00fF
C3442 VDD.n2885 GND 0.00fF
C3443 VDD.n2886 GND 0.00fF
C3444 VDD.n2887 GND 0.00fF
C3445 VDD.n2888 GND 0.00fF
C3446 VDD.n2889 GND 0.00fF
C3447 VDD.n2890 GND 0.00fF
C3448 VDD.n2891 GND 0.00fF
C3449 VDD.n2892 GND 0.00fF
C3450 VDD.n2893 GND 0.00fF
C3451 VDD.n2894 GND 0.00fF
C3452 VDD.n2895 GND 0.00fF
C3453 VDD.n2896 GND 0.00fF
C3454 VDD.n2897 GND 0.00fF
C3455 VDD.n2898 GND 0.00fF
C3456 VDD.n2899 GND 0.00fF
C3457 VDD.n2900 GND 0.00fF
C3458 VDD.n2901 GND 0.00fF
C3459 VDD.n2902 GND 0.00fF
C3460 VDD.n2903 GND 0.00fF
C3461 VDD.n2904 GND 0.00fF
C3462 VDD.n2905 GND 0.00fF
C3463 VDD.n2906 GND 0.00fF
C3464 VDD.n2907 GND 0.00fF
C3465 VDD.n2908 GND 0.00fF
C3466 VDD.n2909 GND 0.00fF
C3467 VDD.n2910 GND 0.00fF
C3468 VDD.n2911 GND 0.00fF
C3469 VDD.n2912 GND 0.00fF
C3470 VDD.n2913 GND 0.00fF
C3471 VDD.n2914 GND 0.00fF
C3472 VDD.n2915 GND 0.00fF
C3473 VDD.n2916 GND 0.00fF
C3474 VDD.n2917 GND 0.00fF
C3475 VDD.n2918 GND 0.01fF
C3476 VDD.n2919 GND 0.00fF
C3477 VDD.n2920 GND 0.01fF
C3478 VDD.n2921 GND 0.00fF
C3479 VDD.n2922 GND 0.00fF
C3480 VDD.n2923 GND 0.00fF
C3481 VDD.n2924 GND 0.00fF
C3482 VDD.n2925 GND 0.01fF
C3483 VDD.n2926 GND 0.00fF
C3484 VDD.n2927 GND 0.01fF
C3485 VDD.n2928 GND 0.00fF
C3486 VDD.n2929 GND 0.00fF
C3487 VDD.n2930 GND 0.00fF
C3488 VDD.n2931 GND 0.00fF
C3489 VDD.n2932 GND 0.01fF
C3490 VDD.n2933 GND 0.00fF
C3491 VDD.n2934 GND 0.01fF
C3492 VDD.n2935 GND 0.00fF
C3493 VDD.n2936 GND 0.00fF
C3494 VDD.n2937 GND 0.00fF
C3495 VDD.n2938 GND 0.00fF
C3496 VDD.n2939 GND 0.01fF
C3497 VDD.n2940 GND 0.00fF
C3498 VDD.n2941 GND 0.01fF
C3499 VDD.n2942 GND 0.00fF
C3500 VDD.n2943 GND 0.00fF
C3501 VDD.n2944 GND 0.01fF
C3502 VDD.n2945 GND 0.01fF
C3503 VDD.n2946 GND 0.04fF
C3504 VDD.n2947 GND 0.01fF
C3505 VDD.n2948 GND 0.01fF
C3506 VDD.n2949 GND 0.01fF
C3507 VDD.n2950 GND 0.00fF
C3508 VDD.n2951 GND 0.00fF
C3509 VDD.n2952 GND 0.01fF
C3510 VDD.n2953 GND 0.00fF
C3511 VDD.n2954 GND 0.04fF
C3512 VDD.n2955 GND 0.01fF
C3513 VDD.n2956 GND 0.00fF
C3514 VDD.n2957 GND 0.01fF
C3515 VDD.n2958 GND 0.01fF
C3516 VDD.n2959 GND 0.00fF
C3517 VDD.n2960 GND 0.01fF
C3518 VDD.n2961 GND 0.01fF
C3519 VDD.n2962 GND 0.00fF
C3520 VDD.n2963 GND 0.01fF
C3521 VDD.n2964 GND 0.01fF
C3522 VDD.n2965 GND 0.00fF
C3523 VDD.n2966 GND 0.01fF
C3524 VDD.n2967 GND 0.01fF
C3525 VDD.n2968 GND 0.00fF
C3526 VDD.n2969 GND 0.01fF
C3527 VDD.n2970 GND 0.01fF
C3528 VDD.n2971 GND 0.00fF
C3529 VDD.n2972 GND 0.01fF
C3530 VDD.n2973 GND 0.01fF
C3531 VDD.n2974 GND 0.00fF
C3532 VDD.n2975 GND 0.01fF
C3533 VDD.n2976 GND 0.01fF
C3534 VDD.n2977 GND 0.00fF
C3535 VDD.n2978 GND 0.00fF
C3536 VDD.n2979 GND 0.01fF
C3537 VDD.n2980 GND 0.01fF
C3538 VDD.n2981 GND 0.01fF
C3539 VDD.n2982 GND 0.00fF
C3540 VDD.n2984 GND 0.00fF
C3541 VDD.n2985 GND 0.00fF
C3542 VDD.n2986 GND 0.00fF
C3543 VDD.n2987 GND 0.00fF
C3544 VDD.n2988 GND 0.00fF
C3545 VDD.n2989 GND 0.01fF
C3546 VDD.n2990 GND 0.01fF
C3547 VDD.n2991 GND 0.00fF
C3548 VDD.n2993 GND 0.01fF
C3549 VDD.n2995 GND 0.00fF
C3550 VDD.n2996 GND 0.00fF
C3551 VDD.n2997 GND 0.00fF
C3552 VDD.n2998 GND 0.00fF
C3553 VDD.n2999 GND 0.00fF
C3554 VDD.n3000 GND 0.00fF
C3555 VDD.n3001 GND 0.01fF
C3556 VDD.n3002 GND 0.01fF
C3557 VDD.n3004 GND 0.00fF
C3558 VDD.n3005 GND 0.00fF
C3559 VDD.n3006 GND 0.00fF
C3560 VDD.n3007 GND 0.01fF
C3561 VDD.n3008 GND 0.00fF
C3562 VDD.n3009 GND 0.00fF
C3563 VDD.n3010 GND 0.02fF
C3564 VDD.n3013 GND 0.01fF
C3565 VDD.n3014 GND 0.02fF
C3566 VDD.n3016 GND 0.01fF
C3567 VDD.n3017 GND 0.02fF
C3568 VDD.n3018 GND 0.01fF
C3569 VDD.n3019 GND 0.03fF
C3570 VDD.n3020 GND 0.01fF
C3571 VDD.n3021 GND 0.02fF
C3572 VDD.n3023 GND 0.01fF
C3573 VDD.n3025 GND 0.00fF
C3574 VDD.n3026 GND 0.00fF
C3575 VDD.n3027 GND 0.00fF
C3576 VDD.n3028 GND 0.00fF
C3577 VDD.n3029 GND 0.00fF
C3578 VDD.n3030 GND 0.00fF
C3579 VDD.n3031 GND 0.01fF
C3580 VDD.n3032 GND 0.01fF
C3581 VDD.n3034 GND 0.00fF
C3582 VDD.n3035 GND 0.00fF
C3583 VDD.n3036 GND 0.00fF
C3584 VDD.n3037 GND 0.00fF
C3585 VDD.n3038 GND 0.00fF
C3586 VDD.n3039 GND 0.00fF
C3587 VDD.n3040 GND 0.01fF
C3588 VDD.n3041 GND 0.00fF
C3589 VDD.n3042 GND 0.00fF
C3590 VDD.n3043 GND 0.00fF
C3591 VDD.n3044 GND 0.00fF
C3592 VDD.n3045 GND 0.00fF
C3593 VDD.n3046 GND 0.01fF
C3594 VDD.n3047 GND 0.01fF
C3595 VDD.n3048 GND 0.00fF
C3596 VDD.n3050 GND 0.00fF
C3597 VDD.n3051 GND 0.00fF
C3598 VDD.n3052 GND 0.00fF
C3599 VDD.n3053 GND 0.00fF
C3600 VDD.n3054 GND 0.00fF
C3601 VDD.n3055 GND 0.01fF
C3602 VDD.n3056 GND 0.01fF
C3603 VDD.n3057 GND 0.00fF
C3604 VDD.n3059 GND 0.94fF
C3605 VDD.n3060 GND 0.04fF
C3606 VDD.n3061 GND 0.02fF
C3607 VDD.n3062 GND 0.05fF
C3608 VDD.n3063 GND 0.04fF
C3609 VDD.n3064 GND 0.67fF
C3610 VDD.n3065 GND 0.04fF
C3611 VDD.n3066 GND 0.02fF
C3612 VDD.n3067 GND 0.01fF
C3613 VDD.n3068 GND 0.02fF
C3614 VDD.n3069 GND 0.01fF
C3615 VDD.n3070 GND 0.01fF
C3616 VDD.n3071 GND 0.04fF
C3617 VDD.t1 GND 0.35fF $ **FLOATING
C3618 VDD.n3072 GND 0.37fF
C3619 VDD.n3073 GND 0.02fF
C3620 VDD.n3074 GND 0.01fF
C3621 VDD.n3075 GND 0.03fF
C3622 VDD.t37 GND 0.04fF $ **FLOATING
C3623 VDD.n3076 GND 0.04fF
C3624 VDD.n3077 GND 0.02fF
C3625 VDD.n3078 GND 0.01fF
C3626 VDD.n3079 GND 0.03fF
C3627 VDD.n3080 GND 0.66fF
C3628 VDD.n3081 GND 0.02fF
C3629 VDD.n3082 GND 0.01fF
C3630 VDD.n3083 GND 0.04fF
C3631 VDD.n3084 GND 0.03fF
C3632 VDD.n3087 GND 0.35fF
C3633 VDD.n3088 GND 0.02fF
C3634 VDD.n3089 GND 0.01fF
C3635 VDD.n3090 GND 0.01fF
C3636 VDD.n3091 GND 0.01fF
C3637 VDD.n3092 GND 0.00fF
C3638 VDD.n3093 GND 0.00fF
C3639 VDD.n3094 GND 0.00fF
C3640 VDD.n3095 GND 0.00fF
C3641 VDD.n3096 GND 0.00fF
C3642 VDD.n3097 GND 0.01fF
C3643 VDD.n3098 GND 0.00fF
C3644 VDD.n3100 GND 0.01fF
C3645 VDD.n3101 GND 0.00fF
C3646 VDD.n3102 GND 0.01fF
C3647 VDD.n3103 GND 0.00fF
C3648 VDD.n3104 GND 0.01fF
C3649 VDD.n3105 GND 0.00fF
C3650 VDD.n3106 GND 0.00fF
C3651 VDD.n3107 GND 0.00fF
C3652 VDD.n3108 GND 0.00fF
C3653 VDD.n3109 GND 0.01fF
C3654 VDD.n3110 GND 0.00fF
C3655 VDD.n3112 GND 0.01fF
C3656 VDD.n3113 GND 0.00fF
C3657 VDD.n3114 GND 0.01fF
C3658 VDD.n3115 GND 0.00fF
C3659 VDD.n3116 GND 0.01fF
C3660 VDD.n3117 GND 0.00fF
C3661 VDD.n3118 GND 0.00fF
C3662 VDD.n3119 GND 0.00fF
C3663 VDD.n3120 GND 0.00fF
C3664 VDD.n3121 GND 0.01fF
C3665 VDD.n3122 GND 0.00fF
C3666 VDD.n3124 GND 0.01fF
C3667 VDD.n3125 GND 0.00fF
C3668 VDD.n3126 GND 0.01fF
C3669 VDD.n3127 GND 0.00fF
C3670 VDD.n3128 GND 0.01fF
C3671 VDD.n3129 GND 0.00fF
C3672 VDD.n3130 GND 0.00fF
C3673 VDD.n3131 GND 0.00fF
C3674 VDD.n3132 GND 0.00fF
C3675 VDD.n3133 GND 0.01fF
C3676 VDD.n3134 GND 0.00fF
C3677 VDD.n3136 GND 0.01fF
C3678 VDD.n3137 GND 0.00fF
C3679 VDD.n3138 GND 0.01fF
C3680 VDD.n3139 GND 0.00fF
C3681 VDD.n3140 GND 0.00fF
C3682 VDD.n3141 GND 0.01fF
C3683 VDD.n3143 GND 0.00fF
C3684 VDD.n3144 GND 0.01fF
C3685 VDD.n3145 GND 0.00fF
C3686 VDD.n3146 GND 0.01fF
C3687 VDD.n3147 GND 0.00fF
C3688 VDD.n3148 GND 0.00fF
C3689 VDD.n3149 GND 0.00fF
C3690 VDD.n3150 GND 0.01fF
C3691 VDD.n3151 GND 0.00fF
C3692 VDD.n3152 GND 0.00fF
C3693 VDD.n3153 GND 0.01fF
C3694 VDD.n3155 GND 0.00fF
C3695 VDD.n3156 GND 0.01fF
C3696 VDD.n3157 GND 0.00fF
C3697 VDD.n3158 GND 0.01fF
C3698 VDD.n3159 GND 0.00fF
C3699 VDD.n3160 GND 0.00fF
C3700 VDD.n3161 GND 0.00fF
C3701 VDD.n3162 GND 0.01fF
C3702 VDD.n3163 GND 0.00fF
C3703 VDD.n3164 GND 0.00fF
C3704 VDD.n3165 GND 0.01fF
C3705 VDD.n3167 GND 0.00fF
C3706 VDD.n3168 GND 0.01fF
C3707 VDD.n3169 GND 0.00fF
C3708 VDD.n3170 GND 0.01fF
C3709 VDD.n3171 GND 0.00fF
C3710 VDD.n3172 GND 0.00fF
C3711 VDD.n3173 GND 0.00fF
C3712 VDD.n3174 GND 0.01fF
C3713 VDD.n3175 GND 0.00fF
C3714 VDD.n3176 GND 0.00fF
C3715 VDD.n3177 GND 0.01fF
C3716 VDD.n3179 GND 0.00fF
C3717 VDD.n3180 GND 0.02fF
C3718 VDD.n3181 GND 0.00fF
C3719 VDD.n3182 GND 0.01fF
C3720 VDD.n3183 GND 0.00fF
C3721 VDD.n3184 GND 0.00fF
C3722 VDD.n3185 GND 0.01fF
C3723 VDD.n3186 GND 0.01fF
C3724 VDD.n3187 GND 0.04fF
C3725 VDD.n3189 GND 0.02fF
C3726 VDD.n3190 GND 0.01fF
C3727 VDD.n3191 GND 0.02fF
C3728 VDD.n3192 GND 0.02fF
C3729 VDD.n3193 GND 0.01fF
C3730 VDD.n3194 GND 0.01fF
C3731 VDD.n3195 GND 0.01fF
C3732 VDD.n3196 GND 0.01fF
C3733 VDD.n3197 GND 0.00fF
C3734 VDD.n3198 GND 0.00fF
C3735 VDD.n3199 GND 0.00fF
C3736 VDD.n3200 GND 0.00fF
C3737 VDD.n3201 GND 0.01fF
C3738 VDD.n3202 GND 0.00fF
C3739 VDD.n3204 GND 0.01fF
C3740 VDD.n3205 GND 0.00fF
C3741 VDD.n3206 GND 0.01fF
C3742 VDD.n3207 GND 0.00fF
C3743 VDD.n3208 GND 0.01fF
C3744 VDD.n3209 GND 0.00fF
C3745 VDD.n3210 GND 0.00fF
C3746 VDD.n3211 GND 0.00fF
C3747 VDD.n3212 GND 0.00fF
C3748 VDD.n3213 GND 0.01fF
C3749 VDD.n3215 GND 0.00fF
C3750 VDD.n3217 GND 0.01fF
C3751 VDD.n3218 GND 0.00fF
C3752 VDD.n3219 GND 0.01fF
C3753 VDD.n3220 GND 0.00fF
C3754 VDD.n3221 GND 0.01fF
C3755 VDD.n3222 GND 0.00fF
C3756 VDD.n3223 GND 0.00fF
C3757 VDD.n3224 GND 0.00fF
C3758 VDD.n3225 GND 0.00fF
C3759 VDD.n3226 GND 0.01fF
C3760 VDD.n3228 GND 0.00fF
C3761 VDD.n3229 GND 0.01fF
C3762 VDD.n3230 GND 0.00fF
C3763 VDD.n3231 GND 0.01fF
C3764 VDD.n3232 GND 0.00fF
C3765 VDD.n3233 GND 0.01fF
C3766 VDD.n3234 GND 0.00fF
C3767 VDD.n3235 GND 0.00fF
C3768 VDD.n3236 GND 0.00fF
C3769 VDD.n3237 GND 0.00fF
C3770 VDD.n3238 GND 0.01fF
C3771 VDD.n3240 GND 0.00fF
C3772 VDD.n3241 GND 0.01fF
C3773 VDD.n3242 GND 0.00fF
C3774 VDD.n3243 GND 0.01fF
C3775 VDD.n3244 GND 0.00fF
C3776 VDD.n3245 GND 0.00fF
C3777 VDD.n3246 GND 0.01fF
C3778 VDD.n3247 GND 0.00fF
C3779 VDD.n3249 GND 0.01fF
C3780 VDD.n3250 GND 0.00fF
C3781 VDD.n3251 GND 0.01fF
C3782 VDD.n3252 GND 0.00fF
C3783 VDD.n3253 GND 0.00fF
C3784 VDD.n3254 GND 0.00fF
C3785 VDD.n3255 GND 0.01fF
C3786 VDD.n3256 GND 0.00fF
C3787 VDD.n3257 GND 0.00fF
C3788 VDD.n3258 GND 0.01fF
C3789 VDD.n3259 GND 0.00fF
C3790 VDD.n3261 GND 0.01fF
C3791 VDD.n3262 GND 0.00fF
C3792 VDD.n3263 GND 0.01fF
C3793 VDD.n3264 GND 0.00fF
C3794 VDD.n3265 GND 0.00fF
C3795 VDD.n3266 GND 0.00fF
C3796 VDD.n3267 GND 0.01fF
C3797 VDD.n3268 GND 0.00fF
C3798 VDD.n3269 GND 0.00fF
C3799 VDD.n3270 GND 0.01fF
C3800 VDD.n3271 GND 0.00fF
C3801 VDD.n3273 GND 0.01fF
C3802 VDD.n3274 GND 0.00fF
C3803 VDD.n3275 GND 0.01fF
C3804 VDD.n3276 GND 0.00fF
C3805 VDD.n3277 GND 0.00fF
C3806 VDD.n3278 GND 0.00fF
C3807 VDD.n3279 GND 0.01fF
C3808 VDD.n3280 GND 0.00fF
C3809 VDD.n3281 GND 0.00fF
C3810 VDD.n3282 GND 0.01fF
C3811 VDD.n3283 GND 0.00fF
C3812 VDD.n3285 GND 0.01fF
C3813 VDD.n3286 GND 0.00fF
C3814 VDD.n3287 GND 0.01fF
C3815 VDD.n3288 GND 0.00fF
C3816 VDD.n3289 GND 0.00fF
C3817 VDD.n3290 GND 0.01fF
C3818 VDD.n3291 GND 0.00fF
C3819 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_13/BULK GND 0.02fF
C3820 VDD.n3292 GND 0.02fF
C3821 VDD.n3293 GND 0.01fF
C3822 VDD.n3294 GND 0.01fF
C3823 VDD.n3295 GND 0.03fF
C3824 VDD.n3296 GND 0.02fF
C3825 VDD.n3297 GND 0.01fF
C3826 VDD.n3298 GND 0.00fF
C3827 VDD.n3299 GND 0.00fF
C3828 VDD.n3300 GND 0.04fF
C3829 VDD.n3301 GND 0.01fF
C3830 VDD.n3302 GND 0.01fF
C3831 VDD.n3303 GND 0.01fF
C3832 VDD.n3304 GND 0.01fF
C3833 VDD.n3305 GND 0.01fF
C3834 VDD.n3306 GND 0.03fF
C3835 VDD.n3307 GND 0.04fF
C3836 VDD.n3308 GND 0.01fF
C3837 VDD.n3309 GND 0.01fF
C3838 VDD.n3310 GND 0.01fF
C3839 VDD.n3311 GND 0.00fF
C3840 VDD.n3312 GND 0.00fF
C3841 VDD.n3313 GND 0.01fF
C3842 VDD.n3314 GND 0.00fF
C3843 VDD.n3315 GND 0.02fF
C3844 VDD.n3316 GND 0.01fF
C3845 VDD.n3317 GND 0.01fF
C3846 VDD.n3318 GND 0.00fF
C3847 VDD.n3319 GND 0.00fF
C3848 VDD.n3320 GND 0.00fF
C3849 VDD.n3321 GND 0.00fF
C3850 VDD.n3322 GND 0.00fF
C3851 VDD.n3323 GND 0.01fF
C3852 VDD.n3325 GND 0.00fF
C3853 VDD.n3326 GND 0.01fF
C3854 VDD.n3327 GND 0.00fF
C3855 VDD.n3328 GND 0.01fF
C3856 VDD.n3329 GND 0.00fF
C3857 VDD.n3330 GND 0.01fF
C3858 VDD.n3331 GND 0.00fF
C3859 VDD.n3332 GND 0.00fF
C3860 VDD.n3333 GND 0.00fF
C3861 VDD.n3334 GND 0.00fF
C3862 VDD.n3335 GND 0.01fF
C3863 VDD.n3336 GND 0.00fF
C3864 VDD.n3338 GND 0.01fF
C3865 VDD.n3339 GND 0.00fF
C3866 VDD.n3340 GND 0.01fF
C3867 VDD.n3341 GND 0.00fF
C3868 VDD.n3342 GND 0.01fF
C3869 VDD.n3343 GND 0.00fF
C3870 VDD.n3344 GND 0.00fF
C3871 VDD.n3345 GND 0.00fF
C3872 VDD.n3346 GND 0.00fF
C3873 VDD.n3347 GND 0.01fF
C3874 VDD.n3349 GND 0.00fF
C3875 VDD.n3351 GND 0.01fF
C3876 VDD.n3352 GND 0.00fF
C3877 VDD.n3353 GND 0.01fF
C3878 VDD.n3354 GND 0.00fF
C3879 VDD.n3355 GND 0.01fF
C3880 VDD.n3356 GND 0.00fF
C3881 VDD.n3357 GND 0.00fF
C3882 VDD.n3358 GND 0.00fF
C3883 VDD.n3359 GND 0.00fF
C3884 VDD.n3360 GND 0.01fF
C3885 VDD.n3361 GND 0.00fF
C3886 VDD.n3363 GND 0.01fF
C3887 VDD.n3364 GND 0.00fF
C3888 VDD.n3365 GND 0.01fF
C3889 VDD.n3366 GND 0.00fF
C3890 VDD.n3367 GND 0.00fF
C3891 VDD.n3369 GND 0.01fF
C3892 VDD.n3370 GND 0.00fF
C3893 VDD.n3372 GND 0.01fF
C3894 VDD.n3373 GND 0.00fF
C3895 VDD.n3374 GND 0.01fF
C3896 VDD.n3375 GND 0.00fF
C3897 VDD.n3376 GND 0.00fF
C3898 VDD.n3377 GND 0.00fF
C3899 VDD.n3378 GND 0.01fF
C3900 VDD.n3379 GND 0.00fF
C3901 VDD.n3380 GND 0.00fF
C3902 VDD.n3381 GND 0.01fF
C3903 VDD.n3383 GND 0.00fF
C3904 VDD.n3385 GND 0.01fF
C3905 VDD.n3386 GND 0.00fF
C3906 VDD.n3387 GND 0.01fF
C3907 VDD.n3388 GND 0.00fF
C3908 VDD.n3389 GND 0.00fF
C3909 VDD.n3390 GND 0.00fF
C3910 VDD.n3391 GND 0.01fF
C3911 VDD.n3392 GND 0.00fF
C3912 VDD.n3393 GND 0.00fF
C3913 VDD.n3394 GND 0.01fF
C3914 VDD.n3395 GND 0.00fF
C3915 VDD.n3397 GND 0.01fF
C3916 VDD.n3398 GND 0.00fF
C3917 VDD.n3399 GND 0.01fF
C3918 VDD.n3400 GND 0.00fF
C3919 VDD.n3401 GND 0.00fF
C3920 VDD.n3402 GND 0.00fF
C3921 VDD.n3403 GND 0.01fF
C3922 VDD.n3404 GND 0.00fF
C3923 VDD.n3405 GND 0.00fF
C3924 VDD.n3406 GND 0.01fF
C3925 VDD.n3408 GND 0.00fF
C3926 VDD.n3409 GND 0.01fF
C3927 VDD.n3410 GND 0.00fF
C3928 VDD.n3411 GND 0.01fF
C3929 VDD.n3412 GND 0.00fF
C3930 VDD.n3413 GND 0.00fF
C3931 VDD.n3414 GND 0.01fF
C3932 VDD.n3415 GND 0.01fF
C3933 VDD.n3416 GND 0.04fF
C3934 VDD.n3417 GND 0.02fF
C3935 VDD.n3418 GND 0.05fF
C3936 VDD.n3419 GND 0.04fF
C3937 VDD.n3420 GND 0.04fF
C3938 VDD.n3421 GND 0.02fF
C3939 VDD.n3422 GND 0.02fF
C3940 VDD.n3423 GND 0.01fF
C3941 VDD.n3424 GND 0.03fF
C3942 VDD.n3425 GND 0.01fF
C3943 VDD.n3426 GND 0.01fF
C3944 VDD.n3427 GND 0.03fF
C3945 VDD.n3428 GND 0.02fF
C3946 VDD.n3429 GND 0.01fF
C3947 VDD.n3430 GND 0.03fF
C3948 VDD.t0 GND 0.04fF $ **FLOATING
C3949 VDD.n3431 GND 0.04fF
C3950 VDD.n3432 GND 0.02fF
C3951 VDD.n3433 GND 0.01fF
C3952 VDD.n3434 GND 0.03fF
C3953 VDD.n3435 GND 0.02fF
C3954 VDD.n3436 GND 0.01fF
C3955 VDD.n3437 GND 0.04fF
C3956 VDD.n3438 GND 0.03fF
C3957 VDD.n3439 GND 0.01fF
C3958 VDD.n3440 GND 0.02fF
C3959 VDD.n3441 GND 0.01fF
C3960 VDD.n3442 GND 0.01fF
C3961 VDD.n3443 GND 0.02fF
C3962 VDD.n3444 GND 0.02fF
C3963 VDD.n3445 GND 0.01fF
C3964 VDD.n3446 GND 0.02fF
C3965 VDD.n3447 GND 0.02fF
C3966 VDD.n3448 GND 0.01fF
C3967 VDD.n3449 GND 0.02fF
C3968 VDD.n3450 GND 0.02fF
C3969 VDD.n3451 GND 0.01fF
C3970 VDD.n3452 GND 0.02fF
C3971 VDD.n3453 GND 0.02fF
C3972 VDD.n3454 GND 0.01fF
C3973 VDD.n3455 GND 0.02fF
C3974 VDD.n3456 GND 0.02fF
C3975 VDD.n3457 GND 0.02fF
C3976 VDD.n3458 GND 0.01fF
C3977 VDD.n3459 GND 0.01fF
C3978 VDD.n3460 GND 0.00fF
C3979 VDD.n3461 GND 0.00fF
C3980 VDD.n3462 GND 0.00fF
C3981 VDD.n3463 GND 0.00fF
C3982 VDD.n3464 GND 0.01fF
C3983 VDD.n3465 GND 0.00fF
C3984 VDD.n3466 GND 0.01fF
C3985 VDD.n3467 GND 0.00fF
C3986 VDD.n3468 GND 0.01fF
C3987 VDD.n3469 GND 0.00fF
C3988 VDD.n3470 GND 0.01fF
C3989 VDD.n3471 GND 0.00fF
C3990 VDD.n3472 GND 0.00fF
C3991 VDD.n3473 GND 0.00fF
C3992 VDD.n3474 GND 0.00fF
C3993 VDD.n3475 GND 0.01fF
C3994 VDD.n3477 GND 0.00fF
C3995 VDD.n3479 GND 0.01fF
C3996 VDD.n3480 GND 0.00fF
C3997 VDD.n3481 GND 0.01fF
C3998 VDD.n3482 GND 0.00fF
C3999 VDD.n3483 GND 0.01fF
C4000 VDD.n3484 GND 0.00fF
C4001 VDD.n3485 GND 0.00fF
C4002 VDD.n3486 GND 0.00fF
C4003 VDD.n3487 GND 0.00fF
C4004 VDD.n3488 GND 0.01fF
C4005 VDD.n3490 GND 0.00fF
C4006 VDD.n3491 GND 0.01fF
C4007 VDD.n3492 GND 0.00fF
C4008 VDD.n3493 GND 0.01fF
C4009 VDD.n3494 GND 0.00fF
C4010 VDD.n3495 GND 0.01fF
C4011 VDD.n3496 GND 0.00fF
C4012 VDD.n3497 GND 0.00fF
C4013 VDD.n3498 GND 0.00fF
C4014 VDD.n3499 GND 0.00fF
C4015 VDD.n3500 GND 0.01fF
C4016 VDD.n3502 GND 0.00fF
C4017 VDD.n3503 GND 0.01fF
C4018 VDD.n3504 GND 0.00fF
C4019 VDD.n3505 GND 0.01fF
C4020 VDD.n3506 GND 0.00fF
C4021 VDD.n3507 GND 0.00fF
C4022 VDD.n3508 GND 0.01fF
C4023 VDD.n3509 GND 0.00fF
C4024 VDD.n3511 GND 0.01fF
C4025 VDD.n3512 GND 0.00fF
C4026 VDD.n3513 GND 0.01fF
C4027 VDD.n3514 GND 0.00fF
C4028 VDD.n3515 GND 0.00fF
C4029 VDD.n3516 GND 0.00fF
C4030 VDD.n3517 GND 0.01fF
C4031 VDD.n3518 GND 0.00fF
C4032 VDD.n3519 GND 0.00fF
C4033 VDD.n3520 GND 0.01fF
C4034 VDD.n3521 GND 0.00fF
C4035 VDD.n3523 GND 0.01fF
C4036 VDD.n3524 GND 0.00fF
C4037 VDD.n3525 GND 0.01fF
C4038 VDD.n3526 GND 0.00fF
C4039 VDD.n3527 GND 0.00fF
C4040 VDD.n3528 GND 0.00fF
C4041 VDD.n3529 GND 0.01fF
C4042 VDD.n3530 GND 0.00fF
C4043 VDD.n3531 GND 0.00fF
C4044 VDD.n3532 GND 0.01fF
C4045 VDD.n3533 GND 0.00fF
C4046 VDD.n3535 GND 0.01fF
C4047 VDD.n3536 GND 0.00fF
C4048 VDD.n3537 GND 0.01fF
C4049 VDD.n3538 GND 0.00fF
C4050 VDD.n3539 GND 0.00fF
C4051 VDD.n3540 GND 0.00fF
C4052 VDD.n3541 GND 0.01fF
C4053 VDD.n3542 GND 0.00fF
C4054 VDD.n3543 GND 0.00fF
C4055 VDD.n3544 GND 0.01fF
C4056 VDD.n3545 GND 0.00fF
C4057 VDD.n3547 GND 0.01fF
C4058 VDD.n3548 GND 0.00fF
C4059 VDD.n3549 GND 0.01fF
C4060 VDD.n3550 GND 0.00fF
C4061 VDD.n3551 GND 0.00fF
C4062 VDD.n3552 GND 0.01fF
C4063 VDD.n3553 GND 0.00fF
C4064 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/BULK GND 0.01fF
C4065 VDD.n3554 GND 0.02fF
C4066 VDD.n3555 GND 0.02fF
C4067 VDD.n3556 GND 0.02fF
C4068 VDD.n3557 GND 0.02fF
C4069 VDD.n3558 GND 0.01fF
C4070 VDD.n3559 GND 0.00fF
C4071 VDD.n3560 GND 0.01fF
C4072 VDD.n3561 GND 0.01fF
C4073 VDD.n3562 GND 0.00fF
C4074 VDD.n3563 GND 0.01fF
C4075 VDD.n3564 GND 0.01fF
C4076 VDD.n3565 GND 0.00fF
C4077 VDD.n3566 GND 0.01fF
C4078 VDD.n3567 GND 0.01fF
C4079 VDD.n3568 GND 0.00fF
C4080 VDD.n3569 GND 0.01fF
C4081 VDD.n3570 GND 0.01fF
C4082 VDD.n3571 GND 0.00fF
C4083 VDD.n3572 GND 0.01fF
C4084 VDD.n3573 GND 0.01fF
C4085 VDD.n3574 GND 0.00fF
C4086 VDD.n3575 GND 0.01fF
C4087 VDD.n3576 GND 0.01fF
C4088 VDD.n3577 GND 0.00fF
C4089 VDD.n3578 GND 0.01fF
C4090 VDD.n3579 GND 0.01fF
C4091 VDD.n3580 GND 0.00fF
C4092 VDD.n3581 GND 0.00fF
C4093 VDD.n3582 GND 0.01fF
C4094 VDD.n3583 GND 0.01fF
C4095 VDD.n3584 GND 0.02fF
C4096 VDD.n3585 GND 0.02fF
C4097 VDD.n3586 GND 0.02fF
C4098 VDD.n3587 GND 0.42fF
C4099 VDD.n3588 GND 0.01fF
C4100 VDD.n3589 GND 0.01fF
C4101 VDD.n3590 GND 0.01fF
C4102 VDD.n3591 GND 0.01fF
C4103 VDD.n3592 GND 0.60fF
C4104 VDD.n3593 GND 0.02fF
C4105 VDD.n3594 GND 0.01fF
C4106 VDD.n3595 GND 0.02fF
C4107 VDD.t41 GND 0.35fF $ **FLOATING
C4108 VDD.n3596 GND 0.38fF
C4109 VDD.n3597 GND 0.02fF
C4110 VDD.n3598 GND 0.01fF
C4111 VDD.n3599 GND 0.02fF
C4112 VDD.t48 GND 0.35fF $ **FLOATING
C4113 VDD.n3600 GND 0.42fF
C4114 VDD.n3601 GND 0.02fF
C4115 VDD.n3602 GND 0.01fF
C4116 VDD.n3603 GND 0.02fF
C4117 VDD.n3604 GND 0.60fF
C4118 VDD.n3605 GND 0.02fF
C4119 VDD.n3606 GND 0.01fF
C4120 VDD.n3607 GND 0.02fF
C4121 VDD.n3608 GND 0.03fF
C4122 VDD.n3609 GND 0.01fF
C4123 VDD.n3610 GND 0.02fF
C4124 VDD.n3611 GND 0.45fF
C4125 VDD.n3612 GND 0.01fF
C4126 VDD.n3613 GND 0.01fF
C4127 VDD.n3614 GND 0.03fF
C4128 VDD.n3615 GND 0.58fF
C4129 VDD.n3616 GND 0.02fF
C4130 VDD.n3617 GND 0.01fF
C4131 VDD.n3618 GND 0.00fF
C4132 VDD.n3619 GND 0.02fF
C4133 VDD.t30 GND 0.04fF $ **FLOATING
C4134 VDD.n3620 GND 0.04fF
C4135 VDD.n3621 GND 0.02fF
C4136 VDD.n3622 GND 0.02fF
C4137 VDD.t31 GND 0.35fF $ **FLOATING
C4138 VDD.n3623 GND 0.38fF
C4139 VDD.n3624 GND 0.02fF
C4140 VDD.n3625 GND 0.01fF
C4141 VDD.n3626 GND 0.02fF
C4142 VDD.n3627 GND 0.01fF
C4143 VDD.n3628 GND 0.02fF
C4144 VDD.n3629 GND 0.02fF
C4145 VDD.n3630 GND 0.02fF
C4146 VDD.n3631 GND 0.01fF
C4147 VDD.n3632 GND 0.07fF
C4148 VDD.n3633 GND 0.05fF
C4149 VDD.n3634 GND 0.02fF
C4150 VDD.n3635 GND 0.03fF
C4151 VDD.n3636 GND 0.00fF
C4152 VDD.n3637 GND 0.01fF
C4153 VDD.n3638 GND 0.01fF
C4154 VDD.n3639 GND 0.01fF
C4155 VDD.n3640 GND 0.03fF
C4156 VDD.n3641 GND 0.01fF
C4157 VDD.n3642 GND 0.00fF
C4158 VDD.n3643 GND 0.01fF
C4159 VDD.n3644 GND 0.01fF
C4160 VDD.n3645 GND 0.03fF
C4161 VDD.n3646 GND 0.05fF
C4162 VDD.n3647 GND 0.10fF
C4163 VDD.n3648 GND 0.04fF
C4164 VDD.n3649 GND 0.04fF
C4165 VDD.n3650 GND 0.03fF
C4166 VDD.n3651 GND 0.01fF
C4167 VDD.n3652 GND 0.00fF
C4168 VDD.n3653 GND 0.00fF
C4169 VDD.n3654 GND 0.01fF
C4170 VDD.n3655 GND 0.01fF
C4171 VDD.n3656 GND 0.01fF
C4172 VDD.n3657 GND 0.03fF
C4173 VDD.n3658 GND 0.01fF
C4174 VDD.n3659 GND 0.01fF
C4175 VDD.n3660 GND 0.00fF
C4176 VDD.n3661 GND 0.01fF
C4177 VDD.n3662 GND 0.01fF
C4178 VDD.n3663 GND 0.05fF
C4179 VDD.n3665 GND 1.53fF
C4180 VDD.n3666 GND 1.52fF
C4181 VDD.n3668 GND 0.03fF
C4182 VDD.n3669 GND 0.01fF
C4183 VDD.n3670 GND 0.05fF
C4184 VDD.n3671 GND 0.02fF
C4185 VDD.n3672 GND 0.00fF
C4186 VDD.n3673 GND 0.01fF
C4187 VDD.n3674 GND 0.01fF
C4188 VDD.n3675 GND 0.05fF
C4189 VDD.n3676 GND 0.07fF
C4190 VDD.n3677 GND 0.20fF
C4191 VDD.n3678 GND 0.03fF
C4192 VDD.n3679 GND 0.00fF
C4193 VDD.n3680 GND 0.01fF
C4194 VDD.n3681 GND 0.01fF
C4195 VDD.n3682 GND 0.01fF
C4196 VDD.n3683 GND 0.03fF
C4197 VDD.n3684 GND 0.01fF
C4198 VDD.n3685 GND 0.01fF
C4199 VDD.n3686 GND 0.00fF
C4200 VDD.n3687 GND 0.00fF
C4201 VDD.n3688 GND 0.01fF
C4202 VDD.n3689 GND 0.01fF
C4203 VDD.n3690 GND 0.04fF
C4204 VDD.n3691 GND 0.05fF
C4205 VDD.n3693 GND 0.20fF
C4206 VDD.n3695 GND 0.20fF
C4207 VDD.n3696 GND 0.00fF
C4208 VDD.n3697 GND 0.19fF
C4209 VDD.n3699 GND 0.09fF
C4210 VDD.n3700 GND 0.09fF
C4211 VDD.n3701 GND 0.09fF
C4212 VDD.n3702 GND 0.09fF
C4213 VDD.n3703 GND 0.00fF
C4214 VDD.n3704 GND 0.09fF
C4215 VDD.n3705 GND 0.02fF
C4216 VDD.n3706 GND 0.01fF
C4217 VDD.n3707 GND 0.01fF
C4218 VDD.n3709 GND 0.01fF
C4219 VDD.n3710 GND 0.01fF
C4220 VDD.n3711 GND 0.01fF
C4221 VDD.n3713 GND 0.01fF
C4222 VDD.n3714 GND 0.01fF
C4223 VDD.n3715 GND 0.01fF
C4224 VDD.n3716 GND 0.01fF
C4225 VDD.n3717 GND 0.01fF
C4226 VDD.n3718 GND 0.01fF
C4227 VDD.n3719 GND 0.01fF
C4228 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/SOURCE GND 0.01fF
C4229 VDD.n3720 GND 0.01fF
C4230 VDD.n3721 GND 0.01fF
C4231 VDD.n3722 GND 0.01fF
C4232 VDD.n3723 GND 0.00fF
C4233 VDD.n3724 GND 0.01fF
C4234 VDD.n3725 GND 0.00fF
C4235 VDD.n3726 GND 0.01fF
C4236 VDD.n3727 GND 0.01fF
C4237 VDD.n3728 GND 0.01fF
C4238 VDD.n3729 GND 0.01fF
C4239 VDD.n3730 GND 0.01fF
C4240 VDD.n3731 GND 0.01fF
C4241 VDD.n3732 GND 0.00fF
C4242 VDD.n3733 GND 0.00fF
C4243 VDD.n3734 GND 0.00fF
C4244 VDD.n3735 GND 0.00fF
C4245 VDD.n3736 GND 0.00fF
C4246 VDD.n3737 GND 0.00fF
C4247 VDD.n3738 GND 0.00fF
C4248 VDD.n3739 GND 0.00fF
C4249 VDD.n3740 GND 0.00fF
C4250 VDD.n3741 GND 0.00fF
C4251 VDD.n3742 GND 0.00fF
C4252 VDD.n3743 GND 0.00fF
C4253 VDD.n3744 GND 0.00fF
C4254 VDD.n3745 GND 0.00fF
C4255 VDD.n3746 GND 0.00fF
C4256 VDD.n3747 GND 0.00fF
C4257 VDD.n3748 GND 0.00fF
C4258 VDD.n3749 GND 0.00fF
C4259 VDD.n3750 GND 0.00fF
C4260 VDD.t47 GND 0.04fF $ **FLOATING
C4261 VDD.n3751 GND 0.13fF
C4262 VDD.n3752 GND 0.00fF
C4263 VDD.n3753 GND 0.04fF
C4264 VDD.n3754 GND 0.07fF
C4265 VDD.n3755 GND 0.00fF
C4266 VDD.n3756 GND 0.00fF
C4267 VDD.n3757 GND 0.00fF
C4268 VDD.n3758 GND 0.00fF
C4269 VDD.n3759 GND 0.00fF
C4270 VDD.n3760 GND 0.00fF
C4271 VDD.n3761 GND 0.00fF
C4272 VDD.n3762 GND 0.00fF
C4273 VDD.n3763 GND 0.00fF
C4274 VDD.n3764 GND 0.00fF
C4275 VDD.n3765 GND 0.00fF
C4276 VDD.n3766 GND 0.00fF
C4277 VDD.n3767 GND 0.00fF
C4278 VDD.n3768 GND 0.00fF
C4279 VDD.n3769 GND 0.00fF
C4280 VDD.n3770 GND 0.00fF
C4281 VDD.n3771 GND 0.00fF
C4282 VDD.n3772 GND 0.01fF
C4283 VDD.n3773 GND 0.01fF
C4284 VDD.n3774 GND 0.00fF
C4285 VDD.n3775 GND 0.00fF
C4286 VDD.n3776 GND 0.00fF
C4287 VDD.n3777 GND 0.00fF
C4288 VDD.n3778 GND 0.00fF
C4289 VDD.n3779 GND 0.00fF
C4290 VDD.n3780 GND 0.00fF
C4291 VDD.n3781 GND 0.00fF
C4292 VDD.n3782 GND 0.00fF
C4293 VDD.n3783 GND 0.00fF
C4294 VDD.n3784 GND 0.00fF
C4295 VDD.n3785 GND 0.00fF
C4296 VDD.n3786 GND 0.00fF
C4297 VDD.n3787 GND 0.00fF
C4298 VDD.n3788 GND 0.00fF
C4299 VDD.n3789 GND 0.00fF
C4300 VDD.n3790 GND 0.00fF
C4301 VDD.n3791 GND 0.00fF
C4302 VDD.n3792 GND 0.00fF
C4303 VDD.t56 GND 0.04fF $ **FLOATING
C4304 VDD.n3793 GND 0.13fF
C4305 VDD.n3794 GND 0.00fF
C4306 VDD.n3795 GND 0.04fF
C4307 VDD.n3796 GND 0.07fF
C4308 VDD.n3797 GND 0.00fF
C4309 VDD.n3798 GND 0.00fF
C4310 VDD.n3799 GND 0.00fF
C4311 VDD.n3800 GND 0.00fF
C4312 VDD.n3801 GND 0.00fF
C4313 VDD.n3802 GND 0.00fF
C4314 VDD.n3803 GND 0.00fF
C4315 VDD.n3804 GND 0.00fF
C4316 VDD.n3805 GND 0.00fF
C4317 VDD.n3806 GND 0.00fF
C4318 VDD.n3807 GND 0.00fF
C4319 VDD.n3808 GND 0.00fF
C4320 VDD.n3809 GND 0.00fF
C4321 VDD.n3810 GND 0.00fF
C4322 VDD.n3811 GND 0.00fF
C4323 VDD.n3812 GND 0.00fF
C4324 VDD.n3813 GND 0.00fF
C4325 VDD.n3814 GND 0.02fF
C4326 VDD.n3816 GND 0.02fF
C4327 VDD.n3817 GND 0.01fF
C4328 VDD.n3818 GND 0.01fF
C4329 VDD.n3820 GND 0.01fF
C4330 VDD.n3821 GND 0.01fF
C4331 VDD.n3822 GND 0.01fF
C4332 VDD.n3824 GND 0.01fF
C4333 VDD.n3825 GND 0.01fF
C4334 VDD.n3826 GND 0.01fF
C4335 VDD.n3827 GND 0.01fF
C4336 VDD.n3828 GND 0.01fF
C4337 VDD.n3829 GND 0.01fF
C4338 VDD.n3830 GND 0.01fF
C4339 VDD.n3831 GND 0.01fF
C4340 VDD.n3832 GND 0.01fF
C4341 VDD.n3833 GND 0.00fF
C4342 VDD.n3834 GND 0.00fF
C4343 VDD.n3835 GND 0.00fF
C4344 VDD.n3836 GND 0.00fF
C4345 VDD.n3837 GND 0.00fF
C4346 VDD.n3838 GND 0.00fF
C4347 VDD.n3839 GND 0.00fF
C4348 VDD.n3840 GND 0.00fF
C4349 VDD.n3841 GND 0.00fF
C4350 VDD.n3842 GND 0.00fF
C4351 VDD.n3843 GND 0.00fF
C4352 VDD.n3844 GND 0.00fF
C4353 VDD.n3845 GND 0.00fF
C4354 VDD.n3846 GND 0.00fF
C4355 VDD.n3847 GND 0.00fF
C4356 VDD.n3848 GND 0.00fF
C4357 VDD.n3849 GND 0.00fF
C4358 VDD.n3850 GND 0.00fF
C4359 VDD.n3851 GND 0.00fF
C4360 VDD.t64 GND 0.04fF $ **FLOATING
C4361 VDD.n3852 GND 0.13fF
C4362 VDD.n3853 GND 0.00fF
C4363 VDD.n3854 GND 0.04fF
C4364 VDD.n3855 GND 0.07fF
C4365 VDD.n3856 GND 0.00fF
C4366 VDD.n3857 GND 0.00fF
C4367 VDD.n3858 GND 0.00fF
C4368 VDD.n3859 GND 0.00fF
C4369 VDD.n3860 GND 0.00fF
C4370 VDD.n3861 GND 0.00fF
C4371 VDD.n3862 GND 0.00fF
C4372 VDD.n3863 GND 0.00fF
C4373 VDD.n3864 GND 0.00fF
C4374 VDD.n3865 GND 0.00fF
C4375 VDD.n3866 GND 0.00fF
C4376 VDD.n3867 GND 0.00fF
C4377 VDD.n3868 GND 0.00fF
C4378 VDD.n3869 GND 0.00fF
C4379 VDD.n3870 GND 0.00fF
C4380 VDD.n3871 GND 0.00fF
C4381 VDD.n3872 GND 0.00fF
C4382 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/SOURCE GND 0.01fF
C4383 VDD.n3873 GND 0.01fF
C4384 VDD.n3874 GND 0.01fF
C4385 VDD.n3875 GND 0.01fF
C4386 VDD.n3876 GND 0.00fF
C4387 VDD.n3877 GND 0.01fF
C4388 VDD.n3878 GND 0.00fF
C4389 VDD.n3879 GND 0.01fF
C4390 VDD.n3880 GND 0.01fF
C4391 VDD.n3881 GND 0.01fF
C4392 VDD.n3882 GND 0.01fF
C4393 VDD.n3883 GND 0.01fF
C4394 VDD.n3884 GND 0.01fF
C4395 VDD.n3885 GND 0.00fF
C4396 VDD.n3886 GND 0.00fF
C4397 VDD.n3887 GND 0.00fF
C4398 VDD.n3888 GND 0.00fF
C4399 VDD.n3889 GND 0.00fF
C4400 VDD.n3890 GND 0.00fF
C4401 VDD.n3891 GND 0.00fF
C4402 VDD.n3892 GND 0.00fF
C4403 VDD.n3893 GND 0.00fF
C4404 VDD.n3894 GND 0.00fF
C4405 VDD.n3895 GND 0.00fF
C4406 VDD.n3896 GND 0.00fF
C4407 VDD.n3897 GND 0.00fF
C4408 VDD.n3898 GND 0.00fF
C4409 VDD.n3899 GND 0.00fF
C4410 VDD.n3900 GND 0.00fF
C4411 VDD.n3901 GND 0.00fF
C4412 VDD.n3902 GND 0.00fF
C4413 VDD.n3903 GND 0.00fF
C4414 VDD.t52 GND 0.04fF $ **FLOATING
C4415 VDD.n3904 GND 0.13fF
C4416 VDD.n3905 GND 0.00fF
C4417 VDD.n3906 GND 0.04fF
C4418 VDD.n3907 GND 0.07fF
C4419 VDD.n3908 GND 0.00fF
C4420 VDD.n3909 GND 0.00fF
C4421 VDD.n3910 GND 0.00fF
C4422 VDD.n3911 GND 0.00fF
C4423 VDD.n3912 GND 0.00fF
C4424 VDD.n3913 GND 0.00fF
C4425 VDD.n3914 GND 0.00fF
C4426 VDD.n3915 GND 0.00fF
C4427 VDD.n3916 GND 0.00fF
C4428 VDD.n3917 GND 0.00fF
C4429 VDD.n3918 GND 0.00fF
C4430 VDD.n3919 GND 0.00fF
C4431 VDD.n3920 GND 0.00fF
C4432 VDD.n3921 GND 0.00fF
C4433 VDD.n3922 GND 0.00fF
C4434 VDD.n3923 GND 0.00fF
C4435 VDD.n3924 GND 0.00fF
C4436 VDD.n3925 GND 0.02fF
C4437 VDD.n3927 GND 0.02fF
C4438 VDD.n3928 GND 0.01fF
C4439 VDD.n3929 GND 0.01fF
C4440 VDD.n3931 GND 0.01fF
C4441 VDD.n3932 GND 0.01fF
C4442 VDD.n3933 GND 0.01fF
C4443 VDD.n3935 GND 0.01fF
C4444 VDD.n3936 GND 0.01fF
C4445 VDD.n3937 GND 0.01fF
C4446 VDD.n3938 GND 0.01fF
C4447 VDD.n3939 GND 0.01fF
C4448 VDD.n3940 GND 0.01fF
C4449 VDD.n3941 GND 0.01fF
C4450 VDD.n3942 GND 0.01fF
C4451 VDD.n3943 GND 0.01fF
C4452 VDD.n3944 GND 0.00fF
C4453 VDD.n3945 GND 0.00fF
C4454 VDD.n3946 GND 0.00fF
C4455 VDD.n3947 GND 0.00fF
C4456 VDD.n3948 GND 0.00fF
C4457 VDD.n3949 GND 0.00fF
C4458 VDD.n3950 GND 0.00fF
C4459 VDD.n3951 GND 0.00fF
C4460 VDD.n3952 GND 0.00fF
C4461 VDD.n3953 GND 0.00fF
C4462 VDD.n3954 GND 0.00fF
C4463 VDD.n3955 GND 0.00fF
C4464 VDD.n3956 GND 0.00fF
C4465 VDD.n3957 GND 0.00fF
C4466 VDD.n3958 GND 0.00fF
C4467 VDD.n3959 GND 0.00fF
C4468 VDD.n3960 GND 0.00fF
C4469 VDD.n3961 GND 0.00fF
C4470 VDD.n3962 GND 0.00fF
C4471 VDD.t66 GND 0.04fF $ **FLOATING
C4472 VDD.n3963 GND 0.13fF
C4473 VDD.n3964 GND 0.00fF
C4474 VDD.n3965 GND 0.04fF
C4475 VDD.n3966 GND 0.07fF
C4476 VDD.n3967 GND 0.00fF
C4477 VDD.n3968 GND 0.00fF
C4478 VDD.n3969 GND 0.00fF
C4479 VDD.n3970 GND 0.00fF
C4480 VDD.n3971 GND 0.00fF
C4481 VDD.n3972 GND 0.00fF
C4482 VDD.n3973 GND 0.00fF
C4483 VDD.n3974 GND 0.00fF
C4484 VDD.n3975 GND 0.00fF
C4485 VDD.n3976 GND 0.00fF
C4486 VDD.n3977 GND 0.00fF
C4487 VDD.n3978 GND 0.00fF
C4488 VDD.n3979 GND 0.00fF
C4489 VDD.n3980 GND 0.00fF
C4490 VDD.n3981 GND 0.00fF
C4491 VDD.n3982 GND 0.00fF
C4492 VDD.n3983 GND 0.00fF
C4493 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/SOURCE GND 0.01fF
C4494 VDD.n3984 GND 0.01fF
C4495 VDD.n3985 GND 0.01fF
C4496 VDD.n3986 GND 0.01fF
C4497 VDD.n3987 GND 0.00fF
C4498 VDD.n3988 GND 0.01fF
C4499 VDD.n3989 GND 0.00fF
C4500 VDD.n3990 GND 0.01fF
C4501 VDD.n3991 GND 0.01fF
C4502 VDD.n3992 GND 0.01fF
C4503 VDD.n3993 GND 0.01fF
C4504 VDD.n3994 GND 0.01fF
C4505 VDD.n3995 GND 0.01fF
C4506 VDD.n3996 GND 0.00fF
C4507 VDD.n3997 GND 0.00fF
C4508 VDD.n3998 GND 0.00fF
C4509 VDD.n3999 GND 0.00fF
C4510 VDD.n4000 GND 0.00fF
C4511 VDD.n4001 GND 0.00fF
C4512 VDD.n4002 GND 0.00fF
C4513 VDD.n4003 GND 0.00fF
C4514 VDD.n4004 GND 0.00fF
C4515 VDD.n4005 GND 0.00fF
C4516 VDD.n4006 GND 0.00fF
C4517 VDD.n4007 GND 0.00fF
C4518 VDD.n4008 GND 0.00fF
C4519 VDD.n4009 GND 0.00fF
C4520 VDD.n4010 GND 0.00fF
C4521 VDD.n4011 GND 0.00fF
C4522 VDD.n4012 GND 0.00fF
C4523 VDD.n4013 GND 0.00fF
C4524 VDD.n4014 GND 0.00fF
C4525 VDD.t63 GND 0.04fF $ **FLOATING
C4526 VDD.n4015 GND 0.13fF
C4527 VDD.n4016 GND 0.00fF
C4528 VDD.n4017 GND 0.04fF
C4529 VDD.n4018 GND 0.07fF
C4530 VDD.n4019 GND 0.00fF
C4531 VDD.n4020 GND 0.00fF
C4532 VDD.n4021 GND 0.00fF
C4533 VDD.n4022 GND 0.00fF
C4534 VDD.n4023 GND 0.00fF
C4535 VDD.n4024 GND 0.00fF
C4536 VDD.n4025 GND 0.00fF
C4537 VDD.n4026 GND 0.00fF
C4538 VDD.n4027 GND 0.00fF
C4539 VDD.n4028 GND 0.00fF
C4540 VDD.n4029 GND 0.00fF
C4541 VDD.n4030 GND 0.00fF
C4542 VDD.n4031 GND 0.00fF
C4543 VDD.n4032 GND 0.00fF
C4544 VDD.n4033 GND 0.00fF
C4545 VDD.n4034 GND 0.00fF
C4546 VDD.n4035 GND 0.00fF
C4547 VDD.n4036 GND 0.02fF
C4548 VDD.n4038 GND 0.02fF
C4549 VDD.n4039 GND 0.01fF
C4550 VDD.n4040 GND 0.01fF
C4551 VDD.n4042 GND 0.01fF
C4552 VDD.n4043 GND 0.01fF
C4553 VDD.n4044 GND 0.01fF
C4554 VDD.n4046 GND 0.01fF
C4555 VDD.n4047 GND 0.01fF
C4556 VDD.n4048 GND 0.01fF
C4557 VDD.n4049 GND 0.01fF
C4558 VDD.n4050 GND 0.01fF
C4559 VDD.n4051 GND 0.01fF
C4560 VDD.n4052 GND 0.01fF
C4561 VDD.n4053 GND 0.01fF
C4562 VDD.n4054 GND 0.01fF
C4563 VDD.n4055 GND 0.00fF
C4564 VDD.n4056 GND 0.00fF
C4565 VDD.n4057 GND 0.00fF
C4566 VDD.n4058 GND 0.00fF
C4567 VDD.n4059 GND 0.00fF
C4568 VDD.n4060 GND 0.00fF
C4569 VDD.n4061 GND 0.00fF
C4570 VDD.n4062 GND 0.00fF
C4571 VDD.n4063 GND 0.00fF
C4572 VDD.n4064 GND 0.00fF
C4573 VDD.n4065 GND 0.00fF
C4574 VDD.n4066 GND 0.00fF
C4575 VDD.n4067 GND 0.00fF
C4576 VDD.n4068 GND 0.00fF
C4577 VDD.n4069 GND 0.00fF
C4578 VDD.n4070 GND 0.00fF
C4579 VDD.n4071 GND 0.00fF
C4580 VDD.n4072 GND 0.00fF
C4581 VDD.n4073 GND 0.00fF
C4582 VDD.t44 GND 0.04fF $ **FLOATING
C4583 VDD.n4074 GND 0.13fF
C4584 VDD.n4075 GND 0.00fF
C4585 VDD.n4076 GND 0.04fF
C4586 VDD.n4077 GND 0.07fF
C4587 VDD.n4078 GND 0.00fF
C4588 VDD.n4079 GND 0.00fF
C4589 VDD.n4080 GND 0.00fF
C4590 VDD.n4081 GND 0.00fF
C4591 VDD.n4082 GND 0.00fF
C4592 VDD.n4083 GND 0.00fF
C4593 VDD.n4084 GND 0.00fF
C4594 VDD.n4085 GND 0.00fF
C4595 VDD.n4086 GND 0.00fF
C4596 VDD.n4087 GND 0.00fF
C4597 VDD.n4088 GND 0.00fF
C4598 VDD.n4089 GND 0.00fF
C4599 VDD.n4090 GND 0.00fF
C4600 VDD.n4091 GND 0.00fF
C4601 VDD.n4092 GND 0.00fF
C4602 VDD.n4093 GND 0.00fF
C4603 VDD.n4094 GND 0.00fF
C4604 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/SOURCE GND 0.01fF
C4605 VDD.n4095 GND 0.01fF
C4606 VDD.n4096 GND 0.01fF
C4607 VDD.n4097 GND 0.01fF
C4608 VDD.n4098 GND 0.00fF
C4609 VDD.n4099 GND 0.01fF
C4610 VDD.n4100 GND 0.00fF
C4611 VDD.n4101 GND 0.01fF
C4612 VDD.n4102 GND 0.01fF
C4613 VDD.n4103 GND 0.01fF
C4614 VDD.n4104 GND 0.01fF
C4615 VDD.n4105 GND 0.01fF
C4616 VDD.n4106 GND 0.01fF
C4617 VDD.n4107 GND 0.00fF
C4618 VDD.n4108 GND 0.00fF
C4619 VDD.n4109 GND 0.00fF
C4620 VDD.n4110 GND 0.00fF
C4621 VDD.n4111 GND 0.00fF
C4622 VDD.n4112 GND 0.00fF
C4623 VDD.n4113 GND 0.00fF
C4624 VDD.n4114 GND 0.00fF
C4625 VDD.n4115 GND 0.00fF
C4626 VDD.n4116 GND 0.00fF
C4627 VDD.n4117 GND 0.00fF
C4628 VDD.n4118 GND 0.00fF
C4629 VDD.n4119 GND 0.00fF
C4630 VDD.n4120 GND 0.00fF
C4631 VDD.n4121 GND 0.00fF
C4632 VDD.n4122 GND 0.00fF
C4633 VDD.n4123 GND 0.00fF
C4634 VDD.n4124 GND 0.00fF
C4635 VDD.n4125 GND 0.00fF
C4636 VDD.t65 GND 0.04fF $ **FLOATING
C4637 VDD.n4126 GND 0.13fF
C4638 VDD.n4127 GND 0.00fF
C4639 VDD.n4128 GND 0.04fF
C4640 VDD.n4129 GND 0.07fF
C4641 VDD.n4130 GND 0.00fF
C4642 VDD.n4131 GND 0.00fF
C4643 VDD.n4132 GND 0.00fF
C4644 VDD.n4133 GND 0.00fF
C4645 VDD.n4134 GND 0.00fF
C4646 VDD.n4135 GND 0.00fF
C4647 VDD.n4136 GND 0.00fF
C4648 VDD.n4137 GND 0.00fF
C4649 VDD.n4138 GND 0.00fF
C4650 VDD.n4139 GND 0.00fF
C4651 VDD.n4140 GND 0.00fF
C4652 VDD.n4141 GND 0.00fF
C4653 VDD.n4142 GND 0.00fF
C4654 VDD.n4143 GND 0.00fF
C4655 VDD.n4144 GND 0.00fF
C4656 VDD.n4145 GND 0.00fF
C4657 VDD.n4146 GND 0.00fF
C4658 VDD.n4147 GND 0.02fF
C4659 VDD.n4149 GND 0.02fF
C4660 VDD.n4150 GND 0.01fF
C4661 VDD.n4151 GND 0.01fF
C4662 VDD.n4153 GND 0.01fF
C4663 VDD.n4154 GND 0.01fF
C4664 VDD.n4155 GND 0.01fF
C4665 VDD.n4157 GND 0.01fF
C4666 VDD.n4158 GND 0.01fF
C4667 VDD.n4159 GND 0.01fF
C4668 VDD.n4160 GND 0.01fF
C4669 VDD.n4161 GND 0.01fF
C4670 VDD.n4162 GND 0.01fF
C4671 VDD.n4163 GND 0.01fF
C4672 VDD.n4164 GND 0.01fF
C4673 VDD.n4165 GND 0.01fF
C4674 VDD.n4166 GND 0.00fF
C4675 VDD.n4167 GND 0.00fF
C4676 VDD.n4168 GND 0.00fF
C4677 VDD.n4169 GND 0.00fF
C4678 VDD.n4170 GND 0.00fF
C4679 VDD.n4171 GND 0.00fF
C4680 VDD.n4172 GND 0.00fF
C4681 VDD.n4173 GND 0.00fF
C4682 VDD.n4174 GND 0.00fF
C4683 VDD.n4175 GND 0.00fF
C4684 VDD.n4176 GND 0.00fF
C4685 VDD.n4177 GND 0.00fF
C4686 VDD.n4178 GND 0.00fF
C4687 VDD.n4179 GND 0.00fF
C4688 VDD.n4180 GND 0.00fF
C4689 VDD.n4181 GND 0.00fF
C4690 VDD.n4182 GND 0.00fF
C4691 VDD.n4183 GND 0.00fF
C4692 VDD.n4184 GND 0.00fF
C4693 VDD.t61 GND 0.04fF $ **FLOATING
C4694 VDD.n4185 GND 0.13fF
C4695 VDD.n4186 GND 0.00fF
C4696 VDD.n4187 GND 0.04fF
C4697 VDD.n4188 GND 0.07fF
C4698 VDD.n4189 GND 0.00fF
C4699 VDD.n4190 GND 0.00fF
C4700 VDD.n4191 GND 0.00fF
C4701 VDD.n4192 GND 0.00fF
C4702 VDD.n4193 GND 0.00fF
C4703 VDD.n4194 GND 0.00fF
C4704 VDD.n4195 GND 0.00fF
C4705 VDD.n4196 GND 0.00fF
C4706 VDD.n4197 GND 0.00fF
C4707 VDD.n4198 GND 0.00fF
C4708 VDD.n4199 GND 0.00fF
C4709 VDD.n4200 GND 0.00fF
C4710 VDD.n4201 GND 0.00fF
C4711 VDD.n4202 GND 0.00fF
C4712 VDD.n4203 GND 0.00fF
C4713 VDD.n4204 GND 0.00fF
C4714 VDD.n4205 GND 0.00fF
C4715 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/SOURCE GND 0.01fF
C4716 VDD.n4206 GND 0.01fF
C4717 VDD.n4207 GND 0.01fF
C4718 VDD.n4208 GND 0.01fF
C4719 VDD.n4209 GND 0.00fF
C4720 VDD.n4210 GND 0.01fF
C4721 VDD.n4211 GND 0.00fF
C4722 VDD.n4212 GND 0.01fF
C4723 VDD.n4213 GND 0.01fF
C4724 VDD.n4214 GND 0.01fF
C4725 VDD.n4215 GND 0.01fF
C4726 VDD.n4216 GND 0.01fF
C4727 VDD.n4217 GND 0.01fF
C4728 VDD.n4218 GND 0.00fF
C4729 VDD.n4219 GND 0.00fF
C4730 VDD.n4220 GND 0.00fF
C4731 VDD.n4221 GND 0.00fF
C4732 VDD.n4222 GND 0.00fF
C4733 VDD.n4223 GND 0.00fF
C4734 VDD.n4224 GND 0.00fF
C4735 VDD.n4225 GND 0.00fF
C4736 VDD.n4226 GND 0.00fF
C4737 VDD.n4227 GND 0.00fF
C4738 VDD.n4228 GND 0.00fF
C4739 VDD.n4229 GND 0.00fF
C4740 VDD.n4230 GND 0.00fF
C4741 VDD.n4231 GND 0.00fF
C4742 VDD.n4232 GND 0.00fF
C4743 VDD.n4233 GND 0.00fF
C4744 VDD.n4234 GND 0.00fF
C4745 VDD.n4235 GND 0.00fF
C4746 VDD.n4236 GND 0.00fF
C4747 VDD.t51 GND 0.04fF $ **FLOATING
C4748 VDD.n4237 GND 0.13fF
C4749 VDD.n4238 GND 0.00fF
C4750 VDD.n4239 GND 0.04fF
C4751 VDD.n4240 GND 0.07fF
C4752 VDD.n4241 GND 0.00fF
C4753 VDD.n4242 GND 0.00fF
C4754 VDD.n4243 GND 0.00fF
C4755 VDD.n4244 GND 0.00fF
C4756 VDD.n4245 GND 0.00fF
C4757 VDD.n4246 GND 0.00fF
C4758 VDD.n4247 GND 0.00fF
C4759 VDD.n4248 GND 0.00fF
C4760 VDD.n4249 GND 0.00fF
C4761 VDD.n4250 GND 0.00fF
C4762 VDD.n4251 GND 0.00fF
C4763 VDD.n4252 GND 0.00fF
C4764 VDD.n4253 GND 0.00fF
C4765 VDD.n4254 GND 0.00fF
C4766 VDD.n4255 GND 0.00fF
C4767 VDD.n4256 GND 0.00fF
C4768 VDD.n4257 GND 0.00fF
C4769 VDD.n4258 GND 0.02fF
C4770 VDD.n4260 GND 0.05fF
C4771 VDD.n4262 GND 0.04fF
C4772 VDD.n4263 GND 0.06fF
C4773 VDD.n4264 GND 0.04fF
C4774 VDD.n4266 GND 0.14fF
C4775 VDD.n4267 GND 0.14fF
C4776 VDD.n4269 GND 0.04fF
C4777 VDD.n4270 GND 0.06fF
C4778 VDD.n4271 GND 0.04fF
C4779 VDD.n4273 GND 0.14fF
C4780 VDD.n4274 GND 0.14fF
C4781 VDD.n4276 GND 0.04fF
C4782 VDD.n4277 GND 0.06fF
C4783 VDD.n4278 GND 0.04fF
C4784 VDD.n4280 GND 0.14fF
C4785 VDD.n4281 GND 0.14fF
C4786 VDD.n4283 GND 0.04fF
C4787 VDD.n4284 GND 0.06fF
C4788 VDD.n4285 GND 0.04fF
C4789 VDD.n4287 GND 0.14fF
C4790 VDD.n4288 GND 0.14fF
C4791 VDD.n4290 GND 0.04fF
C4792 VDD.n4291 GND 0.06fF
C4793 VDD.n4292 GND 0.04fF
C4794 VDD.n4294 GND 0.14fF
C4795 VDD.n4295 GND 0.16fF
C4796 VDD.n4297 GND 0.46fF
C4797 VDD.n4298 GND 0.46fF
C4798 VDD.n4300 GND 0.16fF
C4799 VDD.n4301 GND 0.14fF
C4800 VDD.n4303 GND 0.04fF
C4801 VDD.n4304 GND 0.06fF
C4802 VDD.n4305 GND 0.04fF
C4803 VDD.n4307 GND 0.02fF
C4804 VDD.n4308 GND 0.01fF
C4805 VDD.n4309 GND 0.01fF
C4806 VDD.n4311 GND 0.01fF
C4807 VDD.n4312 GND 0.01fF
C4808 VDD.n4313 GND 0.01fF
C4809 VDD.n4315 GND 0.01fF
C4810 VDD.n4316 GND 0.01fF
C4811 VDD.n4317 GND 0.01fF
C4812 VDD.n4318 GND 0.01fF
C4813 VDD.n4319 GND 0.01fF
C4814 VDD.n4320 GND 0.01fF
C4815 VDD.n4321 GND 0.01fF
C4816 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/SOURCE GND 0.01fF
C4817 VDD.n4322 GND 0.01fF
C4818 VDD.n4323 GND 0.01fF
C4819 VDD.n4324 GND 0.01fF
C4820 VDD.n4325 GND 0.00fF
C4821 VDD.n4326 GND 0.01fF
C4822 VDD.n4327 GND 0.00fF
C4823 VDD.n4328 GND 0.01fF
C4824 VDD.n4329 GND 0.01fF
C4825 VDD.n4330 GND 0.01fF
C4826 VDD.n4331 GND 0.01fF
C4827 VDD.n4332 GND 0.01fF
C4828 VDD.n4333 GND 0.01fF
C4829 VDD.n4334 GND 0.00fF
C4830 VDD.n4335 GND 0.00fF
C4831 VDD.n4336 GND 0.00fF
C4832 VDD.n4337 GND 0.00fF
C4833 VDD.n4338 GND 0.00fF
C4834 VDD.n4339 GND 0.00fF
C4835 VDD.n4340 GND 0.00fF
C4836 VDD.n4341 GND 0.00fF
C4837 VDD.n4342 GND 0.00fF
C4838 VDD.n4343 GND 0.00fF
C4839 VDD.n4344 GND 0.00fF
C4840 VDD.n4345 GND 0.00fF
C4841 VDD.n4346 GND 0.00fF
C4842 VDD.n4347 GND 0.00fF
C4843 VDD.n4348 GND 0.00fF
C4844 VDD.n4349 GND 0.00fF
C4845 VDD.n4350 GND 0.00fF
C4846 VDD.n4351 GND 0.00fF
C4847 VDD.n4352 GND 0.00fF
C4848 VDD.t58 GND 0.04fF $ **FLOATING
C4849 VDD.n4353 GND 0.13fF
C4850 VDD.n4354 GND 0.00fF
C4851 VDD.n4355 GND 0.04fF
C4852 VDD.n4356 GND 0.07fF
C4853 VDD.n4357 GND 0.00fF
C4854 VDD.n4358 GND 0.00fF
C4855 VDD.n4359 GND 0.00fF
C4856 VDD.n4360 GND 0.00fF
C4857 VDD.n4361 GND 0.00fF
C4858 VDD.n4362 GND 0.00fF
C4859 VDD.n4363 GND 0.00fF
C4860 VDD.n4364 GND 0.00fF
C4861 VDD.n4365 GND 0.00fF
C4862 VDD.n4366 GND 0.00fF
C4863 VDD.n4367 GND 0.00fF
C4864 VDD.n4368 GND 0.00fF
C4865 VDD.n4369 GND 0.00fF
C4866 VDD.n4370 GND 0.00fF
C4867 VDD.n4371 GND 0.00fF
C4868 VDD.n4372 GND 0.00fF
C4869 VDD.n4373 GND 0.00fF
C4870 VDD.n4374 GND 0.01fF
C4871 VDD.n4375 GND 0.01fF
C4872 VDD.n4376 GND 0.00fF
C4873 VDD.n4377 GND 0.00fF
C4874 VDD.n4378 GND 0.00fF
C4875 VDD.n4379 GND 0.00fF
C4876 VDD.n4380 GND 0.00fF
C4877 VDD.n4381 GND 0.00fF
C4878 VDD.n4382 GND 0.00fF
C4879 VDD.n4383 GND 0.00fF
C4880 VDD.n4384 GND 0.00fF
C4881 VDD.n4385 GND 0.00fF
C4882 VDD.n4386 GND 0.00fF
C4883 VDD.n4387 GND 0.00fF
C4884 VDD.n4388 GND 0.00fF
C4885 VDD.n4389 GND 0.00fF
C4886 VDD.n4390 GND 0.00fF
C4887 VDD.n4391 GND 0.00fF
C4888 VDD.n4392 GND 0.00fF
C4889 VDD.n4393 GND 0.00fF
C4890 VDD.n4394 GND 0.00fF
C4891 VDD.t62 GND 0.04fF $ **FLOATING
C4892 VDD.n4395 GND 0.13fF
C4893 VDD.n4396 GND 0.00fF
C4894 VDD.n4397 GND 0.04fF
C4895 VDD.n4398 GND 0.07fF
C4896 VDD.n4399 GND 0.00fF
C4897 VDD.n4400 GND 0.00fF
C4898 VDD.n4401 GND 0.00fF
C4899 VDD.n4402 GND 0.00fF
C4900 VDD.n4403 GND 0.00fF
C4901 VDD.n4404 GND 0.00fF
C4902 VDD.n4405 GND 0.00fF
C4903 VDD.n4406 GND 0.00fF
C4904 VDD.n4407 GND 0.00fF
C4905 VDD.n4408 GND 0.00fF
C4906 VDD.n4409 GND 0.00fF
C4907 VDD.n4410 GND 0.00fF
C4908 VDD.n4411 GND 0.00fF
C4909 VDD.n4412 GND 0.00fF
C4910 VDD.n4413 GND 0.00fF
C4911 VDD.n4414 GND 0.00fF
C4912 VDD.n4415 GND 0.00fF
C4913 VDD.n4416 GND 0.02fF
C4914 VDD.n4418 GND 0.14fF
C4915 VDD.n4419 GND 0.14fF
C4916 VDD.n4421 GND 0.04fF
C4917 VDD.n4422 GND 0.06fF
C4918 VDD.n4423 GND 0.04fF
C4919 VDD.n4425 GND 0.02fF
C4920 VDD.n4426 GND 0.01fF
C4921 VDD.n4427 GND 0.01fF
C4922 VDD.n4429 GND 0.01fF
C4923 VDD.n4430 GND 0.01fF
C4924 VDD.n4431 GND 0.01fF
C4925 VDD.n4433 GND 0.01fF
C4926 VDD.n4434 GND 0.01fF
C4927 VDD.n4435 GND 0.01fF
C4928 VDD.n4436 GND 0.01fF
C4929 VDD.n4437 GND 0.01fF
C4930 VDD.n4438 GND 0.01fF
C4931 VDD.n4439 GND 0.01fF
C4932 VDD.n4440 GND 0.01fF
C4933 VDD.n4441 GND 0.01fF
C4934 VDD.n4442 GND 0.00fF
C4935 VDD.n4443 GND 0.00fF
C4936 VDD.n4444 GND 0.00fF
C4937 VDD.n4445 GND 0.00fF
C4938 VDD.n4446 GND 0.00fF
C4939 VDD.n4447 GND 0.00fF
C4940 VDD.n4448 GND 0.00fF
C4941 VDD.n4449 GND 0.00fF
C4942 VDD.n4450 GND 0.00fF
C4943 VDD.n4451 GND 0.00fF
C4944 VDD.n4452 GND 0.00fF
C4945 VDD.n4453 GND 0.00fF
C4946 VDD.n4454 GND 0.00fF
C4947 VDD.n4455 GND 0.00fF
C4948 VDD.n4456 GND 0.00fF
C4949 VDD.n4457 GND 0.00fF
C4950 VDD.n4458 GND 0.00fF
C4951 VDD.n4459 GND 0.00fF
C4952 VDD.n4460 GND 0.00fF
C4953 VDD.t42 GND 0.04fF $ **FLOATING
C4954 VDD.n4461 GND 0.13fF
C4955 VDD.n4462 GND 0.00fF
C4956 VDD.n4463 GND 0.04fF
C4957 VDD.n4464 GND 0.07fF
C4958 VDD.n4465 GND 0.00fF
C4959 VDD.n4466 GND 0.00fF
C4960 VDD.n4467 GND 0.00fF
C4961 VDD.n4468 GND 0.00fF
C4962 VDD.n4469 GND 0.00fF
C4963 VDD.n4470 GND 0.00fF
C4964 VDD.n4471 GND 0.00fF
C4965 VDD.n4472 GND 0.00fF
C4966 VDD.n4473 GND 0.00fF
C4967 VDD.n4474 GND 0.00fF
C4968 VDD.n4475 GND 0.00fF
C4969 VDD.n4476 GND 0.00fF
C4970 VDD.n4477 GND 0.00fF
C4971 VDD.n4478 GND 0.00fF
C4972 VDD.n4479 GND 0.00fF
C4973 VDD.n4480 GND 0.00fF
C4974 VDD.n4481 GND 0.00fF
C4975 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/SOURCE GND 0.01fF
C4976 VDD.n4482 GND 0.01fF
C4977 VDD.n4483 GND 0.01fF
C4978 VDD.n4484 GND 0.01fF
C4979 VDD.n4485 GND 0.00fF
C4980 VDD.n4486 GND 0.01fF
C4981 VDD.n4487 GND 0.00fF
C4982 VDD.n4488 GND 0.01fF
C4983 VDD.n4489 GND 0.01fF
C4984 VDD.n4490 GND 0.01fF
C4985 VDD.n4491 GND 0.01fF
C4986 VDD.n4492 GND 0.01fF
C4987 VDD.n4493 GND 0.01fF
C4988 VDD.n4494 GND 0.00fF
C4989 VDD.n4495 GND 0.00fF
C4990 VDD.n4496 GND 0.00fF
C4991 VDD.n4497 GND 0.00fF
C4992 VDD.n4498 GND 0.00fF
C4993 VDD.n4499 GND 0.00fF
C4994 VDD.n4500 GND 0.00fF
C4995 VDD.n4501 GND 0.00fF
C4996 VDD.n4502 GND 0.00fF
C4997 VDD.n4503 GND 0.00fF
C4998 VDD.n4504 GND 0.00fF
C4999 VDD.n4505 GND 0.00fF
C5000 VDD.n4506 GND 0.00fF
C5001 VDD.n4507 GND 0.00fF
C5002 VDD.n4508 GND 0.00fF
C5003 VDD.n4509 GND 0.00fF
C5004 VDD.n4510 GND 0.00fF
C5005 VDD.n4511 GND 0.00fF
C5006 VDD.n4512 GND 0.00fF
C5007 VDD.t49 GND 0.04fF $ **FLOATING
C5008 VDD.n4513 GND 0.13fF
C5009 VDD.n4514 GND 0.00fF
C5010 VDD.n4515 GND 0.04fF
C5011 VDD.n4516 GND 0.07fF
C5012 VDD.n4517 GND 0.00fF
C5013 VDD.n4518 GND 0.00fF
C5014 VDD.n4519 GND 0.00fF
C5015 VDD.n4520 GND 0.00fF
C5016 VDD.n4521 GND 0.00fF
C5017 VDD.n4522 GND 0.00fF
C5018 VDD.n4523 GND 0.00fF
C5019 VDD.n4524 GND 0.00fF
C5020 VDD.n4525 GND 0.00fF
C5021 VDD.n4526 GND 0.00fF
C5022 VDD.n4527 GND 0.00fF
C5023 VDD.n4528 GND 0.00fF
C5024 VDD.n4529 GND 0.00fF
C5025 VDD.n4530 GND 0.00fF
C5026 VDD.n4531 GND 0.00fF
C5027 VDD.n4532 GND 0.00fF
C5028 VDD.n4533 GND 0.00fF
C5029 VDD.n4534 GND 0.02fF
C5030 VDD.n4536 GND 0.35fF
C5031 VDD.n4537 GND 0.35fF
C5032 VDD.n4539 GND 0.04fF
C5033 VDD.n4540 GND 0.06fF
C5034 VDD.n4541 GND 0.04fF
C5035 VDD.n4543 GND 0.02fF
C5036 VDD.n4544 GND 0.01fF
C5037 VDD.n4545 GND 0.01fF
C5038 VDD.n4547 GND 0.01fF
C5039 VDD.n4548 GND 0.01fF
C5040 VDD.n4549 GND 0.01fF
C5041 VDD.n4551 GND 0.01fF
C5042 VDD.n4552 GND 0.01fF
C5043 VDD.n4553 GND 0.01fF
C5044 VDD.n4554 GND 0.01fF
C5045 VDD.n4555 GND 0.01fF
C5046 VDD.n4556 GND 0.01fF
C5047 VDD.n4557 GND 0.01fF
C5048 VDD.n4558 GND 0.01fF
C5049 VDD.n4559 GND 0.01fF
C5050 VDD.n4560 GND 0.00fF
C5051 VDD.n4561 GND 0.00fF
C5052 VDD.n4562 GND 0.00fF
C5053 VDD.n4563 GND 0.00fF
C5054 VDD.n4564 GND 0.00fF
C5055 VDD.n4565 GND 0.00fF
C5056 VDD.n4566 GND 0.00fF
C5057 VDD.n4567 GND 0.00fF
C5058 VDD.n4568 GND 0.00fF
C5059 VDD.n4569 GND 0.00fF
C5060 VDD.n4570 GND 0.00fF
C5061 VDD.n4571 GND 0.00fF
C5062 VDD.n4572 GND 0.00fF
C5063 VDD.n4573 GND 0.00fF
C5064 VDD.n4574 GND 0.00fF
C5065 VDD.n4575 GND 0.00fF
C5066 VDD.n4576 GND 0.00fF
C5067 VDD.n4577 GND 0.00fF
C5068 VDD.n4578 GND 0.00fF
C5069 VDD.t45 GND 0.04fF $ **FLOATING
C5070 VDD.n4579 GND 0.13fF
C5071 VDD.n4580 GND 0.00fF
C5072 VDD.n4581 GND 0.04fF
C5073 VDD.n4582 GND 0.07fF
C5074 VDD.n4583 GND 0.00fF
C5075 VDD.n4584 GND 0.00fF
C5076 VDD.n4585 GND 0.00fF
C5077 VDD.n4586 GND 0.00fF
C5078 VDD.n4587 GND 0.00fF
C5079 VDD.n4588 GND 0.00fF
C5080 VDD.n4589 GND 0.00fF
C5081 VDD.n4590 GND 0.00fF
C5082 VDD.n4591 GND 0.00fF
C5083 VDD.n4592 GND 0.00fF
C5084 VDD.n4593 GND 0.00fF
C5085 VDD.n4594 GND 0.00fF
C5086 VDD.n4595 GND 0.00fF
C5087 VDD.n4596 GND 0.00fF
C5088 VDD.n4597 GND 0.00fF
C5089 VDD.n4598 GND 0.00fF
C5090 VDD.n4599 GND 0.00fF
C5091 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/SOURCE GND 0.01fF
C5092 VDD.n4600 GND 0.01fF
C5093 VDD.n4601 GND 0.01fF
C5094 VDD.n4602 GND 0.01fF
C5095 VDD.n4603 GND 0.00fF
C5096 VDD.n4604 GND 0.01fF
C5097 VDD.n4605 GND 0.00fF
C5098 VDD.n4606 GND 0.01fF
C5099 VDD.n4607 GND 0.01fF
C5100 VDD.n4608 GND 0.01fF
C5101 VDD.n4609 GND 0.01fF
C5102 VDD.n4610 GND 0.01fF
C5103 VDD.n4611 GND 0.01fF
C5104 VDD.n4612 GND 0.00fF
C5105 VDD.n4613 GND 0.00fF
C5106 VDD.n4614 GND 0.00fF
C5107 VDD.n4615 GND 0.00fF
C5108 VDD.n4616 GND 0.00fF
C5109 VDD.n4617 GND 0.00fF
C5110 VDD.n4618 GND 0.00fF
C5111 VDD.n4619 GND 0.00fF
C5112 VDD.n4620 GND 0.00fF
C5113 VDD.n4621 GND 0.00fF
C5114 VDD.n4622 GND 0.00fF
C5115 VDD.n4623 GND 0.00fF
C5116 VDD.n4624 GND 0.00fF
C5117 VDD.n4625 GND 0.00fF
C5118 VDD.n4626 GND 0.00fF
C5119 VDD.n4627 GND 0.00fF
C5120 VDD.n4628 GND 0.00fF
C5121 VDD.n4629 GND 0.00fF
C5122 VDD.n4630 GND 0.00fF
C5123 VDD.t54 GND 0.04fF $ **FLOATING
C5124 VDD.n4631 GND 0.13fF
C5125 VDD.n4632 GND 0.00fF
C5126 VDD.n4633 GND 0.04fF
C5127 VDD.n4634 GND 0.07fF
C5128 VDD.n4635 GND 0.00fF
C5129 VDD.n4636 GND 0.00fF
C5130 VDD.n4637 GND 0.00fF
C5131 VDD.n4638 GND 0.00fF
C5132 VDD.n4639 GND 0.00fF
C5133 VDD.n4640 GND 0.00fF
C5134 VDD.n4641 GND 0.00fF
C5135 VDD.n4642 GND 0.00fF
C5136 VDD.n4643 GND 0.00fF
C5137 VDD.n4644 GND 0.00fF
C5138 VDD.n4645 GND 0.00fF
C5139 VDD.n4646 GND 0.00fF
C5140 VDD.n4647 GND 0.00fF
C5141 VDD.n4648 GND 0.00fF
C5142 VDD.n4649 GND 0.00fF
C5143 VDD.n4650 GND 0.00fF
C5144 VDD.n4651 GND 0.00fF
C5145 VDD.n4652 GND 0.02fF
C5146 VDD.n4654 GND 0.14fF
C5147 VDD.n4655 GND 0.14fF
C5148 VDD.n4657 GND 0.04fF
C5149 VDD.n4658 GND 0.06fF
C5150 VDD.n4659 GND 0.04fF
C5151 VDD.n4661 GND 0.05fF
C5152 VDD.n4663 GND 0.01fF
C5153 VDD.n4664 GND 0.01fF
C5154 VDD.n4665 GND 0.00fF
C5155 VDD.n4666 GND 0.00fF
C5156 VDD.n4667 GND 0.00fF
C5157 VDD.n4668 GND 0.00fF
C5158 VDD.n4669 GND 0.00fF
C5159 VDD.n4670 GND 0.00fF
C5160 VDD.n4671 GND 0.00fF
C5161 VDD.n4672 GND 0.00fF
C5162 VDD.n4673 GND 0.00fF
C5163 VDD.n4674 GND 0.00fF
C5164 VDD.n4675 GND 0.00fF
C5165 VDD.n4676 GND 0.00fF
C5166 VDD.n4677 GND 0.00fF
C5167 VDD.n4678 GND 0.00fF
C5168 VDD.n4679 GND 0.00fF
C5169 VDD.n4680 GND 0.00fF
C5170 VDD.n4681 GND 0.00fF
C5171 VDD.n4682 GND 0.00fF
C5172 VDD.n4683 GND 0.00fF
C5173 VDD.t57 GND 0.04fF $ **FLOATING
C5174 VDD.n4684 GND 0.13fF
C5175 VDD.n4685 GND 0.00fF
C5176 VDD.n4686 GND 0.04fF
C5177 VDD.n4687 GND 0.07fF
C5178 VDD.n4688 GND 0.00fF
C5179 VDD.n4689 GND 0.00fF
C5180 VDD.n4690 GND 0.00fF
C5181 VDD.n4691 GND 0.00fF
C5182 VDD.n4692 GND 0.00fF
C5183 VDD.n4693 GND 0.00fF
C5184 VDD.n4694 GND 0.00fF
C5185 VDD.n4695 GND 0.00fF
C5186 VDD.n4696 GND 0.00fF
C5187 VDD.n4697 GND 0.00fF
C5188 VDD.n4698 GND 0.00fF
C5189 VDD.n4699 GND 0.00fF
C5190 VDD.n4700 GND 0.00fF
C5191 VDD.n4701 GND 0.00fF
C5192 VDD.n4702 GND 0.00fF
C5193 VDD.n4703 GND 0.00fF
C5194 VDD.n4704 GND 0.00fF
C5195 VDD.n4705 GND 0.02fF
C5196 VDD.n4706 GND 0.01fF
C5197 VDD.n4707 GND 0.01fF
C5198 VDD.n4708 GND 0.01fF
C5199 VDD.n4709 GND 0.01fF
C5200 VDD.n4710 GND 0.00fF
C5201 VDD.n4711 GND 0.01fF
C5202 VDD.n4712 GND 0.00fF
C5203 VDD.n4713 GND 0.01fF
C5204 VDD.n4714 GND 0.01fF
C5205 VDD.n4715 GND 0.01fF
C5206 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/SOURCE GND 0.01fF
C5207 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n0 GND 0.01fF
C5208 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1 GND 0.00fF
C5209 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n2 GND 0.00fF
C5210 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t2 GND 0.08fF $ **FLOATING
C5211 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t4 GND 0.08fF $ **FLOATING
C5212 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n3 GND 0.21fF
C5213 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n4 GND 0.00fF
C5214 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n5 GND 0.01fF
C5215 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n6 GND 0.09fF
C5216 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n7 GND 0.14fF
C5217 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n8 GND 0.08fF
C5218 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n9 GND 0.06fF
C5219 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n10 GND 0.01fF
C5220 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n11 GND 0.01fF
C5221 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n12 GND 0.00fF
C5222 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n13 GND 0.00fF
C5223 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n14 GND 0.01fF
C5224 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n15 GND 0.01fF
C5225 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n16 GND 0.00fF
C5226 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n17 GND 0.00fF
C5227 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n18 GND 0.00fF
C5228 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n19 GND 0.00fF
C5229 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n20 GND 0.00fF
C5230 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n21 GND 0.06fF
C5231 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n22 GND 0.03fF
C5232 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n23 GND 0.05fF
C5233 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n24 GND 0.05fF
C5234 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n25 GND 0.01fF
C5235 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n26 GND 0.01fF
C5236 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n27 GND 0.00fF
C5237 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n28 GND 0.01fF
C5238 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n29 GND 0.01fF
C5239 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n30 GND 0.00fF
C5240 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n31 GND 0.00fF
C5241 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n32 GND 0.00fF
C5242 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n33 GND 0.00fF
C5243 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n34 GND 0.00fF
C5244 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n35 GND 0.03fF
C5245 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n36 GND 0.03fF
C5246 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n37 GND 0.05fF
C5247 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n38 GND 0.05fF
C5248 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n39 GND 0.03fF
C5249 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n40 GND 0.01fF
C5250 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n41 GND 0.01fF
C5251 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n42 GND 0.01fF
C5252 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n43 GND 0.00fF
C5253 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n44 GND 0.02fF
C5254 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n45 GND 0.01fF
C5255 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n46 GND 0.00fF
C5256 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n47 GND 0.00fF
C5257 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n48 GND 0.03fF
C5258 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n49 GND 0.03fF
C5259 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n50 GND 0.01fF
C5260 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n51 GND 0.01fF
C5261 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/GATE GND 0.02fF
C5262 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n52 GND 0.01fF
C5263 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n53 GND 0.00fF
C5264 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t3 GND 0.10fF $ **FLOATING
C5265 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n54 GND 0.07fF
C5266 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n55 GND 0.02fF
C5267 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n56 GND 0.02fF
C5268 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n57 GND 0.01fF
C5269 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n58 GND 0.01fF
C5270 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n59 GND 0.01fF
C5271 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n60 GND 0.00fF
C5272 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n61 GND 0.03fF
C5273 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n62 GND 0.01fF
C5274 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n63 GND 0.01fF
C5275 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n64 GND 0.01fF
C5276 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n65 GND 0.01fF
C5277 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n66 GND 0.00fF
C5278 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t1 GND 0.10fF $ **FLOATING
C5279 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n67 GND 0.08fF
C5280 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n68 GND 0.03fF
C5281 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n69 GND 0.05fF
C5282 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n70 GND 0.01fF
C5283 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n71 GND 0.07fF
C5284 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n72 GND 0.26fF
C5285 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n73 GND 0.10fF
C5286 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n74 GND 0.07fF
C5287 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n75 GND 0.05fF
C5288 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n76 GND 0.05fF
C5289 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n77 GND 0.04fF
C5290 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n78 GND 0.40fF
C5291 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t0 GND 0.61fF $ **FLOATING
C5292 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n79 GND 6.53fF
C5293 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n80 GND 2.07fF
C5294 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n81 GND 0.05fF
C5295 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n82 GND 0.05fF
C5296 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n83 GND 0.10fF
C5297 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n84 GND 0.12fF
C5298 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n85 GND 0.08fF
C5299 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n86 GND 0.15fF
C5300 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n87 GND 0.08fF
C5301 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n88 GND 0.06fF
C5302 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n89 GND 0.85fF
C5303 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n90 GND 0.79fF
C5304 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n91 GND 0.03fF
C5305 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n92 GND 0.01fF
C5306 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n93 GND 0.00fF
C5307 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_1/GATE GND 0.02fF
C5308 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n94 GND 0.07fF
C5309 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n95 GND 0.02fF
C5310 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n96 GND 0.01fF
C5311 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n97 GND 0.00fF
C5312 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n98 GND 0.02fF
C5313 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n99 GND 0.01fF
C5314 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n100 GND 0.01fF
C5315 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n101 GND 0.01fF
C5316 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n102 GND 0.00fF
C5317 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n103 GND 0.00fF
C5318 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n104 GND 0.01fF
C5319 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n105 GND 0.01fF
C5320 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n106 GND 0.01fF
C5321 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n107 GND 0.01fF
C5322 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n108 GND 0.01fF
C5323 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n109 GND 0.01fF
C5324 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n110 GND 0.00fF
C5325 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n111 GND 0.00fF
C5326 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n112 GND 0.01fF
C5327 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n113 GND 0.00fF
C5328 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n114 GND 0.07fF
C5329 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n115 GND 0.02fF
C5330 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n116 GND 0.02fF
C5331 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n117 GND 0.03fF
C5332 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n118 GND 0.01fF
C5333 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n119 GND 0.01fF
C5334 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n120 GND 0.01fF
C5335 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n121 GND 0.01fF
C5336 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n122 GND 0.01fF
C5337 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n123 GND 0.03fF
C5338 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n124 GND 0.01fF
C5339 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n125 GND 0.01fF
C5340 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n126 GND 0.01fF
C5341 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n127 GND 0.01fF
C5342 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n128 GND 0.01fF
C5343 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n129 GND 0.00fF
C5344 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n130 GND 0.01fF
C5345 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n131 GND 0.01fF
C5346 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n132 GND 0.01fF
C5347 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n133 GND 0.04fF
C5348 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n134 GND 0.00fF
C5349 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n135 GND 0.01fF
C5350 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n136 GND 0.01fF
C5351 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n137 GND 0.01fF
C5352 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n138 GND 0.01fF
C5353 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n139 GND 0.00fF
C5354 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n140 GND 0.00fF
C5355 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n141 GND 0.00fF
C5356 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n142 GND 0.00fF
C5357 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n143 GND 0.03fF
C5358 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n144 GND 0.01fF
C5359 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n146 GND 0.02fF
C5360 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n147 GND 0.01fF
C5361 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n148 GND 0.01fF
C5362 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n149 GND 0.00fF
C5363 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n150 GND 0.00fF
C5364 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n151 GND 0.00fF
C5365 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n152 GND 0.01fF
C5366 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n153 GND 0.08fF
C5367 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n154 GND 0.03fF
C5368 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n155 GND 0.04fF
C5369 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n156 GND 0.01fF
C5370 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n157 GND 0.00fF
C5371 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n158 GND 0.00fF
C5372 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n159 GND 0.00fF
C5373 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n160 GND 0.00fF
C5374 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n161 GND 0.01fF
C5375 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n162 GND 0.01fF
C5376 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n163 GND 0.01fF
C5377 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n164 GND 0.00fF
C5378 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n165 GND 0.00fF
C5379 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n166 GND 0.03fF
C5380 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n167 GND 0.00fF
C5381 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n168 GND 0.01fF
C5382 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n169 GND 0.01fF
C5383 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n170 GND 0.01fF
C5384 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_2/GATE GND 0.01fF
C5385 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n171 GND 0.07fF
C5386 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n172 GND 0.02fF
C5387 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n173 GND 0.01fF
C5388 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n174 GND 0.00fF
C5389 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n175 GND 0.02fF
C5390 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n176 GND 0.01fF
C5391 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n177 GND 0.01fF
C5392 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n178 GND 0.01fF
C5393 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n179 GND 0.01fF
C5394 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n180 GND 0.00fF
C5395 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n181 GND 0.00fF
C5396 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n182 GND 0.00fF
C5397 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n183 GND 0.01fF
C5398 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n184 GND 0.01fF
C5399 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n186 GND 0.00fF
C5400 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n187 GND 0.01fF
C5401 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n188 GND 0.01fF
C5402 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n189 GND 0.01fF
C5403 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n190 GND 0.01fF
C5404 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n191 GND 0.00fF
C5405 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n192 GND 0.00fF
C5406 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n193 GND 0.00fF
C5407 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n194 GND 0.00fF
C5408 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n195 GND 0.03fF
C5409 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n196 GND 0.01fF
C5410 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n198 GND 0.02fF
C5411 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n199 GND 0.01fF
C5412 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n200 GND 0.01fF
C5413 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n201 GND 0.00fF
C5414 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n202 GND 0.00fF
C5415 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n203 GND 0.00fF
C5416 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n204 GND 0.01fF
C5417 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n205 GND 0.08fF
C5418 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n206 GND 0.03fF
C5419 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n207 GND 0.04fF
C5420 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n208 GND 0.01fF
C5421 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n209 GND 0.00fF
C5422 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n210 GND 0.00fF
C5423 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n211 GND 0.00fF
C5424 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n212 GND 0.00fF
C5425 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n213 GND 0.01fF
C5426 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n214 GND 0.01fF
C5427 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n215 GND 0.01fF
C5428 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n216 GND 0.00fF
C5429 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n217 GND 0.00fF
C5430 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n218 GND 0.03fF
C5431 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n219 GND 0.00fF
C5432 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n220 GND 0.01fF
C5433 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n221 GND 0.01fF
C5434 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n222 GND 0.01fF
C5435 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_4/GATE GND 0.01fF
C5436 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n223 GND 0.07fF
C5437 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n224 GND 0.02fF
C5438 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n225 GND 0.01fF
C5439 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n226 GND 0.00fF
C5440 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n227 GND 0.02fF
C5441 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n228 GND 0.01fF
C5442 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n229 GND 0.01fF
C5443 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n230 GND 0.01fF
C5444 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n231 GND 0.01fF
C5445 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n232 GND 0.00fF
C5446 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n233 GND 0.00fF
C5447 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n234 GND 0.00fF
C5448 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n235 GND 0.01fF
C5449 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n236 GND 0.01fF
C5450 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n238 GND 0.00fF
C5451 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n239 GND 0.01fF
C5452 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n240 GND 0.01fF
C5453 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n241 GND 0.01fF
C5454 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n242 GND 0.01fF
C5455 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n243 GND 0.00fF
C5456 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n244 GND 0.00fF
C5457 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n245 GND 0.00fF
C5458 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n246 GND 0.00fF
C5459 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n247 GND 0.03fF
C5460 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n248 GND 0.01fF
C5461 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n250 GND 0.02fF
C5462 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n251 GND 0.01fF
C5463 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n252 GND 0.01fF
C5464 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n253 GND 0.00fF
C5465 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n254 GND 0.00fF
C5466 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n255 GND 0.00fF
C5467 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n256 GND 0.01fF
C5468 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n257 GND 0.08fF
C5469 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n258 GND 0.03fF
C5470 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n259 GND 0.04fF
C5471 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n260 GND 0.01fF
C5472 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n261 GND 0.00fF
C5473 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n262 GND 0.00fF
C5474 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n263 GND 0.00fF
C5475 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n264 GND 0.00fF
C5476 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n265 GND 0.01fF
C5477 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n266 GND 0.01fF
C5478 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n267 GND 0.01fF
C5479 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n268 GND 0.00fF
C5480 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n269 GND 0.00fF
C5481 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n270 GND 0.03fF
C5482 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n271 GND 0.00fF
C5483 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n272 GND 0.01fF
C5484 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n273 GND 0.01fF
C5485 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n274 GND 0.01fF
C5486 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n275 GND 0.01fF
C5487 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n276 GND 0.00fF
C5488 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n277 GND 0.07fF
C5489 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n278 GND 0.02fF
C5490 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n279 GND 0.02fF
C5491 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n280 GND 0.01fF
C5492 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n281 GND 0.01fF
C5493 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n282 GND 0.01fF
C5494 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n283 GND 0.01fF
C5495 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n284 GND 0.00fF
C5496 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n285 GND 0.00fF
C5497 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n286 GND 0.00fF
C5498 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n287 GND 0.01fF
C5499 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n288 GND 0.01fF
C5500 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n290 GND 0.04fF
C5501 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n291 GND 0.01fF
C5502 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n292 GND 0.01fF
C5503 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n293 GND 0.01fF
C5504 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n294 GND 0.02fF
C5505 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n295 GND 0.01fF
C5506 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n296 GND 0.01fF
C5507 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n297 GND 0.10fF
C5508 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n298 GND 0.10fF
C5509 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n299 GND 0.01fF
C5510 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n300 GND 0.01fF
C5511 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n301 GND 0.01fF
C5512 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n302 GND 0.01fF
C5513 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n303 GND 0.02fF
C5514 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n304 GND 0.01fF
C5515 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n305 GND 0.01fF
C5516 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n306 GND 0.23fF
C5517 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n307 GND 0.23fF
C5518 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n308 GND 0.01fF
C5519 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n309 GND 0.01fF
C5520 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n310 GND 0.01fF
C5521 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n311 GND 0.01fF
C5522 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n312 GND 0.02fF
C5523 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n313 GND 0.01fF
C5524 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n314 GND 0.01fF
C5525 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n315 GND 0.09fF
C5526 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n316 GND 0.09fF
C5527 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n317 GND 0.01fF
C5528 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n318 GND 0.02fF
C5529 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n319 GND 0.03fF
C5530 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n320 GND 0.01fF
C5531 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n321 GND 0.13fF
C5532 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n322 GND 0.30fF
C5533 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n323 GND 0.03fF
C5534 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n324 GND 0.01fF
C5535 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n325 GND 0.00fF
C5536 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n326 GND 0.01fF
C5537 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n327 GND 0.00fF
C5538 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t9 GND 0.10fF $ **FLOATING
C5539 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n328 GND 0.07fF
C5540 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n329 GND 0.02fF
C5541 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n330 GND 0.02fF
C5542 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n331 GND 0.01fF
C5543 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n332 GND 0.01fF
C5544 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n333 GND 0.01fF
C5545 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n334 GND 0.00fF
C5546 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n335 GND 0.00fF
C5547 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n336 GND 0.01fF
C5548 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n337 GND 0.01fF
C5549 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n338 GND 0.01fF
C5550 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n339 GND 0.01fF
C5551 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n340 GND 0.01fF
C5552 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n341 GND 0.01fF
C5553 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n342 GND 0.00fF
C5554 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n343 GND 0.00fF
C5555 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n344 GND 0.01fF
C5556 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n345 GND 0.00fF
C5557 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t11 GND 0.10fF $ **FLOATING
C5558 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n346 GND 0.07fF
C5559 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n347 GND 0.02fF
C5560 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n348 GND 0.02fF
C5561 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n349 GND 0.03fF
C5562 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n350 GND 0.01fF
C5563 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n351 GND 0.03fF
C5564 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n352 GND 0.01fF
C5565 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n353 GND 0.01fF
C5566 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n354 GND 0.01fF
C5567 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n355 GND 0.01fF
C5568 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n356 GND 0.01fF
C5569 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n357 GND 0.01fF
C5570 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n358 GND 0.01fF
C5571 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n359 GND 0.01fF
C5572 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n360 GND 0.01fF
C5573 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n361 GND 0.00fF
C5574 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n362 GND 0.01fF
C5575 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n363 GND 0.01fF
C5576 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n364 GND 0.01fF
C5577 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n365 GND 0.04fF
C5578 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n366 GND 0.03fF
C5579 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n367 GND 0.01fF
C5580 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n368 GND 0.00fF
C5581 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n369 GND 0.01fF
C5582 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n370 GND 0.01fF
C5583 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n371 GND 0.01fF
C5584 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n372 GND 0.01fF
C5585 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n373 GND 0.00fF
C5586 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n374 GND 0.00fF
C5587 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n375 GND 0.00fF
C5588 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n376 GND 0.00fF
C5589 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n378 GND 0.02fF
C5590 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n379 GND 0.01fF
C5591 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n380 GND 0.01fF
C5592 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n381 GND 0.00fF
C5593 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n382 GND 0.00fF
C5594 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n383 GND 0.00fF
C5595 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n384 GND 0.01fF
C5596 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t13 GND 0.10fF $ **FLOATING
C5597 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n385 GND 0.08fF
C5598 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n386 GND 0.03fF
C5599 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n387 GND 0.04fF
C5600 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n388 GND 0.01fF
C5601 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n389 GND 0.00fF
C5602 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n390 GND 0.00fF
C5603 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n391 GND 0.00fF
C5604 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n392 GND 0.00fF
C5605 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n393 GND 0.01fF
C5606 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n394 GND 0.01fF
C5607 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n395 GND 0.01fF
C5608 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n396 GND 0.00fF
C5609 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n397 GND 0.01fF
C5610 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n398 GND 0.03fF
C5611 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n399 GND 0.00fF
C5612 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n400 GND 0.01fF
C5613 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n401 GND 0.01fF
C5614 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n402 GND 0.01fF
C5615 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n403 GND 0.01fF
C5616 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n404 GND 0.01fF
C5617 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n405 GND 0.00fF
C5618 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t18 GND 0.10fF $ **FLOATING
C5619 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n406 GND 0.07fF
C5620 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n407 GND 0.02fF
C5621 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n408 GND 0.02fF
C5622 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n409 GND 0.01fF
C5623 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n410 GND 0.01fF
C5624 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n411 GND 0.01fF
C5625 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n412 GND 0.01fF
C5626 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n413 GND 0.00fF
C5627 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n414 GND 0.00fF
C5628 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n415 GND 0.00fF
C5629 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n416 GND 0.01fF
C5630 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n417 GND 0.01fF
C5631 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n419 GND 0.03fF
C5632 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n420 GND 0.01fF
C5633 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n421 GND 0.00fF
C5634 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n422 GND 0.01fF
C5635 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n423 GND 0.01fF
C5636 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n424 GND 0.01fF
C5637 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n425 GND 0.01fF
C5638 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n426 GND 0.00fF
C5639 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n427 GND 0.00fF
C5640 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n428 GND 0.00fF
C5641 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n429 GND 0.00fF
C5642 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n431 GND 0.02fF
C5643 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n432 GND 0.01fF
C5644 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n433 GND 0.01fF
C5645 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n434 GND 0.00fF
C5646 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n435 GND 0.00fF
C5647 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n436 GND 0.00fF
C5648 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n437 GND 0.01fF
C5649 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t16 GND 0.10fF $ **FLOATING
C5650 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n438 GND 0.08fF
C5651 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n439 GND 0.03fF
C5652 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n440 GND 0.04fF
C5653 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n441 GND 0.01fF
C5654 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n442 GND 0.00fF
C5655 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n443 GND 0.00fF
C5656 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n444 GND 0.00fF
C5657 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n445 GND 0.00fF
C5658 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n446 GND 0.01fF
C5659 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n447 GND 0.01fF
C5660 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n448 GND 0.01fF
C5661 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n449 GND 0.00fF
C5662 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n450 GND 0.01fF
C5663 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n451 GND 0.03fF
C5664 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n452 GND 0.00fF
C5665 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n453 GND 0.01fF
C5666 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n454 GND 0.01fF
C5667 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n455 GND 0.01fF
C5668 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n456 GND 0.01fF
C5669 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n457 GND 0.01fF
C5670 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n458 GND 0.00fF
C5671 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t20 GND 0.10fF $ **FLOATING
C5672 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n459 GND 0.07fF
C5673 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n460 GND 0.02fF
C5674 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n461 GND 0.02fF
C5675 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n462 GND 0.01fF
C5676 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n463 GND 0.01fF
C5677 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n464 GND 0.01fF
C5678 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n465 GND 0.01fF
C5679 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n466 GND 0.00fF
C5680 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n467 GND 0.00fF
C5681 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n468 GND 0.00fF
C5682 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n469 GND 0.01fF
C5683 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n470 GND 0.01fF
C5684 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n472 GND 0.03fF
C5685 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n473 GND 0.01fF
C5686 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n474 GND 0.00fF
C5687 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n475 GND 0.01fF
C5688 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n476 GND 0.01fF
C5689 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n477 GND 0.01fF
C5690 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n478 GND 0.01fF
C5691 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n479 GND 0.00fF
C5692 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n480 GND 0.00fF
C5693 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n481 GND 0.00fF
C5694 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n482 GND 0.00fF
C5695 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n484 GND 0.02fF
C5696 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n485 GND 0.01fF
C5697 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n486 GND 0.01fF
C5698 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n487 GND 0.00fF
C5699 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n488 GND 0.00fF
C5700 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n489 GND 0.00fF
C5701 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n490 GND 0.01fF
C5702 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t10 GND 0.10fF $ **FLOATING
C5703 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n491 GND 0.08fF
C5704 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n492 GND 0.03fF
C5705 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n493 GND 0.04fF
C5706 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n494 GND 0.01fF
C5707 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n495 GND 0.00fF
C5708 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n496 GND 0.00fF
C5709 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n497 GND 0.00fF
C5710 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n498 GND 0.00fF
C5711 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n499 GND 0.01fF
C5712 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n500 GND 0.01fF
C5713 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n501 GND 0.01fF
C5714 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n502 GND 0.00fF
C5715 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n503 GND 0.01fF
C5716 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n504 GND 0.03fF
C5717 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n505 GND 0.00fF
C5718 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n506 GND 0.01fF
C5719 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n507 GND 0.01fF
C5720 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n508 GND 0.01fF
C5721 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n509 GND 0.01fF
C5722 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t7 GND 0.10fF $ **FLOATING
C5723 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n510 GND 0.07fF
C5724 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n511 GND 0.02fF
C5725 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n512 GND 0.01fF
C5726 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n513 GND 0.00fF
C5727 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n514 GND 0.02fF
C5728 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n515 GND 0.01fF
C5729 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n516 GND 0.01fF
C5730 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n517 GND 0.01fF
C5731 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n518 GND 0.01fF
C5732 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n519 GND 0.00fF
C5733 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n520 GND 0.00fF
C5734 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n521 GND 0.00fF
C5735 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n522 GND 0.01fF
C5736 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n523 GND 0.01fF
C5737 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n525 GND 0.04fF
C5738 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n526 GND 0.01fF
C5739 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n527 GND 0.01fF
C5740 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n528 GND 0.01fF
C5741 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n529 GND 0.02fF
C5742 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n530 GND 0.01fF
C5743 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n531 GND 0.01fF
C5744 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n532 GND 0.10fF
C5745 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n533 GND 0.10fF
C5746 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n534 GND 0.01fF
C5747 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n535 GND 0.01fF
C5748 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n536 GND 0.01fF
C5749 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n537 GND 0.01fF
C5750 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n538 GND 0.02fF
C5751 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n539 GND 0.01fF
C5752 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n540 GND 0.01fF
C5753 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n541 GND 0.23fF
C5754 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n542 GND 0.23fF
C5755 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n543 GND 0.01fF
C5756 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n544 GND 0.01fF
C5757 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n545 GND 0.01fF
C5758 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n546 GND 0.01fF
C5759 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n547 GND 0.02fF
C5760 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n548 GND 0.01fF
C5761 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n549 GND 0.01fF
C5762 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n550 GND 0.09fF
C5763 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n551 GND 0.09fF
C5764 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n552 GND 0.01fF
C5765 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n553 GND 0.02fF
C5766 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n554 GND 0.03fF
C5767 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n555 GND 0.01fF
C5768 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n556 GND 0.13fF
C5769 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n557 GND 0.04fF
C5770 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n558 GND 0.33fF
C5771 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n559 GND 0.03fF
C5772 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n560 GND 0.01fF
C5773 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n561 GND 0.00fF
C5774 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_8/GATE GND 0.02fF
C5775 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n562 GND 0.07fF
C5776 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n563 GND 0.02fF
C5777 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n564 GND 0.01fF
C5778 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n565 GND 0.00fF
C5779 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n566 GND 0.02fF
C5780 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n567 GND 0.01fF
C5781 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n568 GND 0.01fF
C5782 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n569 GND 0.01fF
C5783 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n570 GND 0.00fF
C5784 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n571 GND 0.00fF
C5785 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n572 GND 0.01fF
C5786 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n573 GND 0.01fF
C5787 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n574 GND 0.01fF
C5788 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n575 GND 0.01fF
C5789 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n576 GND 0.01fF
C5790 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n577 GND 0.01fF
C5791 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n578 GND 0.00fF
C5792 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n579 GND 0.00fF
C5793 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n580 GND 0.01fF
C5794 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n581 GND 0.00fF
C5795 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n582 GND 0.07fF
C5796 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n583 GND 0.02fF
C5797 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n584 GND 0.02fF
C5798 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n585 GND 0.03fF
C5799 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n586 GND 0.01fF
C5800 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n587 GND 0.01fF
C5801 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n588 GND 0.01fF
C5802 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n589 GND 0.01fF
C5803 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n590 GND 0.01fF
C5804 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n591 GND 0.03fF
C5805 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n592 GND 0.01fF
C5806 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n593 GND 0.01fF
C5807 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n594 GND 0.01fF
C5808 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n595 GND 0.01fF
C5809 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n596 GND 0.01fF
C5810 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n597 GND 0.00fF
C5811 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n598 GND 0.01fF
C5812 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n599 GND 0.01fF
C5813 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n600 GND 0.01fF
C5814 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n601 GND 0.04fF
C5815 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n602 GND 0.00fF
C5816 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n603 GND 0.01fF
C5817 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n604 GND 0.01fF
C5818 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n605 GND 0.01fF
C5819 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n606 GND 0.01fF
C5820 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n607 GND 0.00fF
C5821 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n608 GND 0.00fF
C5822 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n609 GND 0.00fF
C5823 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n610 GND 0.00fF
C5824 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n611 GND 0.03fF
C5825 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n612 GND 0.01fF
C5826 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n614 GND 0.02fF
C5827 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n615 GND 0.01fF
C5828 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n616 GND 0.01fF
C5829 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n617 GND 0.00fF
C5830 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n618 GND 0.00fF
C5831 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n619 GND 0.00fF
C5832 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n620 GND 0.01fF
C5833 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n621 GND 0.08fF
C5834 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n622 GND 0.03fF
C5835 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n623 GND 0.04fF
C5836 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n624 GND 0.01fF
C5837 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n625 GND 0.00fF
C5838 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n626 GND 0.00fF
C5839 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n627 GND 0.00fF
C5840 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n628 GND 0.00fF
C5841 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n629 GND 0.01fF
C5842 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n630 GND 0.01fF
C5843 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n631 GND 0.01fF
C5844 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n632 GND 0.00fF
C5845 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n633 GND 0.01fF
C5846 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n634 GND 0.03fF
C5847 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n635 GND 0.00fF
C5848 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n636 GND 0.01fF
C5849 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n637 GND 0.01fF
C5850 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n638 GND 0.01fF
C5851 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE GND 0.01fF
C5852 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n639 GND 0.01fF
C5853 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n640 GND 0.07fF
C5854 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n641 GND 0.02fF
C5855 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n642 GND 0.01fF
C5856 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n643 GND 0.00fF
C5857 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n644 GND 0.02fF
C5858 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n645 GND 0.01fF
C5859 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n646 GND 0.01fF
C5860 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n647 GND 0.01fF
C5861 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n648 GND 0.01fF
C5862 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n649 GND 0.00fF
C5863 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n650 GND 0.00fF
C5864 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n651 GND 0.00fF
C5865 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n652 GND 0.01fF
C5866 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n653 GND 0.01fF
C5867 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n655 GND 0.00fF
C5868 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n656 GND 0.01fF
C5869 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n657 GND 0.01fF
C5870 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n658 GND 0.01fF
C5871 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n659 GND 0.01fF
C5872 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n660 GND 0.00fF
C5873 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n661 GND 0.00fF
C5874 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n662 GND 0.00fF
C5875 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n663 GND 0.00fF
C5876 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n664 GND 0.03fF
C5877 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n665 GND 0.01fF
C5878 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n667 GND 0.02fF
C5879 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n668 GND 0.01fF
C5880 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n669 GND 0.01fF
C5881 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n670 GND 0.00fF
C5882 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n671 GND 0.00fF
C5883 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n672 GND 0.00fF
C5884 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n673 GND 0.01fF
C5885 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n674 GND 0.08fF
C5886 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n675 GND 0.03fF
C5887 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n676 GND 0.04fF
C5888 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n677 GND 0.01fF
C5889 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n678 GND 0.00fF
C5890 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n679 GND 0.00fF
C5891 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n680 GND 0.00fF
C5892 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n681 GND 0.00fF
C5893 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n682 GND 0.01fF
C5894 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n683 GND 0.01fF
C5895 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n684 GND 0.01fF
C5896 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n685 GND 0.00fF
C5897 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n686 GND 0.01fF
C5898 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n687 GND 0.03fF
C5899 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n688 GND 0.00fF
C5900 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n689 GND 0.01fF
C5901 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n690 GND 0.01fF
C5902 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n691 GND 0.01fF
C5903 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n692 GND 0.01fF
C5904 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n693 GND 0.01fF
C5905 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n694 GND 0.00fF
C5906 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n695 GND 0.07fF
C5907 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n696 GND 0.02fF
C5908 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n697 GND 0.02fF
C5909 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n698 GND 0.01fF
C5910 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n699 GND 0.01fF
C5911 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n700 GND 0.01fF
C5912 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n701 GND 0.01fF
C5913 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n702 GND 0.00fF
C5914 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n703 GND 0.00fF
C5915 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n704 GND 0.00fF
C5916 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n705 GND 0.01fF
C5917 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n706 GND 0.01fF
C5918 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n708 GND 0.00fF
C5919 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n709 GND 0.01fF
C5920 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n710 GND 0.01fF
C5921 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n711 GND 0.01fF
C5922 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n712 GND 0.01fF
C5923 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n713 GND 0.00fF
C5924 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n714 GND 0.00fF
C5925 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n715 GND 0.00fF
C5926 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n716 GND 0.00fF
C5927 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n717 GND 0.03fF
C5928 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n718 GND 0.01fF
C5929 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n720 GND 0.02fF
C5930 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n721 GND 0.01fF
C5931 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n722 GND 0.01fF
C5932 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n723 GND 0.00fF
C5933 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n724 GND 0.00fF
C5934 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n725 GND 0.00fF
C5935 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n726 GND 0.01fF
C5936 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n727 GND 0.08fF
C5937 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n728 GND 0.03fF
C5938 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n729 GND 0.04fF
C5939 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n730 GND 0.01fF
C5940 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n731 GND 0.00fF
C5941 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n732 GND 0.00fF
C5942 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n733 GND 0.00fF
C5943 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n734 GND 0.00fF
C5944 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n735 GND 0.01fF
C5945 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n736 GND 0.01fF
C5946 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n737 GND 0.01fF
C5947 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n738 GND 0.00fF
C5948 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n739 GND 0.01fF
C5949 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n740 GND 0.03fF
C5950 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n741 GND 0.00fF
C5951 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n742 GND 0.01fF
C5952 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n743 GND 0.01fF
C5953 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n744 GND 0.01fF
C5954 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_11/GATE GND 0.01fF
C5955 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n745 GND 0.01fF
C5956 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n746 GND 0.07fF
C5957 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n747 GND 0.02fF
C5958 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n748 GND 0.01fF
C5959 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n749 GND 0.00fF
C5960 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n750 GND 0.02fF
C5961 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n751 GND 0.01fF
C5962 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n752 GND 0.01fF
C5963 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n753 GND 0.01fF
C5964 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n754 GND 0.01fF
C5965 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n755 GND 0.00fF
C5966 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n756 GND 0.00fF
C5967 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n757 GND 0.00fF
C5968 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n758 GND 0.01fF
C5969 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n759 GND 0.01fF
C5970 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n761 GND 0.00fF
C5971 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n762 GND 0.01fF
C5972 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n763 GND 0.01fF
C5973 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n764 GND 0.01fF
C5974 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n765 GND 0.01fF
C5975 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n766 GND 0.00fF
C5976 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n767 GND 0.00fF
C5977 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n768 GND 0.00fF
C5978 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n769 GND 0.00fF
C5979 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n770 GND 0.03fF
C5980 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n771 GND 0.01fF
C5981 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n773 GND 0.02fF
C5982 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n774 GND 0.01fF
C5983 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n775 GND 0.01fF
C5984 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n776 GND 0.00fF
C5985 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n777 GND 0.00fF
C5986 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n778 GND 0.00fF
C5987 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n779 GND 0.01fF
C5988 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n780 GND 0.08fF
C5989 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n781 GND 0.03fF
C5990 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n782 GND 0.04fF
C5991 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n783 GND 0.01fF
C5992 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n784 GND 0.00fF
C5993 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n785 GND 0.00fF
C5994 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n786 GND 0.00fF
C5995 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n787 GND 0.00fF
C5996 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n788 GND 0.01fF
C5997 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n789 GND 0.01fF
C5998 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n790 GND 0.01fF
C5999 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n791 GND 0.00fF
C6000 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n792 GND 0.01fF
C6001 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n793 GND 0.03fF
C6002 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n794 GND 0.00fF
C6003 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n795 GND 0.01fF
C6004 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n796 GND 0.01fF
C6005 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n797 GND 0.01fF
C6006 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_12/GATE GND 0.01fF
C6007 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n798 GND 0.01fF
C6008 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n799 GND 0.01fF
C6009 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n800 GND 0.00fF
C6010 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n801 GND 0.07fF
C6011 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n802 GND 0.02fF
C6012 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n803 GND 0.02fF
C6013 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n804 GND 0.01fF
C6014 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n805 GND 0.01fF
C6015 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n806 GND 0.01fF
C6016 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n807 GND 0.01fF
C6017 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n808 GND 0.00fF
C6018 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n809 GND 0.00fF
C6019 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n810 GND 0.00fF
C6020 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n811 GND 0.01fF
C6021 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n812 GND 0.01fF
C6022 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n814 GND 0.04fF
C6023 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n815 GND 0.01fF
C6024 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n816 GND 0.01fF
C6025 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n817 GND 0.01fF
C6026 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n818 GND 0.02fF
C6027 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n819 GND 0.01fF
C6028 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n820 GND 0.01fF
C6029 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n821 GND 0.10fF
C6030 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n822 GND 0.10fF
C6031 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n823 GND 0.01fF
C6032 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n824 GND 0.01fF
C6033 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n825 GND 0.01fF
C6034 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n826 GND 0.01fF
C6035 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n827 GND 0.02fF
C6036 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n828 GND 0.01fF
C6037 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n829 GND 0.01fF
C6038 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n830 GND 0.10fF
C6039 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n831 GND 0.10fF
C6040 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n832 GND 0.01fF
C6041 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n833 GND 0.01fF
C6042 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n834 GND 0.01fF
C6043 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n835 GND 0.01fF
C6044 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n836 GND 0.02fF
C6045 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n837 GND 0.01fF
C6046 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n838 GND 0.01fF
C6047 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n839 GND 0.10fF
C6048 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n840 GND 0.10fF
C6049 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n841 GND 0.01fF
C6050 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n842 GND 0.01fF
C6051 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n843 GND 0.01fF
C6052 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n844 GND 0.01fF
C6053 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n845 GND 0.02fF
C6054 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n846 GND 0.01fF
C6055 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n847 GND 0.01fF
C6056 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n848 GND 0.09fF
C6057 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n849 GND 0.09fF
C6058 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n850 GND 0.01fF
C6059 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n851 GND 0.02fF
C6060 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n852 GND 0.03fF
C6061 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n853 GND 0.01fF
C6062 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n854 GND 0.13fF
C6063 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n855 GND 0.04fF
C6064 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n856 GND 0.32fF
C6065 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n857 GND 0.03fF
C6066 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n858 GND 0.01fF
C6067 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n859 GND 0.00fF
C6068 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n860 GND 0.01fF
C6069 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n861 GND 0.00fF
C6070 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t8 GND 0.10fF $ **FLOATING
C6071 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n862 GND 0.07fF
C6072 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n863 GND 0.02fF
C6073 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n864 GND 0.02fF
C6074 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n865 GND 0.01fF
C6075 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n866 GND 0.01fF
C6076 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n867 GND 0.01fF
C6077 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n868 GND 0.00fF
C6078 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n869 GND 0.00fF
C6079 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n870 GND 0.01fF
C6080 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n871 GND 0.01fF
C6081 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n872 GND 0.01fF
C6082 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n873 GND 0.01fF
C6083 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n874 GND 0.01fF
C6084 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n875 GND 0.01fF
C6085 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n876 GND 0.00fF
C6086 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n877 GND 0.00fF
C6087 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n878 GND 0.01fF
C6088 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n879 GND 0.00fF
C6089 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t14 GND 0.10fF $ **FLOATING
C6090 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n880 GND 0.07fF
C6091 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n881 GND 0.02fF
C6092 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n882 GND 0.02fF
C6093 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n883 GND 0.03fF
C6094 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n884 GND 0.01fF
C6095 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n885 GND 0.01fF
C6096 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n886 GND 0.01fF
C6097 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n887 GND 0.01fF
C6098 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n888 GND 0.01fF
C6099 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n889 GND 0.03fF
C6100 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n890 GND 0.01fF
C6101 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n891 GND 0.01fF
C6102 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n892 GND 0.01fF
C6103 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n893 GND 0.01fF
C6104 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n894 GND 0.01fF
C6105 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n895 GND 0.00fF
C6106 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n896 GND 0.01fF
C6107 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n897 GND 0.01fF
C6108 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n898 GND 0.01fF
C6109 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n899 GND 0.04fF
C6110 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n900 GND 0.04fF
C6111 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n901 GND 0.01fF
C6112 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n902 GND 0.02fF
C6113 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n903 GND 0.01fF
C6114 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n904 GND 0.00fF
C6115 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t5 GND 0.10fF $ **FLOATING
C6116 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n905 GND 0.08fF
C6117 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n906 GND 0.03fF
C6118 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n907 GND 0.04fF
C6119 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n908 GND 0.01fF
C6120 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n909 GND 0.00fF
C6121 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n910 GND 0.03fF
C6122 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n911 GND 0.00fF
C6123 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n912 GND 0.01fF
C6124 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n913 GND 0.00fF
C6125 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n914 GND 0.01fF
C6126 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n915 GND 0.01fF
C6127 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n916 GND 0.00fF
C6128 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n917 GND 0.01fF
C6129 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n918 GND 0.00fF
C6130 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n919 GND 0.01fF
C6131 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n920 GND 0.04fF
C6132 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n921 GND 0.01fF
C6133 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n922 GND 0.01fF
C6134 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n923 GND 0.01fF
C6135 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n924 GND 0.01fF
C6136 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n925 GND 0.00fF
C6137 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t19 GND 0.10fF $ **FLOATING
C6138 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n926 GND 0.07fF
C6139 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n927 GND 0.02fF
C6140 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n928 GND 0.02fF
C6141 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n929 GND 0.01fF
C6142 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n930 GND 0.01fF
C6143 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n931 GND 0.01fF
C6144 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n932 GND 0.01fF
C6145 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n933 GND 0.00fF
C6146 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n934 GND 0.00fF
C6147 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n935 GND 0.01fF
C6148 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n936 GND 0.01fF
C6149 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n938 GND 0.04fF
C6150 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n939 GND 0.01fF
C6151 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n940 GND 0.02fF
C6152 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n941 GND 0.01fF
C6153 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n942 GND 0.00fF
C6154 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t15 GND 0.10fF $ **FLOATING
C6155 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n943 GND 0.08fF
C6156 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n944 GND 0.03fF
C6157 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n945 GND 0.04fF
C6158 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n946 GND 0.00fF
C6159 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n947 GND 0.03fF
C6160 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n948 GND 0.00fF
C6161 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n949 GND 0.01fF
C6162 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n950 GND 0.00fF
C6163 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n951 GND 0.01fF
C6164 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n952 GND 0.01fF
C6165 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n953 GND 0.01fF
C6166 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n954 GND 0.00fF
C6167 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n955 GND 0.01fF
C6168 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n956 GND 0.00fF
C6169 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n957 GND 0.01fF
C6170 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n958 GND 0.04fF
C6171 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n959 GND 0.01fF
C6172 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n960 GND 0.01fF
C6173 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n961 GND 0.01fF
C6174 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n962 GND 0.01fF
C6175 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n963 GND 0.00fF
C6176 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t6 GND 0.10fF $ **FLOATING
C6177 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n964 GND 0.07fF
C6178 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n965 GND 0.02fF
C6179 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n966 GND 0.02fF
C6180 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n967 GND 0.01fF
C6181 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n968 GND 0.01fF
C6182 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n969 GND 0.01fF
C6183 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n970 GND 0.01fF
C6184 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n971 GND 0.00fF
C6185 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n972 GND 0.00fF
C6186 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n973 GND 0.01fF
C6187 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n974 GND 0.01fF
C6188 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n976 GND 0.04fF
C6189 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n977 GND 0.01fF
C6190 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n978 GND 0.02fF
C6191 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n979 GND 0.01fF
C6192 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n980 GND 0.00fF
C6193 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t17 GND 0.10fF $ **FLOATING
C6194 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n981 GND 0.08fF
C6195 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n982 GND 0.03fF
C6196 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n983 GND 0.04fF
C6197 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n984 GND 0.00fF
C6198 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n985 GND 0.03fF
C6199 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n986 GND 0.00fF
C6200 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n987 GND 0.01fF
C6201 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n988 GND 0.00fF
C6202 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n989 GND 0.01fF
C6203 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n990 GND 0.01fF
C6204 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n991 GND 0.01fF
C6205 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n992 GND 0.00fF
C6206 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n993 GND 0.01fF
C6207 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n994 GND 0.00fF
C6208 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n995 GND 0.01fF
C6209 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n996 GND 0.04fF
C6210 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n997 GND 0.01fF
C6211 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n998 GND 0.01fF
C6212 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n999 GND 0.01fF
C6213 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.t12 GND 0.10fF $ **FLOATING
C6214 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1000 GND 0.07fF
C6215 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1001 GND 0.02fF
C6216 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1002 GND 0.01fF
C6217 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1003 GND 0.00fF
C6218 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1004 GND 0.02fF
C6219 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1005 GND 0.01fF
C6220 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1006 GND 0.01fF
C6221 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1007 GND 0.01fF
C6222 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1008 GND 0.01fF
C6223 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1009 GND 0.00fF
C6224 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1010 GND 0.00fF
C6225 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1011 GND 0.01fF
C6226 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1012 GND 0.01fF
C6227 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1013 GND 0.01fF
C6228 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1014 GND 0.07fF
C6229 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1015 GND 0.03fF
C6230 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1016 GND 0.10fF
C6231 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1017 GND 0.11fF
C6232 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1018 GND 0.03fF
C6233 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1019 GND 0.03fF
C6234 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1020 GND 0.23fF
C6235 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1021 GND 0.24fF
C6236 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1022 GND 0.03fF
C6237 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1023 GND 0.03fF
C6238 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1024 GND 0.09fF
C6239 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1025 GND 0.09fF
C6240 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1026 GND 0.01fF
C6241 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1027 GND 0.02fF
C6242 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1028 GND 0.03fF
C6243 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1029 GND 0.01fF
C6244 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1030 GND 0.13fF
C6245 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1031 GND 0.04fF
C6246 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1032 GND 0.59fF
C6247 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1033 GND 2.90fF
C6248 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1034 GND 0.58fF
C6249 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1036 GND 0.03fF
C6250 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1037 GND 0.03fF
C6251 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_5/GATE.n1038 GND 0.10fF
C6252 vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_10/DRAIN GND 0.09fF
.ends
