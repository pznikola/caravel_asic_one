* NGSPICE file created from vco_pmirr.ext - technology: sky130B

.subckt rf_pfet_01v8_aM02W3p00L0p15 GATE DRAIN SOURCE BULK
X0 SOURCE GATE DRAIN BULK sky130_fd_pr__pfet_01v8 ad=1.6856e+12p pd=1.316e+07u as=8.428e+11p ps=6.58e+06u w=3.01e+06u l=150000u
X1 DRAIN GATE SOURCE BULK sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.01e+06u l=150000u
.ends

.subckt vco_pmirr_base rf_pfet_01v8_aM02W3p00L0p15_10/SOURCE rf_pfet_01v8_aM02W3p00L0p15_1/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_10/DRAIN rf_pfet_01v8_aM02W3p00L0p15_2/DRAIN rf_pfet_01v8_aM02W3p00L0p15_11/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_5/SOURCE rf_pfet_01v8_aM02W3p00L0p15_12/DRAIN rf_pfet_01v8_aM02W3p00L0p15_4/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_5/DRAIN rf_pfet_01v8_aM02W3p00L0p15_10/GATE rf_pfet_01v8_aM02W3p00L0p15_4/GATE
+ rf_pfet_01v8_aM02W3p00L0p15_4/SOURCE rf_pfet_01v8_aM02W3p00L0p15_8/DRAIN rf_pfet_01v8_aM02W3p00L0p15_1/GATE
+ rf_pfet_01v8_aM02W3p00L0p15_9/DRAIN rf_pfet_01v8_aM02W3p00L0p15_9/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK
+ rf_pfet_01v8_aM02W3p00L0p15_8/GATE rf_pfet_01v8_aM02W3p00L0p15_11/GATE rf_pfet_01v8_aM02W3p00L0p15_5/GATE
+ rf_pfet_01v8_aM02W3p00L0p15_8/SOURCE rf_pfet_01v8_aM02W3p00L0p15_2/GATE rf_pfet_01v8_aM02W3p00L0p15_12/SOURCE
+ rf_pfet_01v8_aM02W3p00L0p15_2/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/GATE rf_pfet_01v8_aM02W3p00L0p15_1/SOURCE
+ rf_pfet_01v8_aM02W3p00L0p15_11/SOURCE rf_pfet_01v8_aM02W3p00L0p15_12/GATE
Xrf_pfet_01v8_aM02W3p00L0p15_8 rf_pfet_01v8_aM02W3p00L0p15_8/GATE rf_pfet_01v8_aM02W3p00L0p15_8/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_8/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_9 rf_pfet_01v8_aM02W3p00L0p15_9/GATE rf_pfet_01v8_aM02W3p00L0p15_9/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_9/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_10 rf_pfet_01v8_aM02W3p00L0p15_10/GATE rf_pfet_01v8_aM02W3p00L0p15_10/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_10/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_11 rf_pfet_01v8_aM02W3p00L0p15_11/GATE rf_pfet_01v8_aM02W3p00L0p15_11/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_11/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_12 rf_pfet_01v8_aM02W3p00L0p15_12/GATE rf_pfet_01v8_aM02W3p00L0p15_12/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_12/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_13 rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK
+ rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_0 rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK
+ rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_1 rf_pfet_01v8_aM02W3p00L0p15_1/GATE rf_pfet_01v8_aM02W3p00L0p15_1/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_1/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_3 rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK
+ rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_2 rf_pfet_01v8_aM02W3p00L0p15_2/GATE rf_pfet_01v8_aM02W3p00L0p15_2/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_2/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_4 rf_pfet_01v8_aM02W3p00L0p15_4/GATE rf_pfet_01v8_aM02W3p00L0p15_4/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_4/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_5 rf_pfet_01v8_aM02W3p00L0p15_5/GATE rf_pfet_01v8_aM02W3p00L0p15_5/DRAIN
+ rf_pfet_01v8_aM02W3p00L0p15_5/SOURCE rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_6 rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK
+ rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
Xrf_pfet_01v8_aM02W3p00L0p15_7 rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK
+ rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15_9/BULK rf_pfet_01v8_aM02W3p00L0p15
.ends

.subckt sky130_fd_pr__res_high_po_2p85_5ZUK6C a_n415_n912# a_n285_350# a_n285_n782#
X0 a_n285_n782# a_n285_350# a_n415_n912# sky130_fd_pr__res_high_po_2p85 l=3.5e+06u
.ends

.subckt vco_pmirr IND_CT VBIAS VDD GND
Xvco_pmirr_base_0 VDD IND_CT vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE IND_CT
+ IND_CT VDD IND_CT IND_CT IND_CT vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE
+ vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE VDD IND_CT vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE
+ IND_CT VDD VDD vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE
+ vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE VDD vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE
+ VDD VDD vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE VDD VDD vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE
+ vco_pmirr_base
Xsky130_fd_pr__res_high_po_2p85_5ZUK6C_0 GND vco_pmirr_base_0/rf_pfet_01v8_aM02W3p00L0p15_9/GATE
+ VBIAS sky130_fd_pr__res_high_po_2p85_5ZUK6C
.ends

