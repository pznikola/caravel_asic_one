magic
tech sky130B
magscale 1 2
timestamp 1654419893
<< pwell >>
rect -96 -34 814 1130
<< nmos >>
rect 302 92 332 422
rect 388 92 418 422
<< ndiff >>
rect 246 410 302 422
rect 246 376 257 410
rect 291 376 302 410
rect 246 342 302 376
rect 246 308 257 342
rect 291 308 302 342
rect 246 274 302 308
rect 246 240 257 274
rect 291 240 302 274
rect 246 206 302 240
rect 246 172 257 206
rect 291 172 302 206
rect 246 138 302 172
rect 246 104 257 138
rect 291 104 302 138
rect 246 92 302 104
rect 332 410 388 422
rect 332 376 343 410
rect 377 376 388 410
rect 332 342 388 376
rect 332 308 343 342
rect 377 308 388 342
rect 332 274 388 308
rect 332 240 343 274
rect 377 240 388 274
rect 332 206 388 240
rect 332 172 343 206
rect 377 172 388 206
rect 332 138 388 172
rect 332 104 343 138
rect 377 104 388 138
rect 332 92 388 104
rect 418 410 474 422
rect 418 376 429 410
rect 463 376 474 410
rect 418 342 474 376
rect 418 308 429 342
rect 463 308 474 342
rect 418 274 474 308
rect 418 240 429 274
rect 463 240 474 274
rect 418 206 474 240
rect 418 172 429 206
rect 463 172 474 206
rect 418 138 474 172
rect 418 104 429 138
rect 463 104 474 138
rect 418 92 474 104
<< ndiffc >>
rect 257 376 291 410
rect 257 308 291 342
rect 257 240 291 274
rect 257 172 291 206
rect 257 104 291 138
rect 343 376 377 410
rect 343 308 377 342
rect 343 240 377 274
rect 343 172 377 206
rect 343 104 377 138
rect 429 376 463 410
rect 429 308 463 342
rect 429 240 463 274
rect 429 172 463 206
rect 429 104 463 138
<< psubdiff >>
rect 134 376 192 422
rect 134 342 146 376
rect 180 342 192 376
rect 134 308 192 342
rect 134 274 146 308
rect 180 274 192 308
rect 134 240 192 274
rect 134 206 146 240
rect 180 206 192 240
rect 134 172 192 206
rect 134 138 146 172
rect 180 138 192 172
rect 134 92 192 138
rect 528 376 586 422
rect 528 342 540 376
rect 574 342 586 376
rect 528 308 586 342
rect 528 274 540 308
rect 574 274 586 308
rect 528 240 586 274
rect 528 206 540 240
rect 574 206 586 240
rect 528 172 586 206
rect 528 138 540 172
rect 574 138 586 172
rect 528 92 586 138
<< psubdiffcont >>
rect 146 342 180 376
rect 146 274 180 308
rect 146 206 180 240
rect 146 138 180 172
rect 540 342 574 376
rect 540 274 574 308
rect 540 206 574 240
rect 540 138 574 172
<< poly >>
rect 259 494 461 514
rect 259 460 275 494
rect 309 460 343 494
rect 377 460 411 494
rect 445 460 461 494
rect 259 444 461 460
rect 302 422 332 444
rect 388 422 418 444
rect 302 70 332 92
rect 388 70 418 92
rect 259 54 461 70
rect 259 20 275 54
rect 309 20 343 54
rect 377 20 411 54
rect 445 20 461 54
rect 259 0 461 20
<< polycont >>
rect 275 460 309 494
rect 343 460 377 494
rect 411 460 445 494
rect 275 20 309 54
rect 343 20 377 54
rect 411 20 445 54
<< xpolycontact >>
rect -44 648 26 1080
rect 694 648 764 1080
rect -44 16 26 448
rect 694 16 764 448
<< xpolyres >>
rect -44 448 26 648
rect 694 448 764 648
<< locali >>
rect 259 460 271 494
rect 309 460 343 494
rect 377 460 411 494
rect 449 460 461 494
rect 257 410 291 426
rect 146 382 180 392
rect 146 310 180 342
rect 146 240 180 274
rect 146 172 180 204
rect 146 122 180 132
rect 257 342 291 348
rect 257 274 291 276
rect 257 238 291 240
rect 257 166 291 172
rect 257 88 291 104
rect 343 410 377 426
rect 343 342 377 348
rect 343 274 377 276
rect 343 238 377 240
rect 343 166 377 172
rect 343 88 377 104
rect 429 410 463 426
rect 429 342 463 348
rect 429 274 463 276
rect 429 238 463 240
rect 429 166 463 172
rect 540 382 574 392
rect 540 310 574 342
rect 540 240 574 274
rect 540 172 574 204
rect 540 122 574 132
rect 429 88 463 104
rect 259 20 271 54
rect 309 20 343 54
rect 377 20 411 54
rect 449 20 461 54
<< viali >>
rect -28 665 10 1062
rect 710 665 748 1062
rect 271 460 275 494
rect 275 460 305 494
rect 343 460 377 494
rect 415 460 445 494
rect 445 460 449 494
rect -28 34 10 431
rect 146 376 180 382
rect 146 348 180 376
rect 146 308 180 310
rect 146 276 180 308
rect 146 206 180 238
rect 146 204 180 206
rect 146 138 180 166
rect 146 132 180 138
rect 257 376 291 382
rect 257 348 291 376
rect 257 308 291 310
rect 257 276 291 308
rect 257 206 291 238
rect 257 204 291 206
rect 257 138 291 166
rect 257 132 291 138
rect 343 376 377 382
rect 343 348 377 376
rect 343 308 377 310
rect 343 276 377 308
rect 343 206 377 238
rect 343 204 377 206
rect 343 138 377 166
rect 343 132 377 138
rect 429 376 463 382
rect 429 348 463 376
rect 429 308 463 310
rect 429 276 463 308
rect 429 206 463 238
rect 429 204 463 206
rect 429 138 463 166
rect 429 132 463 138
rect 540 376 574 382
rect 540 348 574 376
rect 540 308 574 310
rect 540 276 574 308
rect 540 206 574 238
rect 540 204 574 206
rect 540 138 574 166
rect 540 132 574 138
rect 271 20 275 54
rect 275 20 305 54
rect 343 20 377 54
rect 415 20 445 54
rect 445 20 449 54
rect 710 34 748 431
<< metal1 >>
rect -4220 1062 4980 2920
rect -4220 920 -28 1062
rect -34 665 -28 920
rect 10 920 710 1062
rect 10 665 16 920
rect -34 653 16 665
rect 704 665 710 920
rect 748 920 4980 1062
rect 748 665 754 920
rect 704 653 754 665
rect 259 494 461 514
rect 259 460 271 494
rect 305 460 343 494
rect 377 460 415 494
rect 449 460 461 494
rect 259 448 461 460
rect -54 16 -44 448
rect 26 16 36 448
rect 134 382 192 410
rect 134 348 146 382
rect 180 348 192 382
rect 134 310 192 348
rect 134 276 146 310
rect 180 276 192 310
rect 134 238 192 276
rect 134 204 146 238
rect 180 204 192 238
rect 134 166 192 204
rect 134 132 146 166
rect 180 132 192 166
rect 134 104 192 132
rect 248 382 300 410
rect 248 348 257 382
rect 291 348 300 382
rect 248 310 300 348
rect 248 276 257 310
rect 291 276 300 310
rect 248 238 300 276
rect 248 226 257 238
rect 291 226 300 238
rect 248 166 300 174
rect 248 162 257 166
rect 291 162 300 166
rect 248 104 300 110
rect 334 404 386 410
rect 334 348 343 352
rect 377 348 386 352
rect 334 340 386 348
rect 334 276 343 288
rect 377 276 386 288
rect 334 238 386 276
rect 334 204 343 238
rect 377 204 386 238
rect 334 166 386 204
rect 334 132 343 166
rect 377 132 386 166
rect 334 104 386 132
rect 420 382 472 410
rect 420 348 429 382
rect 463 348 472 382
rect 420 310 472 348
rect 420 276 429 310
rect 463 276 472 310
rect 420 238 472 276
rect 420 226 429 238
rect 463 226 472 238
rect 420 166 472 174
rect 420 162 429 166
rect 463 162 472 166
rect 420 104 472 110
rect 528 382 586 410
rect 528 348 540 382
rect 574 348 586 382
rect 528 310 586 348
rect 528 276 540 310
rect 574 276 586 310
rect 528 238 586 276
rect 528 204 540 238
rect 574 204 586 238
rect 528 166 586 204
rect 528 132 540 166
rect 574 132 586 166
rect 528 104 586 132
rect 146 -70 180 104
rect 259 54 461 66
rect 259 20 271 54
rect 305 20 343 54
rect 377 20 415 54
rect 449 20 461 54
rect 259 0 461 20
rect 259 -60 273 0
rect 447 -60 461 0
rect 140 -130 180 -70
rect 540 -70 574 104
rect 684 16 694 448
rect 764 16 774 448
rect 540 -130 580 -70
rect 140 -2960 580 -130
rect -4220 -4960 4980 -2960
<< via1 >>
rect -44 431 26 448
rect -44 34 -28 431
rect -28 34 10 431
rect 10 34 26 431
rect -44 16 26 34
rect 248 204 257 226
rect 257 204 291 226
rect 291 204 300 226
rect 248 174 300 204
rect 248 132 257 162
rect 257 132 291 162
rect 291 132 300 162
rect 248 110 300 132
rect 334 382 386 404
rect 334 352 343 382
rect 343 352 377 382
rect 377 352 386 382
rect 334 310 386 340
rect 334 288 343 310
rect 343 288 377 310
rect 377 288 386 310
rect 420 204 429 226
rect 429 204 463 226
rect 463 204 472 226
rect 420 174 472 204
rect 420 132 429 162
rect 429 132 463 162
rect 463 132 472 162
rect 420 110 472 132
rect 273 -60 447 0
rect 694 431 764 448
rect 694 34 710 431
rect 710 34 748 431
rect 748 34 764 431
rect 694 16 764 34
<< metal2 >>
rect -44 448 26 458
rect -50 16 -44 410
rect 694 448 764 458
rect 26 404 612 410
rect 26 352 334 404
rect 386 352 612 404
rect 26 340 612 352
rect 26 288 334 340
rect 386 288 612 340
rect 26 282 612 288
rect 26 16 30 282
rect 108 226 694 232
rect 108 174 248 226
rect 300 174 420 226
rect 472 174 694 226
rect 108 162 694 174
rect 108 110 248 162
rect 300 110 420 162
rect 472 110 694 162
rect 108 104 694 110
rect -50 -240 30 16
rect 690 16 694 104
rect 764 16 770 232
rect -60 -260 30 -240
rect -60 -330 -50 -260
rect 20 -330 30 -260
rect -60 -340 30 -330
rect 270 0 450 10
rect 270 -60 273 0
rect 447 -60 450 0
rect 270 -460 450 -60
rect 690 -240 770 16
rect 690 -260 780 -240
rect 690 -330 700 -260
rect 770 -330 780 -260
rect 690 -340 780 -330
rect -4220 -2460 4980 -460
<< via2 >>
rect -50 -330 20 -260
rect 700 -330 770 -260
<< metal3 >>
rect -1135 832 -176 860
rect -1135 28 -260 832
rect -196 28 -176 832
rect -1135 0 -176 28
rect 944 832 1903 860
rect 944 28 964 832
rect 1028 28 1903 832
rect 944 0 1903 28
rect -280 -250 40 -240
rect -280 -340 -270 -250
rect -190 -260 40 -250
rect -190 -330 -50 -260
rect 20 -330 40 -260
rect -190 -340 40 -330
rect -280 -350 40 -340
rect 680 -250 1050 -240
rect 680 -260 960 -250
rect 680 -330 700 -260
rect 770 -330 960 -260
rect 680 -340 960 -330
rect 1040 -340 1050 -250
rect 680 -350 1050 -340
<< via3 >>
rect -260 28 -196 832
rect 964 28 1028 832
rect -270 -340 -190 -250
rect 960 -340 1040 -250
<< mimcap >>
rect -1035 720 -375 760
rect -1035 140 -995 720
rect -415 140 -375 720
rect -1035 100 -375 140
rect 1143 720 1803 760
rect 1143 140 1183 720
rect 1763 140 1803 720
rect 1143 100 1803 140
<< mimcapcontact >>
rect -995 140 -415 720
rect 1183 140 1763 720
<< metal4 >>
rect -3220 480 -1220 3920
rect -280 832 -180 850
rect 950 848 1050 850
rect -996 720 -414 721
rect -996 480 -995 720
rect -3220 380 -995 480
rect -3220 -5960 -1220 380
rect -996 140 -995 380
rect -415 140 -414 720
rect -996 139 -414 140
rect -280 28 -260 832
rect -196 28 -180 832
rect -280 -250 -180 28
rect 948 832 1050 848
rect 948 28 964 832
rect 1028 28 1050 832
rect 1182 720 1764 721
rect 1182 140 1183 720
rect 1763 480 1764 720
rect 1990 480 3990 3920
rect 1763 380 3990 480
rect 1763 140 1764 380
rect 1182 139 1764 140
rect 948 12 1050 28
rect -280 -340 -270 -250
rect -190 -340 -180 -250
rect -280 -350 -180 -340
rect 950 -250 1050 12
rect 950 -340 960 -250
rect 1040 -340 1050 -250
rect 950 -350 1050 -340
rect 1990 -2460 3990 380
rect 1980 -5960 3990 -2460
<< res0p35 >>
rect -46 446 28 650
rect 692 446 766 650
<< labels >>
flabel metal2 4980 -1500 4980 -1500 7 FreeSans 2400 0 0 0 ON
port 1 w
flabel metal1 4980 1860 4980 1860 7 FreeSans 2400 0 0 0 V_bias
port 2 w
flabel metal4 -2270 3920 -2270 3920 5 FreeSans 2400 0 0 0 OUT_P
port 3 s
flabel metal4 2990 3920 2990 3920 5 FreeSans 2400 0 0 0 OUT_N
port 4 s
flabel metal1 4980 -3960 4980 -3960 7 FreeSans 2400 0 0 0 GND
port 5 w
<< end >>
