* NGSPICE file created from capbank_pex.ext - technology: sky130B

.subckt capbank_pex OUT_P OUT_N bit0 bit1 bit2 bit3 bit4 bit5 VDD GND
X0 a_22576_45486.t1 bit4.t0 a_22866_45562.t2 GND.t96 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 OUT_P.t0 a_59376_45486.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X2 a_50176_5966.t2 bit5.t0 a_50466_6042.t1 GND.t161 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_4176_94886.t0 a_n436_94366.t0 GND.t0 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X4 OUT_P.t1 a_4176_55366.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X5 a_13666_15922.t2 bit5.t1 a_13376_15846.t1 GND.t208 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X6 a_4176_15846.t0 a_n436_5446.t8 GND.t15 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X7 a_31776_25726.t3 a_n436_5446.t43 GND.t154 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X8 OUT_P.t2 a_4176_94886.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X9 a_68866_45562.t3 a_n436_44966.t33 GND.t256 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X10 a_50176_45486.t1 bit4.t1 a_50466_45562.t1 GND.t95 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X11 OUT_P.t3 a_50176_55366.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X12 OUT_N.t0 a_68866_35682.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X13 OUT_P.t4 a_31776_45486.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X14 OUT_N.t1 a_59666_55442.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X15 a_13376_35606.t3 a_n436_5446.t65 GND.t263 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X16 a_41266_15922.t2 bit5.t2 a_40976_15846.t1 GND.t156 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X17 a_31776_55366.t1 bit4.t2 a_32066_55442.t1 GND.t94 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X18 a_4466_65322.t1 a_n436_64726.t5 GND.t51 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X19 OUT_P.t5 a_22576_55366.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X20 OUT_N.t2 a_50466_65322.t1 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X21 OUT_N.t3 a_4466_55442.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X22 a_13666_15922.t0 a_n436_5446.t9 GND.t26 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X23 a_4176_35606.t1 bit5.t3 a_4466_35682.t1 GND.t163 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X24 a_22866_25802.t2 bit5.t4 a_22576_25726.t1 GND.t216 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X25 a_4466_75202.t1 bit2.t0 a_4176_75126.t1 GND.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X26 OUT_N.t4 a_4466_94962.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X27 OUT_P.t6 a_13376_65246.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X28 OUT_N.t5 a_32066_45562.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X29 a_13376_55366.t1 bit4.t3 a_13666_55442.t1 GND.t93 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X30 a_4466_6042.t0 a_n436_5446.t10 GND.t27 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X31 a_40976_25726.t0 a_n436_5446.t11 GND.t28 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X32 a_68866_35682.t0 bit5.t5 a_68576_35606.t2 GND.t231 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X33 OUT_P.t7 a_40976_25726.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X34 a_32066_6042.t2 a_n436_5446.t26 GND.t62 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X35 OUT_N.t6 a_22866_55442.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X36 a_22576_35606.t2 a_n436_5446.t27 GND.t97 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X37 a_40976_55366.t1 bit4.t4 a_41266_55442.t0 GND.t92 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X38 a_50466_15922.t1 bit5.t6 a_50176_15846.t1 GND.t162 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X39 a_13376_45486.t2 a_n436_44966.t14 GND.t106 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X40 a_22866_6042.t1 bit5.t7 a_22576_5966.t1 GND.t141 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X41 OUT_N.t7 a_13666_65322.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X42 a_22866_15922.t2 a_n436_5446.t31 GND.t107 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X43 a_32066_25802.t1 bit5.t8 a_31776_25726.t1 GND.t209 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X44 a_50176_35606.t3 a_n436_5446.t57 GND.t185 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X45 a_59376_15846.t1 bit5.t9 a_59666_15922.t2 GND.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X46 a_59376_55366.t3 a_n436_44966.t29 GND.t177 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X47 a_22576_55366.t1 bit4.t5 a_22866_55442.t2 GND.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X48 OUT_N.t8 a_50466_15922.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X49 a_13666_25802.t1 bit5.t10 a_13376_25726.t1 GND.t40 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X50 a_4176_25726.t3 a_n436_5446.t54 GND.t178 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X51 a_31776_35606.t3 a_n436_5446.t42 GND.t152 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X52 OUT_N.t9 a_68866_6042.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X53 a_50176_55366.t1 bit4.t6 a_50466_55442.t1 GND.t90 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X54 OUT_P.t8 a_13376_15846.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X55 OUT_N.t10 a_41266_25802.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X56 a_22576_45486.t3 a_n436_44966.t26 GND.t153 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X57 a_32066_15922.t0 a_n436_5446.t17 GND.t52 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X58 GND.t124 bit3.t0 a_n436_64726.t9 GND.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X59 a_31776_65246.t1 bit3.t1 a_32066_65322.t1 GND.t125 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X60 a_41266_25802.t1 bit5.t11 a_40976_25726.t2 GND.t214 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X61 a_59666_35682.t2 bit5.t12 a_59376_35606.t2 GND.t215 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X62 a_68576_15846.t1 bit5.t13 a_68866_15922.t0 GND.t225 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X63 a_4466_75202.t3 a_n436_74606.t9 GND.t179 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X64 a_50176_45486.t3 a_n436_44966.t30 GND.t180 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X65 a_13666_25802.t3 a_n436_5446.t55 GND.t181 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X66 a_4176_45486.t1 bit4.t7 a_4466_45562.t1 GND.t89 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X67 a_68576_55366.t3 a_n436_44966.t31 GND.t182 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X68 a_68576_5966.t0 a_n436_5446.t18 GND.t53 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X69 a_59666_15922.t0 a_n436_5446.t19 GND.t54 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X70 OUT_N.t11 a_13666_15922.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X71 OUT_P.t9 a_4176_85006.t0 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X72 a_59666_6042.t0 a_n436_5446.t20 GND.t55 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X73 a_13376_65246.t3 bit3.t2 a_13666_65322.t3 GND.t126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X74 a_13666_6042.t1 bit5.t14 a_13376_5966.t1 GND.t226 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X75 a_40976_35606.t0 a_n436_5446.t21 GND.t56 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X76 a_68866_45562.t1 bit4.t8 a_68576_45486.t1 GND.t88 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X77 a_31776_45486.t0 a_n436_44966.t3 GND.t29 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X78 OUT_P.t10 a_50176_5966.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X79 a_41266_15922.t0 a_n436_5446.t12 GND.t30 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X80 a_50466_25802.t1 bit5.t15 a_50176_25726.t1 GND.t229 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X81 a_40976_65246.t1 bit3.t3 a_41266_65322.t2 GND.t127 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X82 OUT_P.t11 a_68576_65246.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X83 OUT_N.t12 a_4466_85082.t0 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X84 a_22866_25802.t0 a_n436_5446.t13 GND.t31 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X85 a_59376_25726.t1 bit5.t16 a_59666_25802.t0 GND.t230 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X86 a_13666_85082.t2 bit1.t0 a_13376_85006.t3 GND.t257 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X87 a_59376_65246.t3 a_n436_64726.t16 GND.t183 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X88 a_13376_5966.t3 a_n436_5446.t56 GND.t184 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X89 a_4466_15922.t2 bit5.t17 a_4176_15846.t2 GND.t212 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X90 a_22576_65246.t1 bit3.t4 a_22866_65322.t1 GND.t128 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X91 OUT_P.t12 a_40976_55366.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X92 OUT_N.t13 a_68866_65322.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X93 a_40976_45486.t3 a_n436_44966.t27 GND.t157 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X94 OUT_P.t13 a_59376_5966.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X95 a_4176_35606.t3 a_n436_5446.t44 GND.t158 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X96 OUT_P.t14 a_31776_75126.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X97 a_50466_15922.t3 a_n436_5446.t45 GND.t159 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X98 a_50176_65246.t1 bit3.t5 a_50466_65322.t2 GND.t129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X99 OUT_P.t15 a_4176_35606.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X100 OUT_P.t16 a_50176_35606.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X101 a_32066_25802.t3 a_n436_5446.t46 GND.t160 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X102 OUT_N.t14 a_59666_35682.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X103 GND.t18 bit2.t1 a_n436_74606.t3 GND.t17 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X104 a_31776_75126.t2 bit2.t2 a_32066_75202.t1 GND.t19 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X105 a_50466_6042.t3 a_n436_5446.t58 GND.t186 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X106 a_59666_45562.t1 bit4.t9 a_59376_45486.t1 GND.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X107 a_68576_25726.t2 bit5.t18 a_68866_25802.t2 GND.t213 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X108 a_4466_85082.t1 a_n436_84486.t4 GND.t187 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X109 OUT_P.t17 a_40976_5966.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X110 a_68576_65246.t3 a_n436_64726.t17 GND.t188 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X111 a_13666_35682.t3 a_n436_5446.t59 GND.t189 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X112 a_4176_55366.t1 bit4.t10 a_4466_55442.t1 GND.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X113 OUT_P.t18 a_22576_35606.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X114 OUT_P.t19 a_68576_15846.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X115 OUT_N.t15 a_32066_75202.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X116 a_41266_6042.t2 bit5.t19 a_40976_5966.t1 GND.t227 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X117 OUT_N.t16 a_50466_45562.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X118 OUT_N.t17 a_4466_35682.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X119 a_59666_25802.t2 a_n436_5446.t29 GND.t103 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X120 a_13376_75126.t1 bit2.t3 a_13666_75202.t2 GND.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X121 OUT_P.t20 a_68576_5966.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X122 OUT_P.t21 a_13376_45486.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X123 OUT_P.t22 a_59376_25726.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X124 OUT_N.t18 a_41266_55442.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X125 a_4176_45486.t2 a_n436_44966.t13 GND.t104 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X126 a_68866_55442.t2 bit4.t11 a_68576_55366.t1 GND.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X127 OUT_N.t19 a_68866_15922.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X128 a_41266_25802.t2 a_n436_5446.t30 GND.t105 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X129 OUT_N.t20 a_22866_35682.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X130 OUT_P.t23 a_31776_25726.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X131 a_68576_5966.t2 bit5.t20 a_68866_6042.t2 GND.t228 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X132 a_22866_35682.t3 a_n436_5446.t51 GND.t172 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X133 OUT_N.t21 a_13666_45562.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X134 a_13666_45562.t3 a_n436_44966.t28 GND.t173 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X135 a_4466_25802.t1 bit5.t21 a_4176_25726.t0 GND.t210 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X136 a_22576_75126.t2 bit2.t4 a_22866_75202.t1 GND.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X137 OUT_N.t22 a_32066_25802.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X138 a_50466_25802.t3 a_n436_5446.t52 GND.t174 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X139 VDD.t9 bit0.t0 a_n436_94366.t1 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X140 a_32066_35682.t3 a_n436_5446.t53 GND.t175 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X141 a_59666_55442.t2 bit4.t12 a_59376_55366.t1 GND.t84 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X142 a_4466_94962.t3 a_n436_94366.t3 GND.t176 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X143 a_13376_5966.t0 bit5.t22 a_13666_6042.t0 GND.t211 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X144 a_22866_45562.t0 a_n436_44966.t0 GND.t8 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X145 GND.t222 bit5.t23 a_n436_5446.t24 GND.t221 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X146 a_4466_15922.t0 a_n436_5446.t4 GND.t9 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X147 a_4176_65246.t2 bit3.t6 a_4466_65322.t3 GND.t130 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X148 a_59666_35682.t0 a_n436_5446.t5 GND.t10 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X149 a_68866_55442.t0 a_n436_44966.t1 GND.t11 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X150 a_31776_5966.t0 a_n436_5446.t6 GND.t12 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X151 a_68866_65322.t1 bit3.t7 a_68576_65246.t1 GND.t131 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X152 a_41266_35682.t0 a_n436_5446.t7 GND.t13 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X153 a_32066_45562.t0 a_n436_44966.t2 GND.t14 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X154 a_22866_35682.t1 bit5.t24 a_22576_35606.t0 GND.t223 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X155 a_4466_85082.t2 bit1.t1 a_4176_85006.t2 GND.t258 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X156 OUT_P.t24 a_68576_45486.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X157 a_31776_15846.t1 bit5.t25 a_32066_15922.t2 GND.t224 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X158 OUT_N.t23 a_13666_6042.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X159 a_59666_45562.t2 a_n436_44966.t10 GND.t98 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X160 OUT_P.t25 a_59376_55366.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X161 OUT_P.t26 a_4176_65246.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X162 OUT_N.t24 a_41266_6042.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X163 a_13376_15846.t0 bit5.t26 a_13666_15922.t1 GND.t217 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X164 OUT_N.t25 a_68866_45562.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X165 OUT_P.t27 a_40976_35606.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X166 OUT_P.t28 a_50176_65246.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X167 a_50466_35682.t2 a_n436_5446.t28 GND.t99 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X168 a_13376_55366.t2 a_n436_44966.t11 GND.t100 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X169 OUT_P.t29 a_31776_55366.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X170 OUT_N.t26 a_59666_65322.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X171 a_40976_5966.t0 bit5.t27 a_41266_6042.t1 GND.t218 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X172 a_41266_45562.t2 a_n436_44966.t12 GND.t101 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X173 a_32066_35682.t1 bit5.t28 a_31776_35606.t1 GND.t219 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X174 a_40976_15846.t0 bit5.t29 a_41266_15922.t1 GND.t220 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X175 a_4466_94962.t0 bit0.t1 a_4176_94886.t1 GND.t102 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X176 a_59666_65322.t2 bit3.t8 a_59376_65246.t1 GND.t132 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X177 OUT_N.t27 a_22866_6042.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X178 OUT_P.t30 a_22576_65246.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X179 OUT_N.t28 a_4466_65322.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X180 a_4466_25802.t2 a_n436_5446.t32 GND.t108 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X181 a_68866_6042.t1 bit5.t30 a_68576_5966.t1 GND.t232 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X182 a_4176_75126.t0 bit2.t5 a_4466_75202.t0 GND.t22 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X183 OUT_N.t29 a_32066_55442.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X184 OUT_P.t31 a_13376_75126.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X185 a_13666_35682.t1 bit5.t31 a_13376_35606.t1 GND.t233 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X186 OUT_N.t30 a_50466_6042.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X187 a_22576_15846.t2 bit5.t32 a_22866_15922.t1 GND.t234 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X188 a_68866_65322.t2 a_n436_64726.t7 GND.t109 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X189 a_22576_55366.t2 a_n436_44966.t15 GND.t110 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X190 OUT_N.t31 a_22866_65322.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X191 OUT_N.t32 a_41266_35682.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X192 a_50466_45562.t2 a_n436_44966.t16 GND.t111 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X193 a_41266_35682.t2 bit5.t33 a_40976_35606.t2 GND.t235 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X194 OUT_P.t32 a_4176_15846.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X195 a_50176_15846.t0 bit5.t34 a_50466_15922.t0 GND.t236 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X196 OUT_N.t33 a_32066_6042.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X197 OUT_P.t33 a_50176_15846.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X198 OUT_N.t34 a_13666_75202.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X199 a_50176_55366.t2 a_n436_44966.t17 GND.t112 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X200 a_22866_6042.t2 a_n436_5446.t33 GND.t113 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X201 a_22866_45562.t1 bit4.t13 a_22576_45486.t0 GND.t83 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X202 a_31776_25726.t0 bit5.t35 a_32066_25802.t0 GND.t237 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X203 OUT_N.t35 a_59666_15922.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X204 OUT_N.t36 a_59666_6042.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X205 OUT_N.t37 a_50466_25802.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X206 OUT_P.t34 a_22576_15846.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X207 OUT_N.t38 a_4466_15922.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X208 a_59376_15846.t2 a_n436_5446.t34 GND.t117 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X209 a_31776_55366.t2 a_n436_44966.t18 GND.t118 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X210 a_13376_25726.t0 bit5.t36 a_13666_25802.t0 GND.t190 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X211 OUT_P.t35 a_13376_25726.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X212 a_50466_35682.t1 bit5.t37 a_50176_35606.t1 GND.t191 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X213 a_13376_65246.t1 a_n436_64726.t8 GND.t119 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X214 a_59666_6042.t2 bit5.t38 a_59376_5966.t1 GND.t192 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X215 a_32066_45562.t2 bit4.t14 a_31776_45486.t2 GND.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X216 OUT_N.t39 a_22866_15922.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X217 a_40976_25726.t1 bit5.t39 a_41266_25802.t0 GND.t193 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X218 a_59376_35606.t1 bit5.t40 a_59666_35682.t1 GND.t194 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X219 OUT_P.t36 a_13376_5966.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X220 a_4466_35682.t2 a_n436_5446.t35 GND.t120 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X221 OUT_N.t40 a_13666_25802.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X222 a_68576_15846.t2 a_n436_5446.t36 GND.t121 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X223 a_40976_55366.t2 a_n436_44966.t19 GND.t122 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X224 a_13666_45562.t1 bit4.t15 a_13376_45486.t1 GND.t81 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X225 a_22576_25726.t0 bit5.t41 a_22866_25802.t1 GND.t195 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X226 a_22576_65246.t3 a_n436_64726.t10 GND.t133 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X227 a_59376_5966.t3 a_n436_5446.t37 GND.t134 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X228 GND.t260 bit1.t2 a_n436_84486.t2 GND.t259 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X229 a_41266_45562.t1 bit4.t16 a_40976_45486.t1 GND.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X230 a_50176_25726.t0 bit5.t42 a_50466_25802.t0 GND.t196 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X231 a_68576_35606.t1 bit5.t43 a_68866_35682.t1 GND.t197 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X232 OUT_N.t41 a_4466_6042.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X233 OUT_P.t37 a_22576_5966.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X234 a_50176_65246.t3 a_n436_64726.t11 GND.t135 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X235 a_22866_55442.t1 bit4.t17 a_22576_55366.t0 GND.t79 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X236 a_4466_45562.t3 a_n436_44966.t20 GND.t136 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X237 a_13376_85006.t2 bit1.t3 a_13666_85082.t1 GND.t261 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X238 a_4176_15846.t1 bit5.t44 a_4466_15922.t1 GND.t198 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X239 OUT_P.t38 a_40976_65246.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X240 a_59376_25726.t3 a_n436_5446.t38 GND.t137 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X241 OUT_P.t39 a_59376_35606.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X242 a_4176_55366.t3 a_n436_44966.t21 GND.t138 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X243 a_31776_65246.t3 a_n436_64726.t12 GND.t139 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X244 OUT_P.t40 a_4176_45486.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X245 a_50466_45562.t0 bit4.t18 a_50176_45486.t0 GND.t78 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X246 a_13376_75126.t3 a_n436_74606.t5 GND.t140 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X247 OUT_P.t41 a_50176_45486.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X248 OUT_P.t42 a_31776_5966.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X249 a_68866_15922.t1 bit5.t45 a_68576_15846.t0 GND.t199 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X250 OUT_P.t43 a_31776_35606.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X251 OUT_N.t42 a_59666_45562.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X252 VDD.t5 bit4.t19 a_n436_44966.t9 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X253 a_32066_55442.t2 bit4.t20 a_31776_55366.t0 GND.t77 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X254 a_59376_45486.t0 bit4.t21 a_59666_45562.t0 GND.t76 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X255 a_13666_55442.t0 a_n436_44966.t7 GND.t57 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X256 OUT_P.t44 a_68576_25726.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X257 a_4466_35682.t0 bit5.t46 a_4176_35606.t0 GND.t200 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X258 OUT_N.t43 a_50466_55442.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X259 OUT_P.t45 a_22576_45486.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X260 OUT_N.t44 a_4466_45562.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X261 a_68576_25726.t0 a_n436_5446.t22 GND.t58 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X262 a_41266_6042.t0 a_n436_5446.t23 GND.t59 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X263 a_4466_6042.t2 bit5.t47 a_4176_5966.t2 GND.t238 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X264 a_40976_65246.t2 a_n436_64726.t6 GND.t60 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X265 a_13666_55442.t2 bit4.t22 a_13376_55366.t0 GND.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X266 OUT_P.t46 a_13376_55366.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X267 OUT_N.t45 a_32066_35682.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X268 OUT_N.t46 a_41266_65322.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X269 a_32066_6042.t1 bit5.t48 a_31776_5966.t2 GND.t239 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X270 a_22576_75126.t0 a_n436_74606.t2 GND.t61 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X271 OUT_P.t47 a_40976_15846.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X272 GND.t115 bit0.t2 a_n436_94366.t2 GND.t114 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X273 OUT_N.t47 a_22866_45562.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X274 OUT_N.t48 a_68866_25802.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X275 a_41266_55442.t1 bit4.t23 a_40976_55366.t0 GND.t74 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X276 a_68576_45486.t0 bit4.t24 a_68866_45562.t0 GND.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X277 a_22866_55442.t0 a_n436_44966.t4 GND.t41 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X278 a_22866_65322.t0 bit3.t9 a_22576_65246.t0 GND.t32 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X279 OUT_N.t49 a_13666_55442.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X280 a_59666_15922.t1 bit5.t49 a_59376_15846.t0 GND.t240 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X281 a_4176_5966.t0 a_n436_5446.t14 GND.t42 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X282 a_4176_25726.t1 bit5.t50 a_4466_25802.t0 GND.t241 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X283 a_59376_5966.t0 bit5.t51 a_59666_6042.t1 GND.t242 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X284 a_59376_35606.t0 a_n436_5446.t15 GND.t43 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X285 a_4176_65246.t0 a_n436_64726.t3 GND.t44 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X286 a_31776_75126.t0 a_n436_74606.t1 GND.t45 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X287 a_50466_55442.t0 bit4.t25 a_50176_55366.t0 GND.t72 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X288 a_13376_85006.t0 a_n436_84486.t0 GND.t46 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X289 OUT_P.t48 a_4176_5966.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X290 a_32066_55442.t0 a_n436_44966.t5 GND.t47 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X291 OUT_N.t50 a_41266_15922.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X292 a_68866_25802.t1 bit5.t52 a_68576_25726.t1 GND.t243 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X293 a_32066_65322.t0 bit3.t10 a_31776_65246.t0 GND.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X294 a_59376_55366.t0 bit4.t26 a_59666_55442.t1 GND.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X295 a_13666_65322.t1 a_n436_64726.t4 GND.t48 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X296 a_4466_45562.t0 bit4.t27 a_4176_45486.t0 GND.t70 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X297 a_59666_55442.t0 a_n436_44966.t6 GND.t49 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X298 a_68576_35606.t0 a_n436_5446.t16 GND.t50 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X299 a_13666_65322.t0 bit3.t11 a_13376_65246.t0 GND.t34 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X300 a_59376_45486.t3 a_n436_44966.t22 GND.t142 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X301 a_68866_15922.t3 a_n436_5446.t39 GND.t143 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X302 a_41266_55442.t3 a_n436_44966.t23 GND.t144 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X303 a_41266_65322.t1 bit3.t12 a_40976_65246.t0 GND.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X304 a_68576_55366.t0 bit4.t28 a_68866_55442.t1 GND.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X305 a_22866_65322.t3 a_n436_64726.t13 GND.t145 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X306 OUT_P.t49 a_68576_55366.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X307 a_22576_5966.t3 a_n436_5446.t40 GND.t146 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X308 a_4176_85006.t3 bit1.t4 a_4466_85082.t3 GND.t262 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X309 a_22866_75202.t0 bit2.t6 a_22576_75126.t1 GND.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X310 a_59666_25802.t1 bit5.t53 a_59376_25726.t0 GND.t244 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X311 OUT_P.t50 a_59376_65246.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X312 OUT_P.t51 a_13376_85006.t1 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X313 a_68576_45486.t3 a_n436_44966.t24 GND.t147 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X314 OUT_P.t52 a_4176_75126.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X315 a_4176_75126.t3 a_n436_74606.t6 GND.t148 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X316 a_50466_55442.t3 a_n436_44966.t25 GND.t149 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X317 OUT_P.t53 a_40976_45486.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X318 OUT_N.t51 a_68866_55442.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X319 OUT_P.t54 a_31776_65246.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X320 a_50466_65322.t0 bit3.t13 a_50176_65246.t0 GND.t36 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X321 a_32066_65322.t3 a_n436_64726.t14 GND.t150 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X322 a_13376_15846.t3 a_n436_5446.t41 GND.t151 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X323 a_50466_6042.t0 bit5.t54 a_50176_5966.t1 GND.t245 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X324 OUT_N.t52 a_13666_85082.t0 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X325 a_31776_35606.t0 bit5.t55 a_32066_35682.t0 GND.t246 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X326 a_4176_5966.t1 bit5.t56 a_4466_6042.t1 GND.t247 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X327 VDD.t1 bit3.t14 a_n436_64726.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X328 a_32066_75202.t0 bit2.t7 a_31776_75126.t1 GND.t24 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X329 OUT_P.t55 a_22576_75126.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X330 a_4176_94886.t2 bit0.t3 a_4466_94962.t1 GND.t116 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X331 a_59376_65246.t0 bit3.t15 a_59666_65322.t1 GND.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X332 a_13666_75202.t0 a_n436_74606.t0 GND.t1 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X333 OUT_N.t53 a_4466_75202.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X334 a_31776_5966.t1 bit5.t57 a_32066_6042.t0 GND.t248 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X335 a_59666_65322.t0 a_n436_64726.t0 GND.t2 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X336 a_4466_55442.t0 bit4.t29 a_4176_55366.t0 GND.t68 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X337 OUT_N.t54 a_32066_65322.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X338 OUT_N.t55 a_50466_35682.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X339 a_68866_6042.t0 a_n436_5446.t0 GND.t3 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X340 a_13376_35606.t0 bit5.t58 a_13666_35682.t0 GND.t249 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X341 a_13666_75202.t1 bit2.t8 a_13376_75126.t0 GND.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X342 OUT_P.t56 a_59376_15846.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X343 OUT_N.t56 a_41266_45562.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X344 OUT_P.t57 a_13376_35606.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X345 OUT_N.t57 a_22866_75202.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X346 a_68866_25802.t0 a_n436_5446.t1 GND.t4 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X347 a_41266_65322.t0 a_n436_64726.t1 GND.t5 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X348 a_50176_5966.t0 a_n436_5446.t2 GND.t6 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X349 a_22576_15846.t0 a_n436_5446.t3 GND.t7 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X350 OUT_P.t58 a_4176_25726.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X351 a_40976_35606.t1 bit5.t59 a_41266_35682.t1 GND.t250 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X352 OUT_P.t59 a_50176_25726.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X353 a_68576_65246.t0 bit3.t16 a_68866_65322.t0 GND.t38 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X354 a_22866_75202.t3 a_n436_74606.t7 GND.t164 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X355 OUT_P.t60 a_31776_15846.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X356 OUT_N.t58 a_59666_25802.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X357 a_50176_15846.t3 a_n436_5446.t47 GND.t165 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X358 OUT_N.t59 a_13666_35682.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X359 a_22576_35606.t1 bit5.t60 a_22866_35682.t0 GND.t251 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X360 OUT_P.t61 a_22576_25726.t2 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X361 OUT_N.t60 a_4466_25802.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X362 a_13666_6042.t3 a_n436_5446.t48 GND.t166 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X363 a_4176_85006.t1 a_n436_84486.t1 GND.t167 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X364 a_50466_65322.t3 a_n436_64726.t15 GND.t168 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X365 a_31776_15846.t3 a_n436_5446.t49 GND.t169 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X366 OUT_N.t61 a_32066_15922.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X367 a_50176_35606.t0 bit5.t61 a_50466_35682.t0 GND.t252 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X368 a_22576_5966.t0 bit5.t62 a_22866_6042.t0 GND.t253 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X369 a_32066_75202.t3 a_n436_74606.t8 GND.t170 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X370 a_13376_25726.t3 a_n436_5446.t50 GND.t171 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X371 OUT_N.t62 a_22866_25802.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X372 GND.t67 bit4.t30 a_n436_44966.t8 GND.t66 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X373 a_31776_45486.t1 bit4.t31 a_32066_45562.t1 GND.t65 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X374 VDD.t7 bit2.t9 a_n436_74606.t4 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X375 a_4466_55442.t3 a_n436_44966.t32 GND.t201 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X376 a_13666_85082.t3 a_n436_84486.t5 GND.t202 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X377 a_22866_15922.t0 bit5.t63 a_22576_15846.t1 GND.t254 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X378 a_4466_65322.t0 bit3.t17 a_4176_65246.t1 GND.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X379 a_40976_5966.t3 a_n436_5446.t60 GND.t203 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X380 a_13376_45486.t0 bit4.t32 a_13666_45562.t0 GND.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X381 a_40976_15846.t3 a_n436_5446.t61 GND.t204 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X382 a_68866_35682.t3 a_n436_5446.t62 GND.t205 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X383 a_22576_25726.t3 a_n436_5446.t63 GND.t206 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
X384 a_40976_45486.t0 bit4.t33 a_41266_45562.t0 GND.t63 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X385 VDD.t11 bit1.t5 a_n436_84486.t3 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X386 a_32066_15922.t1 bit5.t64 a_31776_15846.t0 GND.t255 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X387 OUT_P.t62 a_68576_35606.t3 sky130_fd_pr__cap_mim_m3_1 l=3.3e+06u w=3.3e+06u
X388 VDD.t3 bit5.t65 a_n436_5446.t25 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3e+06u l=150000u
X389 a_50176_25726.t3 a_n436_5446.t64 GND.t207 sky130_fd_pr__res_xhigh_po_0p35 l=1e+06u
C0 VDD bit4 0.12fF
C1 VDD bit5 0.12fF
C2 VDD OUT_N 10.91fF
C3 bit0 OUT_N 26.88fF
C4 VDD OUT_P 10.88fF
C5 bit0 OUT_P 26.88fF
C6 bit1 OUT_N 26.89fF
C7 bit1 OUT_P 26.88fF
C8 bit2 OUT_N 26.89fF
C9 bit3 OUT_N 26.91fF
C10 bit2 OUT_P 26.88fF
C11 VDD bit0 0.12fF
C12 bit4 OUT_N 53.81fF
C13 bit3 OUT_P 26.88fF
C14 VDD bit1 0.12fF
C15 bit5 OUT_N 107.63fF
C16 bit4 OUT_P 53.76fF
C17 VDD bit2 0.12fF
C18 bit5 OUT_P 107.52fF
C19 VDD bit3 0.12fF
C20 OUT_N OUT_P 171.08fF
R0 bit4.n119 bit4.t19 552.693
R1 bit4.n2 bit4.t11 300.446
R2 bit4.n0 bit4.t28 300.446
R3 bit4.n9 bit4.t12 300.446
R4 bit4.n7 bit4.t26 300.446
R5 bit4.n16 bit4.t25 300.446
R6 bit4.n14 bit4.t6 300.446
R7 bit4.n23 bit4.t23 300.446
R8 bit4.n21 bit4.t4 300.446
R9 bit4.n30 bit4.t20 300.446
R10 bit4.n28 bit4.t2 300.446
R11 bit4.n37 bit4.t17 300.446
R12 bit4.n35 bit4.t5 300.446
R13 bit4.n44 bit4.t22 300.446
R14 bit4.n42 bit4.t3 300.446
R15 bit4.n53 bit4.t29 300.446
R16 bit4.n51 bit4.t10 300.446
R17 bit4.n65 bit4.t8 300.446
R18 bit4.n63 bit4.t24 300.446
R19 bit4.n72 bit4.t9 300.446
R20 bit4.n70 bit4.t21 300.446
R21 bit4.n79 bit4.t18 300.446
R22 bit4.n77 bit4.t1 300.446
R23 bit4.n86 bit4.t16 300.446
R24 bit4.n84 bit4.t33 300.446
R25 bit4.n93 bit4.t14 300.446
R26 bit4.n91 bit4.t31 300.446
R27 bit4.n100 bit4.t13 300.446
R28 bit4.n98 bit4.t0 300.446
R29 bit4.n107 bit4.t15 300.446
R30 bit4.n105 bit4.t32 300.446
R31 bit4.n114 bit4.t27 300.446
R32 bit4.n112 bit4.t7 300.446
R33 bit4.n119 bit4.t30 279.56
R34 bit4.n120 bit4.n119 120.317
R35 bit4.n52 bit4.n51 27.537
R36 bit4.n5 bit4.n2 27.536
R37 bit4.n12 bit4.n9 27.536
R38 bit4.n19 bit4.n16 27.536
R39 bit4.n26 bit4.n23 27.536
R40 bit4.n33 bit4.n30 27.536
R41 bit4.n40 bit4.n37 27.536
R42 bit4.n47 bit4.n44 27.536
R43 bit4.n68 bit4.n65 27.536
R44 bit4.n75 bit4.n72 27.536
R45 bit4.n82 bit4.n79 27.536
R46 bit4.n89 bit4.n86 27.536
R47 bit4.n96 bit4.n93 27.536
R48 bit4.n103 bit4.n100 27.536
R49 bit4.n110 bit4.n107 27.536
R50 bit4.n117 bit4.n114 27.536
R51 bit4.n1 bit4.n0 24.127
R52 bit4.n8 bit4.n7 24.127
R53 bit4.n15 bit4.n14 24.127
R54 bit4.n22 bit4.n21 24.127
R55 bit4.n29 bit4.n28 24.127
R56 bit4.n36 bit4.n35 24.127
R57 bit4.n43 bit4.n42 24.127
R58 bit4.n54 bit4.n53 24.127
R59 bit4.n64 bit4.n63 24.127
R60 bit4.n71 bit4.n70 24.127
R61 bit4.n78 bit4.n77 24.127
R62 bit4.n85 bit4.n84 24.127
R63 bit4.n92 bit4.n91 24.127
R64 bit4.n99 bit4.n98 24.127
R65 bit4.n106 bit4.n105 24.127
R66 bit4.n113 bit4.n112 24.127
R67 bit4.n4 bit4.n3 8.764
R68 bit4.n11 bit4.n10 8.764
R69 bit4.n18 bit4.n17 8.764
R70 bit4.n25 bit4.n24 8.764
R71 bit4.n32 bit4.n31 8.764
R72 bit4.n39 bit4.n38 8.764
R73 bit4.n46 bit4.n45 8.764
R74 bit4.n50 bit4.n49 8.764
R75 bit4.n67 bit4.n66 8.764
R76 bit4.n74 bit4.n73 8.764
R77 bit4.n81 bit4.n80 8.764
R78 bit4.n88 bit4.n87 8.764
R79 bit4.n95 bit4.n94 8.764
R80 bit4.n102 bit4.n101 8.764
R81 bit4.n109 bit4.n108 8.764
R82 bit4.n116 bit4.n115 8.764
R83 bit4.n6 bit4.n1 4.662
R84 bit4.n13 bit4.n8 4.662
R85 bit4.n20 bit4.n15 4.662
R86 bit4.n27 bit4.n22 4.662
R87 bit4.n34 bit4.n29 4.662
R88 bit4.n41 bit4.n36 4.662
R89 bit4.n48 bit4.n43 4.662
R90 bit4.n69 bit4.n64 4.662
R91 bit4.n76 bit4.n71 4.662
R92 bit4.n83 bit4.n78 4.662
R93 bit4.n90 bit4.n85 4.662
R94 bit4.n97 bit4.n92 4.662
R95 bit4.n104 bit4.n99 4.662
R96 bit4.n111 bit4.n106 4.662
R97 bit4.n118 bit4.n113 4.662
R98 bit4.n55 bit4.n54 4.661
R99 bit4.n5 bit4.n4 3.401
R100 bit4.n12 bit4.n11 3.401
R101 bit4.n19 bit4.n18 3.401
R102 bit4.n26 bit4.n25 3.401
R103 bit4.n33 bit4.n32 3.401
R104 bit4.n40 bit4.n39 3.401
R105 bit4.n47 bit4.n46 3.401
R106 bit4.n68 bit4.n67 3.401
R107 bit4.n75 bit4.n74 3.401
R108 bit4.n82 bit4.n81 3.401
R109 bit4.n89 bit4.n88 3.401
R110 bit4.n96 bit4.n95 3.401
R111 bit4.n103 bit4.n102 3.401
R112 bit4.n110 bit4.n109 3.401
R113 bit4.n117 bit4.n116 3.401
R114 bit4.n52 bit4.n50 3.401
R115 bit4.n128 bit4.n62 1.218
R116 bit4.n56 bit4.n55 0.873
R117 bit4.n128 bit4.n127 0.726
R118 bit4.n55 bit4.n52 0.626
R119 bit4.n6 bit4.n5 0.626
R120 bit4.n13 bit4.n12 0.626
R121 bit4.n20 bit4.n19 0.626
R122 bit4.n27 bit4.n26 0.626
R123 bit4.n34 bit4.n33 0.626
R124 bit4.n41 bit4.n40 0.626
R125 bit4.n48 bit4.n47 0.626
R126 bit4.n69 bit4.n68 0.626
R127 bit4.n76 bit4.n75 0.626
R128 bit4.n83 bit4.n82 0.626
R129 bit4.n90 bit4.n89 0.626
R130 bit4.n97 bit4.n96 0.626
R131 bit4.n104 bit4.n103 0.626
R132 bit4.n111 bit4.n110 0.626
R133 bit4.n118 bit4.n117 0.626
R134 bit4.n62 bit4.n61 0.575
R135 bit4.n61 bit4.n60 0.575
R136 bit4.n60 bit4.n59 0.575
R137 bit4.n59 bit4.n58 0.575
R138 bit4.n58 bit4.n57 0.575
R139 bit4.n57 bit4.n56 0.575
R140 bit4.n127 bit4.n126 0.575
R141 bit4.n126 bit4.n125 0.575
R142 bit4.n125 bit4.n124 0.575
R143 bit4.n124 bit4.n123 0.575
R144 bit4.n123 bit4.n122 0.575
R145 bit4.n122 bit4.n121 0.575
R146 bit4.n121 bit4.n120 0.575
R147 bit4.n62 bit4.n6 0.298
R148 bit4.n61 bit4.n13 0.298
R149 bit4.n60 bit4.n20 0.298
R150 bit4.n59 bit4.n27 0.298
R151 bit4.n58 bit4.n34 0.298
R152 bit4.n57 bit4.n41 0.298
R153 bit4.n56 bit4.n48 0.298
R154 bit4.n127 bit4.n69 0.298
R155 bit4.n126 bit4.n76 0.298
R156 bit4.n125 bit4.n83 0.298
R157 bit4.n124 bit4.n90 0.298
R158 bit4.n123 bit4.n97 0.298
R159 bit4.n122 bit4.n104 0.298
R160 bit4.n121 bit4.n111 0.298
R161 bit4.n120 bit4.n118 0.298
R162 bit4 bit4.n128 0.125
R163 a_22866_45562.n26 a_22866_45562.t1 10.181
R164 a_22866_45562.n18 a_22866_45562.t2 10.181
R165 a_22866_45562.t0 a_22866_45562.n39 9.68
R166 a_22866_45562.n3 a_22866_45562.n2 9.302
R167 a_22866_45562.n13 a_22866_45562.n12 9.302
R168 a_22866_45562.n32 a_22866_45562.n31 9.3
R169 a_22866_45562.n34 a_22866_45562.n33 9.3
R170 a_22866_45562.n7 a_22866_45562.n6 9.3
R171 a_22866_45562.n5 a_22866_45562.n4 9.3
R172 a_22866_45562.n36 a_22866_45562.n35 9
R173 a_22866_45562.n9 a_22866_45562.n8 9
R174 a_22866_45562.n27 a_22866_45562.n25 7.729
R175 a_22866_45562.n19 a_22866_45562.n17 7.729
R176 a_22866_45562.n27 a_22866_45562.n26 6.296
R177 a_22866_45562.n19 a_22866_45562.n18 6.296
R178 a_22866_45562.n30 a_22866_45562.n3 4.508
R179 a_22866_45562.n14 a_22866_45562.n13 4.508
R180 a_22866_45562.n37 a_22866_45562.n36 4.496
R181 a_22866_45562.n21 a_22866_45562.n20 4.496
R182 a_22866_45562.n29 a_22866_45562.n28 4.495
R183 a_22866_45562.n10 a_22866_45562.n9 4.495
R184 a_22866_45562.n14 a_22866_45562.n11 4.494
R185 a_22866_45562.n30 a_22866_45562.n1 4.494
R186 a_22866_45562.n39 a_22866_45562.t3 1.087
R187 a_22866_45562.n25 a_22866_45562.n24 0.536
R188 a_22866_45562.n17 a_22866_45562.n16 0.536
R189 a_22866_45562.n39 a_22866_45562.n38 0.255
R190 a_22866_45562.n28 a_22866_45562.n27 0.151
R191 a_22866_45562.n20 a_22866_45562.n19 0.151
R192 a_22866_45562.n23 a_22866_45562.n22 0.125
R193 a_22866_45562.n34 a_22866_45562.n32 0.028
R194 a_22866_45562.n7 a_22866_45562.n5 0.028
R195 a_22866_45562.n1 a_22866_45562.n0 0.025
R196 a_22866_45562.n20 a_22866_45562.n15 0.024
R197 a_22866_45562.n36 a_22866_45562.n34 0.012
R198 a_22866_45562.n9 a_22866_45562.n7 0.012
R199 a_22866_45562.n29 a_22866_45562.n23 0.011
R200 a_22866_45562.n30 a_22866_45562.n29 0.011
R201 a_22866_45562.n14 a_22866_45562.n10 0.011
R202 a_22866_45562.n38 a_22866_45562.n37 0.01
R203 a_22866_45562.n22 a_22866_45562.n21 0.01
R204 a_22866_45562.n21 a_22866_45562.n14 0.01
R205 a_22866_45562.n37 a_22866_45562.n30 0.01
R206 a_22576_45486.n10 a_22576_45486.t0 10.181
R207 a_22576_45486.n10 a_22576_45486.t1 10.181
R208 a_22576_45486.t3 a_22576_45486.n18 9.68
R209 a_22576_45486.n1 a_22576_45486.n0 9.302
R210 a_22576_45486.n7 a_22576_45486.n6 9.3
R211 a_22576_45486.n5 a_22576_45486.n4 9.3
R212 a_22576_45486.n9 a_22576_45486.n8 9
R213 a_22576_45486.n13 a_22576_45486.n12 7.729
R214 a_22576_45486.n13 a_22576_45486.n10 6.296
R215 a_22576_45486.n16 a_22576_45486.n1 4.508
R216 a_22576_45486.n15 a_22576_45486.n14 4.501
R217 a_22576_45486.n15 a_22576_45486.n9 4.501
R218 a_22576_45486.n16 a_22576_45486.n3 4.494
R219 a_22576_45486.n18 a_22576_45486.t2 1.259
R220 a_22576_45486.n12 a_22576_45486.n11 0.536
R221 a_22576_45486.n18 a_22576_45486.n17 0.415
R222 a_22576_45486.n14 a_22576_45486.n13 0.151
R223 a_22576_45486.n7 a_22576_45486.n5 0.028
R224 a_22576_45486.n3 a_22576_45486.n2 0.025
R225 a_22576_45486.n17 a_22576_45486.n16 0.021
R226 a_22576_45486.n9 a_22576_45486.n7 0.012
R227 a_22576_45486.n16 a_22576_45486.n15 0.006
R228 GND.n6 GND.t114 3941.67
R229 GND.n97 GND.t259 3941.67
R230 GND.n270 GND.t17 3941.67
R231 GND.n607 GND.t123 3941.67
R232 GND.n1927 GND.t66 3941.67
R233 GND.n4557 GND.t221 3941.67
R234 GND.n15 GND.t176 650.171
R235 GND.n55 GND.t0 650.171
R236 GND.n187 GND.t202 650.171
R237 GND.n226 GND.t46 650.171
R238 GND.n106 GND.t187 650.171
R239 GND.n145 GND.t167 650.171
R240 GND.n522 GND.t170 650.171
R241 GND.n561 GND.t45 650.171
R242 GND.n441 GND.t164 650.171
R243 GND.n480 GND.t61 650.171
R244 GND.n360 GND.t1 650.171
R245 GND.n399 GND.t140 650.171
R246 GND.n279 GND.t179 650.171
R247 GND.n318 GND.t148 650.171
R248 GND.n1183 GND.t109 650.171
R249 GND.n1222 GND.t188 650.171
R250 GND.n1102 GND.t2 650.171
R251 GND.n1141 GND.t183 650.171
R252 GND.n1021 GND.t168 650.171
R253 GND.n1060 GND.t135 650.171
R254 GND.n940 GND.t5 650.171
R255 GND.n979 GND.t60 650.171
R256 GND.n859 GND.t150 650.171
R257 GND.n898 GND.t139 650.171
R258 GND.n778 GND.t145 650.171
R259 GND.n817 GND.t133 650.171
R260 GND.n697 GND.t48 650.171
R261 GND.n736 GND.t119 650.171
R262 GND.n616 GND.t51 650.171
R263 GND.n655 GND.t44 650.171
R264 GND.n1838 GND.t11 650.171
R265 GND.n1877 GND.t182 650.171
R266 GND.n1757 GND.t49 650.171
R267 GND.n1796 GND.t177 650.171
R268 GND.n1676 GND.t149 650.171
R269 GND.n1715 GND.t112 650.171
R270 GND.n1595 GND.t144 650.171
R271 GND.n1634 GND.t122 650.171
R272 GND.n1514 GND.t47 650.171
R273 GND.n1553 GND.t118 650.171
R274 GND.n1433 GND.t41 650.171
R275 GND.n1472 GND.t110 650.171
R276 GND.n1352 GND.t57 650.171
R277 GND.n1391 GND.t100 650.171
R278 GND.n1271 GND.t201 650.171
R279 GND.n1310 GND.t138 650.171
R280 GND.n2503 GND.t256 650.171
R281 GND.n2542 GND.t147 650.171
R282 GND.n2422 GND.t98 650.171
R283 GND.n2461 GND.t142 650.171
R284 GND.n2341 GND.t111 650.171
R285 GND.n2380 GND.t180 650.171
R286 GND.n2260 GND.t101 650.171
R287 GND.n2299 GND.t157 650.171
R288 GND.n2179 GND.t14 650.171
R289 GND.n2218 GND.t29 650.171
R290 GND.n2098 GND.t8 650.171
R291 GND.n2137 GND.t153 650.171
R292 GND.n2017 GND.t173 650.171
R293 GND.n2056 GND.t106 650.171
R294 GND.n1936 GND.t136 650.171
R295 GND.n1975 GND.t104 650.171
R296 GND.n3158 GND.t205 650.171
R297 GND.n3197 GND.t50 650.171
R298 GND.n3077 GND.t10 650.171
R299 GND.n3116 GND.t43 650.171
R300 GND.n2996 GND.t99 650.171
R301 GND.n3035 GND.t185 650.171
R302 GND.n2915 GND.t13 650.171
R303 GND.n2954 GND.t56 650.171
R304 GND.n2834 GND.t175 650.171
R305 GND.n2873 GND.t152 650.171
R306 GND.n2753 GND.t172 650.171
R307 GND.n2792 GND.t97 650.171
R308 GND.n2672 GND.t189 650.171
R309 GND.n2711 GND.t263 650.171
R310 GND.n2591 GND.t120 650.171
R311 GND.n2630 GND.t158 650.171
R312 GND.n3813 GND.t4 650.171
R313 GND.n3852 GND.t58 650.171
R314 GND.n3732 GND.t103 650.171
R315 GND.n3771 GND.t137 650.171
R316 GND.n3651 GND.t174 650.171
R317 GND.n3690 GND.t207 650.171
R318 GND.n3570 GND.t105 650.171
R319 GND.n3609 GND.t28 650.171
R320 GND.n3489 GND.t160 650.171
R321 GND.n3528 GND.t154 650.171
R322 GND.n3408 GND.t31 650.171
R323 GND.n3447 GND.t206 650.171
R324 GND.n3327 GND.t181 650.171
R325 GND.n3366 GND.t171 650.171
R326 GND.n3246 GND.t108 650.171
R327 GND.n3285 GND.t178 650.171
R328 GND.n4468 GND.t143 650.171
R329 GND.n4507 GND.t121 650.171
R330 GND.n4387 GND.t54 650.171
R331 GND.n4426 GND.t117 650.171
R332 GND.n4306 GND.t159 650.171
R333 GND.n4345 GND.t165 650.171
R334 GND.n4225 GND.t30 650.171
R335 GND.n4264 GND.t204 650.171
R336 GND.n4144 GND.t52 650.171
R337 GND.n4183 GND.t169 650.171
R338 GND.n4063 GND.t107 650.171
R339 GND.n4102 GND.t7 650.171
R340 GND.n3982 GND.t26 650.171
R341 GND.n4021 GND.t151 650.171
R342 GND.n3901 GND.t9 650.171
R343 GND.n3940 GND.t15 650.171
R344 GND.n5133 GND.t3 650.171
R345 GND.n5172 GND.t53 650.171
R346 GND.n5052 GND.t55 650.171
R347 GND.n5091 GND.t134 650.171
R348 GND.n4971 GND.t186 650.171
R349 GND.n5010 GND.t6 650.171
R350 GND.n4890 GND.t59 650.171
R351 GND.n4929 GND.t203 650.171
R352 GND.n4809 GND.t62 650.171
R353 GND.n4848 GND.t12 650.171
R354 GND.n4728 GND.t113 650.171
R355 GND.n4767 GND.t146 650.171
R356 GND.n4647 GND.t166 650.171
R357 GND.n4686 GND.t184 650.171
R358 GND.n4566 GND.t27 650.171
R359 GND.n4605 GND.t42 650.171
R360 GND.n15 GND.t102 582.13
R361 GND.n55 GND.t116 582.13
R362 GND.n187 GND.t257 582.13
R363 GND.n226 GND.t261 582.13
R364 GND.n106 GND.t258 582.13
R365 GND.n145 GND.t262 582.13
R366 GND.n522 GND.t24 582.13
R367 GND.n561 GND.t19 582.13
R368 GND.n441 GND.t23 582.13
R369 GND.n480 GND.t21 582.13
R370 GND.n360 GND.t25 582.13
R371 GND.n399 GND.t20 582.13
R372 GND.n279 GND.t16 582.13
R373 GND.n318 GND.t22 582.13
R374 GND.n1183 GND.t131 582.13
R375 GND.n1222 GND.t38 582.13
R376 GND.n1102 GND.t132 582.13
R377 GND.n1141 GND.t37 582.13
R378 GND.n1021 GND.t36 582.13
R379 GND.n1060 GND.t129 582.13
R380 GND.n940 GND.t35 582.13
R381 GND.n979 GND.t127 582.13
R382 GND.n859 GND.t33 582.13
R383 GND.n898 GND.t125 582.13
R384 GND.n778 GND.t32 582.13
R385 GND.n817 GND.t128 582.13
R386 GND.n697 GND.t34 582.13
R387 GND.n736 GND.t126 582.13
R388 GND.n616 GND.t39 582.13
R389 GND.n655 GND.t130 582.13
R390 GND.n1838 GND.t85 582.13
R391 GND.n1877 GND.t69 582.13
R392 GND.n1757 GND.t84 582.13
R393 GND.n1796 GND.t71 582.13
R394 GND.n1676 GND.t72 582.13
R395 GND.n1715 GND.t90 582.13
R396 GND.n1595 GND.t74 582.13
R397 GND.n1634 GND.t92 582.13
R398 GND.n1514 GND.t77 582.13
R399 GND.n1553 GND.t94 582.13
R400 GND.n1433 GND.t79 582.13
R401 GND.n1472 GND.t91 582.13
R402 GND.n1352 GND.t75 582.13
R403 GND.n1391 GND.t93 582.13
R404 GND.n1271 GND.t68 582.13
R405 GND.n1310 GND.t86 582.13
R406 GND.n2503 GND.t88 582.13
R407 GND.n2542 GND.t73 582.13
R408 GND.n2422 GND.t87 582.13
R409 GND.n2461 GND.t76 582.13
R410 GND.n2341 GND.t78 582.13
R411 GND.n2380 GND.t95 582.13
R412 GND.n2260 GND.t80 582.13
R413 GND.n2299 GND.t63 582.13
R414 GND.n2179 GND.t82 582.13
R415 GND.n2218 GND.t65 582.13
R416 GND.n2098 GND.t83 582.13
R417 GND.n2137 GND.t96 582.13
R418 GND.n2017 GND.t81 582.13
R419 GND.n2056 GND.t64 582.13
R420 GND.n1936 GND.t70 582.13
R421 GND.n1975 GND.t89 582.13
R422 GND.n3158 GND.t231 582.13
R423 GND.n3197 GND.t197 582.13
R424 GND.n3077 GND.t215 582.13
R425 GND.n3116 GND.t194 582.13
R426 GND.n2996 GND.t191 582.13
R427 GND.n3035 GND.t252 582.13
R428 GND.n2915 GND.t235 582.13
R429 GND.n2954 GND.t250 582.13
R430 GND.n2834 GND.t219 582.13
R431 GND.n2873 GND.t246 582.13
R432 GND.n2753 GND.t223 582.13
R433 GND.n2792 GND.t251 582.13
R434 GND.n2672 GND.t233 582.13
R435 GND.n2711 GND.t249 582.13
R436 GND.n2591 GND.t200 582.13
R437 GND.n2630 GND.t163 582.13
R438 GND.n3813 GND.t243 582.13
R439 GND.n3852 GND.t213 582.13
R440 GND.n3732 GND.t244 582.13
R441 GND.n3771 GND.t230 582.13
R442 GND.n3651 GND.t229 582.13
R443 GND.n3690 GND.t196 582.13
R444 GND.n3570 GND.t214 582.13
R445 GND.n3609 GND.t193 582.13
R446 GND.n3489 GND.t209 582.13
R447 GND.n3528 GND.t237 582.13
R448 GND.n3408 GND.t216 582.13
R449 GND.n3447 GND.t195 582.13
R450 GND.n3327 GND.t40 582.13
R451 GND.n3366 GND.t190 582.13
R452 GND.n3246 GND.t210 582.13
R453 GND.n3285 GND.t241 582.13
R454 GND.n4468 GND.t199 582.13
R455 GND.n4507 GND.t225 582.13
R456 GND.n4387 GND.t240 582.13
R457 GND.n4426 GND.t155 582.13
R458 GND.n4306 GND.t162 582.13
R459 GND.n4345 GND.t236 582.13
R460 GND.n4225 GND.t156 582.13
R461 GND.n4264 GND.t220 582.13
R462 GND.n4144 GND.t255 582.13
R463 GND.n4183 GND.t224 582.13
R464 GND.n4063 GND.t254 582.13
R465 GND.n4102 GND.t234 582.13
R466 GND.n3982 GND.t208 582.13
R467 GND.n4021 GND.t217 582.13
R468 GND.n3901 GND.t212 582.13
R469 GND.n3940 GND.t198 582.13
R470 GND.n5133 GND.t232 582.13
R471 GND.n5172 GND.t228 582.13
R472 GND.n5052 GND.t192 582.13
R473 GND.n5091 GND.t242 582.13
R474 GND.n4971 GND.t245 582.13
R475 GND.n5010 GND.t161 582.13
R476 GND.n4890 GND.t227 582.13
R477 GND.n4929 GND.t218 582.13
R478 GND.n4809 GND.t239 582.13
R479 GND.n4848 GND.t248 582.13
R480 GND.n4728 GND.t141 582.13
R481 GND.n4767 GND.t253 582.13
R482 GND.n4647 GND.t226 582.13
R483 GND.n4686 GND.t211 582.13
R484 GND.n4566 GND.t238 582.13
R485 GND.n4605 GND.t247 582.13
R486 GND.n3 GND.t115 93.671
R487 GND.n94 GND.t260 93.671
R488 GND.n267 GND.t18 93.671
R489 GND.n604 GND.t124 93.671
R490 GND.n1924 GND.t67 93.671
R491 GND.n4554 GND.t222 93.671
R492 GND.n4 GND.n0 73.875
R493 GND.n95 GND.n91 73.875
R494 GND.n268 GND.n264 73.875
R495 GND.n605 GND.n601 73.875
R496 GND.n1925 GND.n1921 73.875
R497 GND.n4555 GND.n4551 73.875
R498 GND.n79 GND.n78 55.353
R499 GND.n39 GND.n38 55.353
R500 GND.n211 GND.n210 55.353
R501 GND.n130 GND.n129 55.353
R502 GND.n546 GND.n545 55.353
R503 GND.n465 GND.n464 55.353
R504 GND.n384 GND.n383 55.353
R505 GND.n303 GND.n302 55.353
R506 GND.n1207 GND.n1206 55.353
R507 GND.n1126 GND.n1125 55.353
R508 GND.n1045 GND.n1044 55.353
R509 GND.n964 GND.n963 55.353
R510 GND.n883 GND.n882 55.353
R511 GND.n802 GND.n801 55.353
R512 GND.n721 GND.n720 55.353
R513 GND.n640 GND.n639 55.353
R514 GND.n1862 GND.n1861 55.353
R515 GND.n1781 GND.n1780 55.353
R516 GND.n1700 GND.n1699 55.353
R517 GND.n1619 GND.n1618 55.353
R518 GND.n1538 GND.n1537 55.353
R519 GND.n1457 GND.n1456 55.353
R520 GND.n1376 GND.n1375 55.353
R521 GND.n1295 GND.n1294 55.353
R522 GND.n2527 GND.n2526 55.353
R523 GND.n2446 GND.n2445 55.353
R524 GND.n2365 GND.n2364 55.353
R525 GND.n2284 GND.n2283 55.353
R526 GND.n2203 GND.n2202 55.353
R527 GND.n2122 GND.n2121 55.353
R528 GND.n2041 GND.n2040 55.353
R529 GND.n1960 GND.n1959 55.353
R530 GND.n3182 GND.n3181 55.353
R531 GND.n3101 GND.n3100 55.353
R532 GND.n3020 GND.n3019 55.353
R533 GND.n2939 GND.n2938 55.353
R534 GND.n2858 GND.n2857 55.353
R535 GND.n2777 GND.n2776 55.353
R536 GND.n2696 GND.n2695 55.353
R537 GND.n2615 GND.n2614 55.353
R538 GND.n3837 GND.n3836 55.353
R539 GND.n3756 GND.n3755 55.353
R540 GND.n3675 GND.n3674 55.353
R541 GND.n3594 GND.n3593 55.353
R542 GND.n3513 GND.n3512 55.353
R543 GND.n3432 GND.n3431 55.353
R544 GND.n3351 GND.n3350 55.353
R545 GND.n3270 GND.n3269 55.353
R546 GND.n4492 GND.n4491 55.353
R547 GND.n4411 GND.n4410 55.353
R548 GND.n4330 GND.n4329 55.353
R549 GND.n4249 GND.n4248 55.353
R550 GND.n4168 GND.n4167 55.353
R551 GND.n4087 GND.n4086 55.353
R552 GND.n4006 GND.n4005 55.353
R553 GND.n3925 GND.n3924 55.353
R554 GND.n5157 GND.n5156 55.353
R555 GND.n5076 GND.n5075 55.353
R556 GND.n4995 GND.n4994 55.353
R557 GND.n4914 GND.n4913 55.353
R558 GND.n4833 GND.n4832 55.353
R559 GND.n4752 GND.n4751 55.353
R560 GND.n4671 GND.n4670 55.353
R561 GND.n4590 GND.n4589 55.353
R562 GND.n71 GND.n70 54.344
R563 GND.n80 GND.n79 54.344
R564 GND.n31 GND.n30 54.344
R565 GND.n40 GND.n39 54.344
R566 GND.n243 GND.n242 54.344
R567 GND.n203 GND.n202 54.344
R568 GND.n212 GND.n211 54.344
R569 GND.n162 GND.n161 54.344
R570 GND.n122 GND.n121 54.344
R571 GND.n131 GND.n130 54.344
R572 GND.n578 GND.n577 54.344
R573 GND.n538 GND.n537 54.344
R574 GND.n547 GND.n546 54.344
R575 GND.n497 GND.n496 54.344
R576 GND.n457 GND.n456 54.344
R577 GND.n466 GND.n465 54.344
R578 GND.n416 GND.n415 54.344
R579 GND.n376 GND.n375 54.344
R580 GND.n385 GND.n384 54.344
R581 GND.n335 GND.n334 54.344
R582 GND.n295 GND.n294 54.344
R583 GND.n304 GND.n303 54.344
R584 GND.n1239 GND.n1238 54.344
R585 GND.n1199 GND.n1198 54.344
R586 GND.n1208 GND.n1207 54.344
R587 GND.n1158 GND.n1157 54.344
R588 GND.n1118 GND.n1117 54.344
R589 GND.n1127 GND.n1126 54.344
R590 GND.n1077 GND.n1076 54.344
R591 GND.n1037 GND.n1036 54.344
R592 GND.n1046 GND.n1045 54.344
R593 GND.n996 GND.n995 54.344
R594 GND.n956 GND.n955 54.344
R595 GND.n965 GND.n964 54.344
R596 GND.n915 GND.n914 54.344
R597 GND.n875 GND.n874 54.344
R598 GND.n884 GND.n883 54.344
R599 GND.n834 GND.n833 54.344
R600 GND.n794 GND.n793 54.344
R601 GND.n803 GND.n802 54.344
R602 GND.n753 GND.n752 54.344
R603 GND.n713 GND.n712 54.344
R604 GND.n722 GND.n721 54.344
R605 GND.n672 GND.n671 54.344
R606 GND.n632 GND.n631 54.344
R607 GND.n641 GND.n640 54.344
R608 GND.n1894 GND.n1893 54.344
R609 GND.n1854 GND.n1853 54.344
R610 GND.n1863 GND.n1862 54.344
R611 GND.n1813 GND.n1812 54.344
R612 GND.n1773 GND.n1772 54.344
R613 GND.n1782 GND.n1781 54.344
R614 GND.n1732 GND.n1731 54.344
R615 GND.n1692 GND.n1691 54.344
R616 GND.n1701 GND.n1700 54.344
R617 GND.n1651 GND.n1650 54.344
R618 GND.n1611 GND.n1610 54.344
R619 GND.n1620 GND.n1619 54.344
R620 GND.n1570 GND.n1569 54.344
R621 GND.n1530 GND.n1529 54.344
R622 GND.n1539 GND.n1538 54.344
R623 GND.n1489 GND.n1488 54.344
R624 GND.n1449 GND.n1448 54.344
R625 GND.n1458 GND.n1457 54.344
R626 GND.n1408 GND.n1407 54.344
R627 GND.n1368 GND.n1367 54.344
R628 GND.n1377 GND.n1376 54.344
R629 GND.n1327 GND.n1326 54.344
R630 GND.n1287 GND.n1286 54.344
R631 GND.n1296 GND.n1295 54.344
R632 GND.n2559 GND.n2558 54.344
R633 GND.n2519 GND.n2518 54.344
R634 GND.n2528 GND.n2527 54.344
R635 GND.n2478 GND.n2477 54.344
R636 GND.n2438 GND.n2437 54.344
R637 GND.n2447 GND.n2446 54.344
R638 GND.n2397 GND.n2396 54.344
R639 GND.n2357 GND.n2356 54.344
R640 GND.n2366 GND.n2365 54.344
R641 GND.n2316 GND.n2315 54.344
R642 GND.n2276 GND.n2275 54.344
R643 GND.n2285 GND.n2284 54.344
R644 GND.n2235 GND.n2234 54.344
R645 GND.n2195 GND.n2194 54.344
R646 GND.n2204 GND.n2203 54.344
R647 GND.n2154 GND.n2153 54.344
R648 GND.n2114 GND.n2113 54.344
R649 GND.n2123 GND.n2122 54.344
R650 GND.n2073 GND.n2072 54.344
R651 GND.n2033 GND.n2032 54.344
R652 GND.n2042 GND.n2041 54.344
R653 GND.n1992 GND.n1991 54.344
R654 GND.n1952 GND.n1951 54.344
R655 GND.n1961 GND.n1960 54.344
R656 GND.n3214 GND.n3213 54.344
R657 GND.n3174 GND.n3173 54.344
R658 GND.n3183 GND.n3182 54.344
R659 GND.n3133 GND.n3132 54.344
R660 GND.n3093 GND.n3092 54.344
R661 GND.n3102 GND.n3101 54.344
R662 GND.n3052 GND.n3051 54.344
R663 GND.n3012 GND.n3011 54.344
R664 GND.n3021 GND.n3020 54.344
R665 GND.n2971 GND.n2970 54.344
R666 GND.n2931 GND.n2930 54.344
R667 GND.n2940 GND.n2939 54.344
R668 GND.n2890 GND.n2889 54.344
R669 GND.n2850 GND.n2849 54.344
R670 GND.n2859 GND.n2858 54.344
R671 GND.n2809 GND.n2808 54.344
R672 GND.n2769 GND.n2768 54.344
R673 GND.n2778 GND.n2777 54.344
R674 GND.n2728 GND.n2727 54.344
R675 GND.n2688 GND.n2687 54.344
R676 GND.n2697 GND.n2696 54.344
R677 GND.n2647 GND.n2646 54.344
R678 GND.n2607 GND.n2606 54.344
R679 GND.n2616 GND.n2615 54.344
R680 GND.n3869 GND.n3868 54.344
R681 GND.n3829 GND.n3828 54.344
R682 GND.n3838 GND.n3837 54.344
R683 GND.n3788 GND.n3787 54.344
R684 GND.n3748 GND.n3747 54.344
R685 GND.n3757 GND.n3756 54.344
R686 GND.n3707 GND.n3706 54.344
R687 GND.n3667 GND.n3666 54.344
R688 GND.n3676 GND.n3675 54.344
R689 GND.n3626 GND.n3625 54.344
R690 GND.n3586 GND.n3585 54.344
R691 GND.n3595 GND.n3594 54.344
R692 GND.n3545 GND.n3544 54.344
R693 GND.n3505 GND.n3504 54.344
R694 GND.n3514 GND.n3513 54.344
R695 GND.n3464 GND.n3463 54.344
R696 GND.n3424 GND.n3423 54.344
R697 GND.n3433 GND.n3432 54.344
R698 GND.n3383 GND.n3382 54.344
R699 GND.n3343 GND.n3342 54.344
R700 GND.n3352 GND.n3351 54.344
R701 GND.n3302 GND.n3301 54.344
R702 GND.n3262 GND.n3261 54.344
R703 GND.n3271 GND.n3270 54.344
R704 GND.n4524 GND.n4523 54.344
R705 GND.n4484 GND.n4483 54.344
R706 GND.n4493 GND.n4492 54.344
R707 GND.n4443 GND.n4442 54.344
R708 GND.n4403 GND.n4402 54.344
R709 GND.n4412 GND.n4411 54.344
R710 GND.n4362 GND.n4361 54.344
R711 GND.n4322 GND.n4321 54.344
R712 GND.n4331 GND.n4330 54.344
R713 GND.n4281 GND.n4280 54.344
R714 GND.n4241 GND.n4240 54.344
R715 GND.n4250 GND.n4249 54.344
R716 GND.n4200 GND.n4199 54.344
R717 GND.n4160 GND.n4159 54.344
R718 GND.n4169 GND.n4168 54.344
R719 GND.n4119 GND.n4118 54.344
R720 GND.n4079 GND.n4078 54.344
R721 GND.n4088 GND.n4087 54.344
R722 GND.n4038 GND.n4037 54.344
R723 GND.n3998 GND.n3997 54.344
R724 GND.n4007 GND.n4006 54.344
R725 GND.n3957 GND.n3956 54.344
R726 GND.n3917 GND.n3916 54.344
R727 GND.n3926 GND.n3925 54.344
R728 GND.n5189 GND.n5188 54.344
R729 GND.n5149 GND.n5148 54.344
R730 GND.n5158 GND.n5157 54.344
R731 GND.n5108 GND.n5107 54.344
R732 GND.n5068 GND.n5067 54.344
R733 GND.n5077 GND.n5076 54.344
R734 GND.n5027 GND.n5026 54.344
R735 GND.n4987 GND.n4986 54.344
R736 GND.n4996 GND.n4995 54.344
R737 GND.n4946 GND.n4945 54.344
R738 GND.n4906 GND.n4905 54.344
R739 GND.n4915 GND.n4914 54.344
R740 GND.n4865 GND.n4864 54.344
R741 GND.n4825 GND.n4824 54.344
R742 GND.n4834 GND.n4833 54.344
R743 GND.n4784 GND.n4783 54.344
R744 GND.n4744 GND.n4743 54.344
R745 GND.n4753 GND.n4752 54.344
R746 GND.n4703 GND.n4702 54.344
R747 GND.n4663 GND.n4662 54.344
R748 GND.n4672 GND.n4671 54.344
R749 GND.n4622 GND.n4621 54.344
R750 GND.n4582 GND.n4581 54.344
R751 GND.n4591 GND.n4590 54.344
R752 GND.n61 GND.n60 47.551
R753 GND.n21 GND.n20 47.551
R754 GND.n225 GND.n224 47.551
R755 GND.n193 GND.n192 47.551
R756 GND.n144 GND.n143 47.551
R757 GND.n112 GND.n111 47.551
R758 GND.n560 GND.n559 47.551
R759 GND.n528 GND.n527 47.551
R760 GND.n479 GND.n478 47.551
R761 GND.n447 GND.n446 47.551
R762 GND.n398 GND.n397 47.551
R763 GND.n366 GND.n365 47.551
R764 GND.n317 GND.n316 47.551
R765 GND.n285 GND.n284 47.551
R766 GND.n1221 GND.n1220 47.551
R767 GND.n1189 GND.n1188 47.551
R768 GND.n1140 GND.n1139 47.551
R769 GND.n1108 GND.n1107 47.551
R770 GND.n1059 GND.n1058 47.551
R771 GND.n1027 GND.n1026 47.551
R772 GND.n978 GND.n977 47.551
R773 GND.n946 GND.n945 47.551
R774 GND.n897 GND.n896 47.551
R775 GND.n865 GND.n864 47.551
R776 GND.n816 GND.n815 47.551
R777 GND.n784 GND.n783 47.551
R778 GND.n735 GND.n734 47.551
R779 GND.n703 GND.n702 47.551
R780 GND.n654 GND.n653 47.551
R781 GND.n622 GND.n621 47.551
R782 GND.n1876 GND.n1875 47.551
R783 GND.n1844 GND.n1843 47.551
R784 GND.n1795 GND.n1794 47.551
R785 GND.n1763 GND.n1762 47.551
R786 GND.n1714 GND.n1713 47.551
R787 GND.n1682 GND.n1681 47.551
R788 GND.n1633 GND.n1632 47.551
R789 GND.n1601 GND.n1600 47.551
R790 GND.n1552 GND.n1551 47.551
R791 GND.n1520 GND.n1519 47.551
R792 GND.n1471 GND.n1470 47.551
R793 GND.n1439 GND.n1438 47.551
R794 GND.n1390 GND.n1389 47.551
R795 GND.n1358 GND.n1357 47.551
R796 GND.n1309 GND.n1308 47.551
R797 GND.n1277 GND.n1276 47.551
R798 GND.n2541 GND.n2540 47.551
R799 GND.n2509 GND.n2508 47.551
R800 GND.n2460 GND.n2459 47.551
R801 GND.n2428 GND.n2427 47.551
R802 GND.n2379 GND.n2378 47.551
R803 GND.n2347 GND.n2346 47.551
R804 GND.n2298 GND.n2297 47.551
R805 GND.n2266 GND.n2265 47.551
R806 GND.n2217 GND.n2216 47.551
R807 GND.n2185 GND.n2184 47.551
R808 GND.n2136 GND.n2135 47.551
R809 GND.n2104 GND.n2103 47.551
R810 GND.n2055 GND.n2054 47.551
R811 GND.n2023 GND.n2022 47.551
R812 GND.n1974 GND.n1973 47.551
R813 GND.n1942 GND.n1941 47.551
R814 GND.n3196 GND.n3195 47.551
R815 GND.n3164 GND.n3163 47.551
R816 GND.n3115 GND.n3114 47.551
R817 GND.n3083 GND.n3082 47.551
R818 GND.n3034 GND.n3033 47.551
R819 GND.n3002 GND.n3001 47.551
R820 GND.n2953 GND.n2952 47.551
R821 GND.n2921 GND.n2920 47.551
R822 GND.n2872 GND.n2871 47.551
R823 GND.n2840 GND.n2839 47.551
R824 GND.n2791 GND.n2790 47.551
R825 GND.n2759 GND.n2758 47.551
R826 GND.n2710 GND.n2709 47.551
R827 GND.n2678 GND.n2677 47.551
R828 GND.n2629 GND.n2628 47.551
R829 GND.n2597 GND.n2596 47.551
R830 GND.n3851 GND.n3850 47.551
R831 GND.n3819 GND.n3818 47.551
R832 GND.n3770 GND.n3769 47.551
R833 GND.n3738 GND.n3737 47.551
R834 GND.n3689 GND.n3688 47.551
R835 GND.n3657 GND.n3656 47.551
R836 GND.n3608 GND.n3607 47.551
R837 GND.n3576 GND.n3575 47.551
R838 GND.n3527 GND.n3526 47.551
R839 GND.n3495 GND.n3494 47.551
R840 GND.n3446 GND.n3445 47.551
R841 GND.n3414 GND.n3413 47.551
R842 GND.n3365 GND.n3364 47.551
R843 GND.n3333 GND.n3332 47.551
R844 GND.n3284 GND.n3283 47.551
R845 GND.n3252 GND.n3251 47.551
R846 GND.n4506 GND.n4505 47.551
R847 GND.n4474 GND.n4473 47.551
R848 GND.n4425 GND.n4424 47.551
R849 GND.n4393 GND.n4392 47.551
R850 GND.n4344 GND.n4343 47.551
R851 GND.n4312 GND.n4311 47.551
R852 GND.n4263 GND.n4262 47.551
R853 GND.n4231 GND.n4230 47.551
R854 GND.n4182 GND.n4181 47.551
R855 GND.n4150 GND.n4149 47.551
R856 GND.n4101 GND.n4100 47.551
R857 GND.n4069 GND.n4068 47.551
R858 GND.n4020 GND.n4019 47.551
R859 GND.n3988 GND.n3987 47.551
R860 GND.n3939 GND.n3938 47.551
R861 GND.n3907 GND.n3906 47.551
R862 GND.n5171 GND.n5170 47.551
R863 GND.n5139 GND.n5138 47.551
R864 GND.n5090 GND.n5089 47.551
R865 GND.n5058 GND.n5057 47.551
R866 GND.n5009 GND.n5008 47.551
R867 GND.n4977 GND.n4976 47.551
R868 GND.n4928 GND.n4927 47.551
R869 GND.n4896 GND.n4895 47.551
R870 GND.n4847 GND.n4846 47.551
R871 GND.n4815 GND.n4814 47.551
R872 GND.n4766 GND.n4765 47.551
R873 GND.n4734 GND.n4733 47.551
R874 GND.n4685 GND.n4684 47.551
R875 GND.n4653 GND.n4652 47.551
R876 GND.n4604 GND.n4603 47.551
R877 GND.n4572 GND.n4571 47.551
R878 GND.n252 GND.n251 25.966
R879 GND.n251 GND.n250 25.966
R880 GND.n171 GND.n170 25.966
R881 GND.n170 GND.n169 25.966
R882 GND.n587 GND.n586 25.966
R883 GND.n586 GND.n585 25.966
R884 GND.n506 GND.n505 25.966
R885 GND.n505 GND.n504 25.966
R886 GND.n425 GND.n424 25.966
R887 GND.n424 GND.n423 25.966
R888 GND.n344 GND.n343 25.966
R889 GND.n343 GND.n342 25.966
R890 GND.n1248 GND.n1247 25.966
R891 GND.n1247 GND.n1246 25.966
R892 GND.n1167 GND.n1166 25.966
R893 GND.n1166 GND.n1165 25.966
R894 GND.n1086 GND.n1085 25.966
R895 GND.n1085 GND.n1084 25.966
R896 GND.n1005 GND.n1004 25.966
R897 GND.n1004 GND.n1003 25.966
R898 GND.n924 GND.n923 25.966
R899 GND.n923 GND.n922 25.966
R900 GND.n843 GND.n842 25.966
R901 GND.n842 GND.n841 25.966
R902 GND.n762 GND.n761 25.966
R903 GND.n761 GND.n760 25.966
R904 GND.n681 GND.n680 25.966
R905 GND.n680 GND.n679 25.966
R906 GND.n1903 GND.n1902 25.966
R907 GND.n1902 GND.n1901 25.966
R908 GND.n1822 GND.n1821 25.966
R909 GND.n1821 GND.n1820 25.966
R910 GND.n1741 GND.n1740 25.966
R911 GND.n1740 GND.n1739 25.966
R912 GND.n1660 GND.n1659 25.966
R913 GND.n1659 GND.n1658 25.966
R914 GND.n1579 GND.n1578 25.966
R915 GND.n1578 GND.n1577 25.966
R916 GND.n1498 GND.n1497 25.966
R917 GND.n1497 GND.n1496 25.966
R918 GND.n1417 GND.n1416 25.966
R919 GND.n1416 GND.n1415 25.966
R920 GND.n1336 GND.n1335 25.966
R921 GND.n1335 GND.n1334 25.966
R922 GND.n2568 GND.n2567 25.966
R923 GND.n2567 GND.n2566 25.966
R924 GND.n2487 GND.n2486 25.966
R925 GND.n2486 GND.n2485 25.966
R926 GND.n2406 GND.n2405 25.966
R927 GND.n2405 GND.n2404 25.966
R928 GND.n2325 GND.n2324 25.966
R929 GND.n2324 GND.n2323 25.966
R930 GND.n2244 GND.n2243 25.966
R931 GND.n2243 GND.n2242 25.966
R932 GND.n2163 GND.n2162 25.966
R933 GND.n2162 GND.n2161 25.966
R934 GND.n2082 GND.n2081 25.966
R935 GND.n2081 GND.n2080 25.966
R936 GND.n2001 GND.n2000 25.966
R937 GND.n2000 GND.n1999 25.966
R938 GND.n3223 GND.n3222 25.966
R939 GND.n3222 GND.n3221 25.966
R940 GND.n3142 GND.n3141 25.966
R941 GND.n3141 GND.n3140 25.966
R942 GND.n3061 GND.n3060 25.966
R943 GND.n3060 GND.n3059 25.966
R944 GND.n2980 GND.n2979 25.966
R945 GND.n2979 GND.n2978 25.966
R946 GND.n2899 GND.n2898 25.966
R947 GND.n2898 GND.n2897 25.966
R948 GND.n2818 GND.n2817 25.966
R949 GND.n2817 GND.n2816 25.966
R950 GND.n2737 GND.n2736 25.966
R951 GND.n2736 GND.n2735 25.966
R952 GND.n2656 GND.n2655 25.966
R953 GND.n2655 GND.n2654 25.966
R954 GND.n3878 GND.n3877 25.966
R955 GND.n3877 GND.n3876 25.966
R956 GND.n3797 GND.n3796 25.966
R957 GND.n3796 GND.n3795 25.966
R958 GND.n3716 GND.n3715 25.966
R959 GND.n3715 GND.n3714 25.966
R960 GND.n3635 GND.n3634 25.966
R961 GND.n3634 GND.n3633 25.966
R962 GND.n3554 GND.n3553 25.966
R963 GND.n3553 GND.n3552 25.966
R964 GND.n3473 GND.n3472 25.966
R965 GND.n3472 GND.n3471 25.966
R966 GND.n3392 GND.n3391 25.966
R967 GND.n3391 GND.n3390 25.966
R968 GND.n3311 GND.n3310 25.966
R969 GND.n3310 GND.n3309 25.966
R970 GND.n4533 GND.n4532 25.966
R971 GND.n4532 GND.n4531 25.966
R972 GND.n4452 GND.n4451 25.966
R973 GND.n4451 GND.n4450 25.966
R974 GND.n4371 GND.n4370 25.966
R975 GND.n4370 GND.n4369 25.966
R976 GND.n4290 GND.n4289 25.966
R977 GND.n4289 GND.n4288 25.966
R978 GND.n4209 GND.n4208 25.966
R979 GND.n4208 GND.n4207 25.966
R980 GND.n4128 GND.n4127 25.966
R981 GND.n4127 GND.n4126 25.966
R982 GND.n4047 GND.n4046 25.966
R983 GND.n4046 GND.n4045 25.966
R984 GND.n3966 GND.n3965 25.966
R985 GND.n3965 GND.n3964 25.966
R986 GND.n5198 GND.n5197 25.966
R987 GND.n5197 GND.n5196 25.966
R988 GND.n5117 GND.n5116 25.966
R989 GND.n5116 GND.n5115 25.966
R990 GND.n5036 GND.n5035 25.966
R991 GND.n5035 GND.n5034 25.966
R992 GND.n4955 GND.n4954 25.966
R993 GND.n4954 GND.n4953 25.966
R994 GND.n4874 GND.n4873 25.966
R995 GND.n4873 GND.n4872 25.966
R996 GND.n4793 GND.n4792 25.966
R997 GND.n4792 GND.n4791 25.966
R998 GND.n4712 GND.n4711 25.966
R999 GND.n4711 GND.n4710 25.966
R1000 GND.n4631 GND.n4630 25.966
R1001 GND.n4630 GND.n4629 25.966
R1002 GND.n53 GND.n52 22.848
R1003 GND.n54 GND.n53 22.848
R1004 GND.n13 GND.n12 22.848
R1005 GND.n14 GND.n13 22.848
R1006 GND.n232 GND.n231 22.848
R1007 GND.n233 GND.n232 22.848
R1008 GND.n185 GND.n184 22.848
R1009 GND.n186 GND.n185 22.848
R1010 GND.n151 GND.n150 22.848
R1011 GND.n152 GND.n151 22.848
R1012 GND.n104 GND.n103 22.848
R1013 GND.n105 GND.n104 22.848
R1014 GND.n567 GND.n566 22.848
R1015 GND.n568 GND.n567 22.848
R1016 GND.n520 GND.n519 22.848
R1017 GND.n521 GND.n520 22.848
R1018 GND.n486 GND.n485 22.848
R1019 GND.n487 GND.n486 22.848
R1020 GND.n439 GND.n438 22.848
R1021 GND.n440 GND.n439 22.848
R1022 GND.n405 GND.n404 22.848
R1023 GND.n406 GND.n405 22.848
R1024 GND.n358 GND.n357 22.848
R1025 GND.n359 GND.n358 22.848
R1026 GND.n324 GND.n323 22.848
R1027 GND.n325 GND.n324 22.848
R1028 GND.n277 GND.n276 22.848
R1029 GND.n278 GND.n277 22.848
R1030 GND.n1228 GND.n1227 22.848
R1031 GND.n1229 GND.n1228 22.848
R1032 GND.n1181 GND.n1180 22.848
R1033 GND.n1182 GND.n1181 22.848
R1034 GND.n1147 GND.n1146 22.848
R1035 GND.n1148 GND.n1147 22.848
R1036 GND.n1100 GND.n1099 22.848
R1037 GND.n1101 GND.n1100 22.848
R1038 GND.n1066 GND.n1065 22.848
R1039 GND.n1067 GND.n1066 22.848
R1040 GND.n1019 GND.n1018 22.848
R1041 GND.n1020 GND.n1019 22.848
R1042 GND.n985 GND.n984 22.848
R1043 GND.n986 GND.n985 22.848
R1044 GND.n938 GND.n937 22.848
R1045 GND.n939 GND.n938 22.848
R1046 GND.n904 GND.n903 22.848
R1047 GND.n905 GND.n904 22.848
R1048 GND.n857 GND.n856 22.848
R1049 GND.n858 GND.n857 22.848
R1050 GND.n823 GND.n822 22.848
R1051 GND.n824 GND.n823 22.848
R1052 GND.n776 GND.n775 22.848
R1053 GND.n777 GND.n776 22.848
R1054 GND.n742 GND.n741 22.848
R1055 GND.n743 GND.n742 22.848
R1056 GND.n695 GND.n694 22.848
R1057 GND.n696 GND.n695 22.848
R1058 GND.n661 GND.n660 22.848
R1059 GND.n662 GND.n661 22.848
R1060 GND.n614 GND.n613 22.848
R1061 GND.n615 GND.n614 22.848
R1062 GND.n1883 GND.n1882 22.848
R1063 GND.n1884 GND.n1883 22.848
R1064 GND.n1836 GND.n1835 22.848
R1065 GND.n1837 GND.n1836 22.848
R1066 GND.n1802 GND.n1801 22.848
R1067 GND.n1803 GND.n1802 22.848
R1068 GND.n1755 GND.n1754 22.848
R1069 GND.n1756 GND.n1755 22.848
R1070 GND.n1721 GND.n1720 22.848
R1071 GND.n1722 GND.n1721 22.848
R1072 GND.n1674 GND.n1673 22.848
R1073 GND.n1675 GND.n1674 22.848
R1074 GND.n1640 GND.n1639 22.848
R1075 GND.n1641 GND.n1640 22.848
R1076 GND.n1593 GND.n1592 22.848
R1077 GND.n1594 GND.n1593 22.848
R1078 GND.n1559 GND.n1558 22.848
R1079 GND.n1560 GND.n1559 22.848
R1080 GND.n1512 GND.n1511 22.848
R1081 GND.n1513 GND.n1512 22.848
R1082 GND.n1478 GND.n1477 22.848
R1083 GND.n1479 GND.n1478 22.848
R1084 GND.n1431 GND.n1430 22.848
R1085 GND.n1432 GND.n1431 22.848
R1086 GND.n1397 GND.n1396 22.848
R1087 GND.n1398 GND.n1397 22.848
R1088 GND.n1350 GND.n1349 22.848
R1089 GND.n1351 GND.n1350 22.848
R1090 GND.n1316 GND.n1315 22.848
R1091 GND.n1317 GND.n1316 22.848
R1092 GND.n1269 GND.n1268 22.848
R1093 GND.n1270 GND.n1269 22.848
R1094 GND.n2548 GND.n2547 22.848
R1095 GND.n2549 GND.n2548 22.848
R1096 GND.n2501 GND.n2500 22.848
R1097 GND.n2502 GND.n2501 22.848
R1098 GND.n2467 GND.n2466 22.848
R1099 GND.n2468 GND.n2467 22.848
R1100 GND.n2420 GND.n2419 22.848
R1101 GND.n2421 GND.n2420 22.848
R1102 GND.n2386 GND.n2385 22.848
R1103 GND.n2387 GND.n2386 22.848
R1104 GND.n2339 GND.n2338 22.848
R1105 GND.n2340 GND.n2339 22.848
R1106 GND.n2305 GND.n2304 22.848
R1107 GND.n2306 GND.n2305 22.848
R1108 GND.n2258 GND.n2257 22.848
R1109 GND.n2259 GND.n2258 22.848
R1110 GND.n2224 GND.n2223 22.848
R1111 GND.n2225 GND.n2224 22.848
R1112 GND.n2177 GND.n2176 22.848
R1113 GND.n2178 GND.n2177 22.848
R1114 GND.n2143 GND.n2142 22.848
R1115 GND.n2144 GND.n2143 22.848
R1116 GND.n2096 GND.n2095 22.848
R1117 GND.n2097 GND.n2096 22.848
R1118 GND.n2062 GND.n2061 22.848
R1119 GND.n2063 GND.n2062 22.848
R1120 GND.n2015 GND.n2014 22.848
R1121 GND.n2016 GND.n2015 22.848
R1122 GND.n1981 GND.n1980 22.848
R1123 GND.n1982 GND.n1981 22.848
R1124 GND.n1934 GND.n1933 22.848
R1125 GND.n1935 GND.n1934 22.848
R1126 GND.n3203 GND.n3202 22.848
R1127 GND.n3204 GND.n3203 22.848
R1128 GND.n3156 GND.n3155 22.848
R1129 GND.n3157 GND.n3156 22.848
R1130 GND.n3122 GND.n3121 22.848
R1131 GND.n3123 GND.n3122 22.848
R1132 GND.n3075 GND.n3074 22.848
R1133 GND.n3076 GND.n3075 22.848
R1134 GND.n3041 GND.n3040 22.848
R1135 GND.n3042 GND.n3041 22.848
R1136 GND.n2994 GND.n2993 22.848
R1137 GND.n2995 GND.n2994 22.848
R1138 GND.n2960 GND.n2959 22.848
R1139 GND.n2961 GND.n2960 22.848
R1140 GND.n2913 GND.n2912 22.848
R1141 GND.n2914 GND.n2913 22.848
R1142 GND.n2879 GND.n2878 22.848
R1143 GND.n2880 GND.n2879 22.848
R1144 GND.n2832 GND.n2831 22.848
R1145 GND.n2833 GND.n2832 22.848
R1146 GND.n2798 GND.n2797 22.848
R1147 GND.n2799 GND.n2798 22.848
R1148 GND.n2751 GND.n2750 22.848
R1149 GND.n2752 GND.n2751 22.848
R1150 GND.n2717 GND.n2716 22.848
R1151 GND.n2718 GND.n2717 22.848
R1152 GND.n2670 GND.n2669 22.848
R1153 GND.n2671 GND.n2670 22.848
R1154 GND.n2636 GND.n2635 22.848
R1155 GND.n2637 GND.n2636 22.848
R1156 GND.n2589 GND.n2588 22.848
R1157 GND.n2590 GND.n2589 22.848
R1158 GND.n3858 GND.n3857 22.848
R1159 GND.n3859 GND.n3858 22.848
R1160 GND.n3811 GND.n3810 22.848
R1161 GND.n3812 GND.n3811 22.848
R1162 GND.n3777 GND.n3776 22.848
R1163 GND.n3778 GND.n3777 22.848
R1164 GND.n3730 GND.n3729 22.848
R1165 GND.n3731 GND.n3730 22.848
R1166 GND.n3696 GND.n3695 22.848
R1167 GND.n3697 GND.n3696 22.848
R1168 GND.n3649 GND.n3648 22.848
R1169 GND.n3650 GND.n3649 22.848
R1170 GND.n3615 GND.n3614 22.848
R1171 GND.n3616 GND.n3615 22.848
R1172 GND.n3568 GND.n3567 22.848
R1173 GND.n3569 GND.n3568 22.848
R1174 GND.n3534 GND.n3533 22.848
R1175 GND.n3535 GND.n3534 22.848
R1176 GND.n3487 GND.n3486 22.848
R1177 GND.n3488 GND.n3487 22.848
R1178 GND.n3453 GND.n3452 22.848
R1179 GND.n3454 GND.n3453 22.848
R1180 GND.n3406 GND.n3405 22.848
R1181 GND.n3407 GND.n3406 22.848
R1182 GND.n3372 GND.n3371 22.848
R1183 GND.n3373 GND.n3372 22.848
R1184 GND.n3325 GND.n3324 22.848
R1185 GND.n3326 GND.n3325 22.848
R1186 GND.n3291 GND.n3290 22.848
R1187 GND.n3292 GND.n3291 22.848
R1188 GND.n3244 GND.n3243 22.848
R1189 GND.n3245 GND.n3244 22.848
R1190 GND.n4513 GND.n4512 22.848
R1191 GND.n4514 GND.n4513 22.848
R1192 GND.n4466 GND.n4465 22.848
R1193 GND.n4467 GND.n4466 22.848
R1194 GND.n4432 GND.n4431 22.848
R1195 GND.n4433 GND.n4432 22.848
R1196 GND.n4385 GND.n4384 22.848
R1197 GND.n4386 GND.n4385 22.848
R1198 GND.n4351 GND.n4350 22.848
R1199 GND.n4352 GND.n4351 22.848
R1200 GND.n4304 GND.n4303 22.848
R1201 GND.n4305 GND.n4304 22.848
R1202 GND.n4270 GND.n4269 22.848
R1203 GND.n4271 GND.n4270 22.848
R1204 GND.n4223 GND.n4222 22.848
R1205 GND.n4224 GND.n4223 22.848
R1206 GND.n4189 GND.n4188 22.848
R1207 GND.n4190 GND.n4189 22.848
R1208 GND.n4142 GND.n4141 22.848
R1209 GND.n4143 GND.n4142 22.848
R1210 GND.n4108 GND.n4107 22.848
R1211 GND.n4109 GND.n4108 22.848
R1212 GND.n4061 GND.n4060 22.848
R1213 GND.n4062 GND.n4061 22.848
R1214 GND.n4027 GND.n4026 22.848
R1215 GND.n4028 GND.n4027 22.848
R1216 GND.n3980 GND.n3979 22.848
R1217 GND.n3981 GND.n3980 22.848
R1218 GND.n3946 GND.n3945 22.848
R1219 GND.n3947 GND.n3946 22.848
R1220 GND.n3899 GND.n3898 22.848
R1221 GND.n3900 GND.n3899 22.848
R1222 GND.n5178 GND.n5177 22.848
R1223 GND.n5179 GND.n5178 22.848
R1224 GND.n5131 GND.n5130 22.848
R1225 GND.n5132 GND.n5131 22.848
R1226 GND.n5097 GND.n5096 22.848
R1227 GND.n5098 GND.n5097 22.848
R1228 GND.n5050 GND.n5049 22.848
R1229 GND.n5051 GND.n5050 22.848
R1230 GND.n5016 GND.n5015 22.848
R1231 GND.n5017 GND.n5016 22.848
R1232 GND.n4969 GND.n4968 22.848
R1233 GND.n4970 GND.n4969 22.848
R1234 GND.n4935 GND.n4934 22.848
R1235 GND.n4936 GND.n4935 22.848
R1236 GND.n4888 GND.n4887 22.848
R1237 GND.n4889 GND.n4888 22.848
R1238 GND.n4854 GND.n4853 22.848
R1239 GND.n4855 GND.n4854 22.848
R1240 GND.n4807 GND.n4806 22.848
R1241 GND.n4808 GND.n4807 22.848
R1242 GND.n4773 GND.n4772 22.848
R1243 GND.n4774 GND.n4773 22.848
R1244 GND.n4726 GND.n4725 22.848
R1245 GND.n4727 GND.n4726 22.848
R1246 GND.n4692 GND.n4691 22.848
R1247 GND.n4693 GND.n4692 22.848
R1248 GND.n4645 GND.n4644 22.848
R1249 GND.n4646 GND.n4645 22.848
R1250 GND.n4611 GND.n4610 22.848
R1251 GND.n4612 GND.n4611 22.848
R1252 GND.n4564 GND.n4563 22.848
R1253 GND.n4565 GND.n4564 22.848
R1254 GND.n56 GND.n54 10.189
R1255 GND.n16 GND.n14 10.189
R1256 GND.n234 GND.n233 10.189
R1257 GND.n188 GND.n186 10.189
R1258 GND.n153 GND.n152 10.189
R1259 GND.n107 GND.n105 10.189
R1260 GND.n569 GND.n568 10.189
R1261 GND.n523 GND.n521 10.189
R1262 GND.n488 GND.n487 10.189
R1263 GND.n442 GND.n440 10.189
R1264 GND.n407 GND.n406 10.189
R1265 GND.n361 GND.n359 10.189
R1266 GND.n326 GND.n325 10.189
R1267 GND.n280 GND.n278 10.189
R1268 GND.n1230 GND.n1229 10.189
R1269 GND.n1184 GND.n1182 10.189
R1270 GND.n1149 GND.n1148 10.189
R1271 GND.n1103 GND.n1101 10.189
R1272 GND.n1068 GND.n1067 10.189
R1273 GND.n1022 GND.n1020 10.189
R1274 GND.n987 GND.n986 10.189
R1275 GND.n941 GND.n939 10.189
R1276 GND.n906 GND.n905 10.189
R1277 GND.n860 GND.n858 10.189
R1278 GND.n825 GND.n824 10.189
R1279 GND.n779 GND.n777 10.189
R1280 GND.n744 GND.n743 10.189
R1281 GND.n698 GND.n696 10.189
R1282 GND.n663 GND.n662 10.189
R1283 GND.n617 GND.n615 10.189
R1284 GND.n1885 GND.n1884 10.189
R1285 GND.n1839 GND.n1837 10.189
R1286 GND.n1804 GND.n1803 10.189
R1287 GND.n1758 GND.n1756 10.189
R1288 GND.n1723 GND.n1722 10.189
R1289 GND.n1677 GND.n1675 10.189
R1290 GND.n1642 GND.n1641 10.189
R1291 GND.n1596 GND.n1594 10.189
R1292 GND.n1561 GND.n1560 10.189
R1293 GND.n1515 GND.n1513 10.189
R1294 GND.n1480 GND.n1479 10.189
R1295 GND.n1434 GND.n1432 10.189
R1296 GND.n1399 GND.n1398 10.189
R1297 GND.n1353 GND.n1351 10.189
R1298 GND.n1318 GND.n1317 10.189
R1299 GND.n1272 GND.n1270 10.189
R1300 GND.n2550 GND.n2549 10.189
R1301 GND.n2504 GND.n2502 10.189
R1302 GND.n2469 GND.n2468 10.189
R1303 GND.n2423 GND.n2421 10.189
R1304 GND.n2388 GND.n2387 10.189
R1305 GND.n2342 GND.n2340 10.189
R1306 GND.n2307 GND.n2306 10.189
R1307 GND.n2261 GND.n2259 10.189
R1308 GND.n2226 GND.n2225 10.189
R1309 GND.n2180 GND.n2178 10.189
R1310 GND.n2145 GND.n2144 10.189
R1311 GND.n2099 GND.n2097 10.189
R1312 GND.n2064 GND.n2063 10.189
R1313 GND.n2018 GND.n2016 10.189
R1314 GND.n1983 GND.n1982 10.189
R1315 GND.n1937 GND.n1935 10.189
R1316 GND.n3205 GND.n3204 10.189
R1317 GND.n3159 GND.n3157 10.189
R1318 GND.n3124 GND.n3123 10.189
R1319 GND.n3078 GND.n3076 10.189
R1320 GND.n3043 GND.n3042 10.189
R1321 GND.n2997 GND.n2995 10.189
R1322 GND.n2962 GND.n2961 10.189
R1323 GND.n2916 GND.n2914 10.189
R1324 GND.n2881 GND.n2880 10.189
R1325 GND.n2835 GND.n2833 10.189
R1326 GND.n2800 GND.n2799 10.189
R1327 GND.n2754 GND.n2752 10.189
R1328 GND.n2719 GND.n2718 10.189
R1329 GND.n2673 GND.n2671 10.189
R1330 GND.n2638 GND.n2637 10.189
R1331 GND.n2592 GND.n2590 10.189
R1332 GND.n3860 GND.n3859 10.189
R1333 GND.n3814 GND.n3812 10.189
R1334 GND.n3779 GND.n3778 10.189
R1335 GND.n3733 GND.n3731 10.189
R1336 GND.n3698 GND.n3697 10.189
R1337 GND.n3652 GND.n3650 10.189
R1338 GND.n3617 GND.n3616 10.189
R1339 GND.n3571 GND.n3569 10.189
R1340 GND.n3536 GND.n3535 10.189
R1341 GND.n3490 GND.n3488 10.189
R1342 GND.n3455 GND.n3454 10.189
R1343 GND.n3409 GND.n3407 10.189
R1344 GND.n3374 GND.n3373 10.189
R1345 GND.n3328 GND.n3326 10.189
R1346 GND.n3293 GND.n3292 10.189
R1347 GND.n3247 GND.n3245 10.189
R1348 GND.n4515 GND.n4514 10.189
R1349 GND.n4469 GND.n4467 10.189
R1350 GND.n4434 GND.n4433 10.189
R1351 GND.n4388 GND.n4386 10.189
R1352 GND.n4353 GND.n4352 10.189
R1353 GND.n4307 GND.n4305 10.189
R1354 GND.n4272 GND.n4271 10.189
R1355 GND.n4226 GND.n4224 10.189
R1356 GND.n4191 GND.n4190 10.189
R1357 GND.n4145 GND.n4143 10.189
R1358 GND.n4110 GND.n4109 10.189
R1359 GND.n4064 GND.n4062 10.189
R1360 GND.n4029 GND.n4028 10.189
R1361 GND.n3983 GND.n3981 10.189
R1362 GND.n3948 GND.n3947 10.189
R1363 GND.n3902 GND.n3900 10.189
R1364 GND.n5180 GND.n5179 10.189
R1365 GND.n5134 GND.n5132 10.189
R1366 GND.n5099 GND.n5098 10.189
R1367 GND.n5053 GND.n5051 10.189
R1368 GND.n5018 GND.n5017 10.189
R1369 GND.n4972 GND.n4970 10.189
R1370 GND.n4937 GND.n4936 10.189
R1371 GND.n4891 GND.n4889 10.189
R1372 GND.n4856 GND.n4855 10.189
R1373 GND.n4810 GND.n4808 10.189
R1374 GND.n4775 GND.n4774 10.189
R1375 GND.n4729 GND.n4727 10.189
R1376 GND.n4694 GND.n4693 10.189
R1377 GND.n4648 GND.n4646 10.189
R1378 GND.n4613 GND.n4612 10.189
R1379 GND.n4567 GND.n4565 10.189
R1380 GND.n62 GND.n61 9.861
R1381 GND.n22 GND.n21 9.861
R1382 GND.n227 GND.n225 9.861
R1383 GND.n194 GND.n193 9.861
R1384 GND.n146 GND.n144 9.861
R1385 GND.n113 GND.n112 9.861
R1386 GND.n562 GND.n560 9.861
R1387 GND.n529 GND.n528 9.861
R1388 GND.n481 GND.n479 9.861
R1389 GND.n448 GND.n447 9.861
R1390 GND.n400 GND.n398 9.861
R1391 GND.n367 GND.n366 9.861
R1392 GND.n319 GND.n317 9.861
R1393 GND.n286 GND.n285 9.861
R1394 GND.n1223 GND.n1221 9.861
R1395 GND.n1190 GND.n1189 9.861
R1396 GND.n1142 GND.n1140 9.861
R1397 GND.n1109 GND.n1108 9.861
R1398 GND.n1061 GND.n1059 9.861
R1399 GND.n1028 GND.n1027 9.861
R1400 GND.n980 GND.n978 9.861
R1401 GND.n947 GND.n946 9.861
R1402 GND.n899 GND.n897 9.861
R1403 GND.n866 GND.n865 9.861
R1404 GND.n818 GND.n816 9.861
R1405 GND.n785 GND.n784 9.861
R1406 GND.n737 GND.n735 9.861
R1407 GND.n704 GND.n703 9.861
R1408 GND.n656 GND.n654 9.861
R1409 GND.n623 GND.n622 9.861
R1410 GND.n1878 GND.n1876 9.861
R1411 GND.n1845 GND.n1844 9.861
R1412 GND.n1797 GND.n1795 9.861
R1413 GND.n1764 GND.n1763 9.861
R1414 GND.n1716 GND.n1714 9.861
R1415 GND.n1683 GND.n1682 9.861
R1416 GND.n1635 GND.n1633 9.861
R1417 GND.n1602 GND.n1601 9.861
R1418 GND.n1554 GND.n1552 9.861
R1419 GND.n1521 GND.n1520 9.861
R1420 GND.n1473 GND.n1471 9.861
R1421 GND.n1440 GND.n1439 9.861
R1422 GND.n1392 GND.n1390 9.861
R1423 GND.n1359 GND.n1358 9.861
R1424 GND.n1311 GND.n1309 9.861
R1425 GND.n1278 GND.n1277 9.861
R1426 GND.n2543 GND.n2541 9.861
R1427 GND.n2510 GND.n2509 9.861
R1428 GND.n2462 GND.n2460 9.861
R1429 GND.n2429 GND.n2428 9.861
R1430 GND.n2381 GND.n2379 9.861
R1431 GND.n2348 GND.n2347 9.861
R1432 GND.n2300 GND.n2298 9.861
R1433 GND.n2267 GND.n2266 9.861
R1434 GND.n2219 GND.n2217 9.861
R1435 GND.n2186 GND.n2185 9.861
R1436 GND.n2138 GND.n2136 9.861
R1437 GND.n2105 GND.n2104 9.861
R1438 GND.n2057 GND.n2055 9.861
R1439 GND.n2024 GND.n2023 9.861
R1440 GND.n1976 GND.n1974 9.861
R1441 GND.n1943 GND.n1942 9.861
R1442 GND.n3198 GND.n3196 9.861
R1443 GND.n3165 GND.n3164 9.861
R1444 GND.n3117 GND.n3115 9.861
R1445 GND.n3084 GND.n3083 9.861
R1446 GND.n3036 GND.n3034 9.861
R1447 GND.n3003 GND.n3002 9.861
R1448 GND.n2955 GND.n2953 9.861
R1449 GND.n2922 GND.n2921 9.861
R1450 GND.n2874 GND.n2872 9.861
R1451 GND.n2841 GND.n2840 9.861
R1452 GND.n2793 GND.n2791 9.861
R1453 GND.n2760 GND.n2759 9.861
R1454 GND.n2712 GND.n2710 9.861
R1455 GND.n2679 GND.n2678 9.861
R1456 GND.n2631 GND.n2629 9.861
R1457 GND.n2598 GND.n2597 9.861
R1458 GND.n3853 GND.n3851 9.861
R1459 GND.n3820 GND.n3819 9.861
R1460 GND.n3772 GND.n3770 9.861
R1461 GND.n3739 GND.n3738 9.861
R1462 GND.n3691 GND.n3689 9.861
R1463 GND.n3658 GND.n3657 9.861
R1464 GND.n3610 GND.n3608 9.861
R1465 GND.n3577 GND.n3576 9.861
R1466 GND.n3529 GND.n3527 9.861
R1467 GND.n3496 GND.n3495 9.861
R1468 GND.n3448 GND.n3446 9.861
R1469 GND.n3415 GND.n3414 9.861
R1470 GND.n3367 GND.n3365 9.861
R1471 GND.n3334 GND.n3333 9.861
R1472 GND.n3286 GND.n3284 9.861
R1473 GND.n3253 GND.n3252 9.861
R1474 GND.n4508 GND.n4506 9.861
R1475 GND.n4475 GND.n4474 9.861
R1476 GND.n4427 GND.n4425 9.861
R1477 GND.n4394 GND.n4393 9.861
R1478 GND.n4346 GND.n4344 9.861
R1479 GND.n4313 GND.n4312 9.861
R1480 GND.n4265 GND.n4263 9.861
R1481 GND.n4232 GND.n4231 9.861
R1482 GND.n4184 GND.n4182 9.861
R1483 GND.n4151 GND.n4150 9.861
R1484 GND.n4103 GND.n4101 9.861
R1485 GND.n4070 GND.n4069 9.861
R1486 GND.n4022 GND.n4020 9.861
R1487 GND.n3989 GND.n3988 9.861
R1488 GND.n3941 GND.n3939 9.861
R1489 GND.n3908 GND.n3907 9.861
R1490 GND.n5173 GND.n5171 9.861
R1491 GND.n5140 GND.n5139 9.861
R1492 GND.n5092 GND.n5090 9.861
R1493 GND.n5059 GND.n5058 9.861
R1494 GND.n5011 GND.n5009 9.861
R1495 GND.n4978 GND.n4977 9.861
R1496 GND.n4930 GND.n4928 9.861
R1497 GND.n4897 GND.n4896 9.861
R1498 GND.n4849 GND.n4847 9.861
R1499 GND.n4816 GND.n4815 9.861
R1500 GND.n4768 GND.n4766 9.861
R1501 GND.n4735 GND.n4734 9.861
R1502 GND.n4687 GND.n4685 9.861
R1503 GND.n4654 GND.n4653 9.861
R1504 GND.n4606 GND.n4604 9.861
R1505 GND.n4573 GND.n4572 9.861
R1506 GND.n63 GND.n62 9.457
R1507 GND.n23 GND.n22 9.457
R1508 GND.n228 GND.n227 9.457
R1509 GND.n195 GND.n194 9.457
R1510 GND.n147 GND.n146 9.457
R1511 GND.n114 GND.n113 9.457
R1512 GND.n563 GND.n562 9.457
R1513 GND.n530 GND.n529 9.457
R1514 GND.n482 GND.n481 9.457
R1515 GND.n449 GND.n448 9.457
R1516 GND.n401 GND.n400 9.457
R1517 GND.n368 GND.n367 9.457
R1518 GND.n320 GND.n319 9.457
R1519 GND.n287 GND.n286 9.457
R1520 GND.n1224 GND.n1223 9.457
R1521 GND.n1191 GND.n1190 9.457
R1522 GND.n1143 GND.n1142 9.457
R1523 GND.n1110 GND.n1109 9.457
R1524 GND.n1062 GND.n1061 9.457
R1525 GND.n1029 GND.n1028 9.457
R1526 GND.n981 GND.n980 9.457
R1527 GND.n948 GND.n947 9.457
R1528 GND.n900 GND.n899 9.457
R1529 GND.n867 GND.n866 9.457
R1530 GND.n819 GND.n818 9.457
R1531 GND.n786 GND.n785 9.457
R1532 GND.n738 GND.n737 9.457
R1533 GND.n705 GND.n704 9.457
R1534 GND.n657 GND.n656 9.457
R1535 GND.n624 GND.n623 9.457
R1536 GND.n1879 GND.n1878 9.457
R1537 GND.n1846 GND.n1845 9.457
R1538 GND.n1798 GND.n1797 9.457
R1539 GND.n1765 GND.n1764 9.457
R1540 GND.n1717 GND.n1716 9.457
R1541 GND.n1684 GND.n1683 9.457
R1542 GND.n1636 GND.n1635 9.457
R1543 GND.n1603 GND.n1602 9.457
R1544 GND.n1555 GND.n1554 9.457
R1545 GND.n1522 GND.n1521 9.457
R1546 GND.n1474 GND.n1473 9.457
R1547 GND.n1441 GND.n1440 9.457
R1548 GND.n1393 GND.n1392 9.457
R1549 GND.n1360 GND.n1359 9.457
R1550 GND.n1312 GND.n1311 9.457
R1551 GND.n1279 GND.n1278 9.457
R1552 GND.n2544 GND.n2543 9.457
R1553 GND.n2511 GND.n2510 9.457
R1554 GND.n2463 GND.n2462 9.457
R1555 GND.n2430 GND.n2429 9.457
R1556 GND.n2382 GND.n2381 9.457
R1557 GND.n2349 GND.n2348 9.457
R1558 GND.n2301 GND.n2300 9.457
R1559 GND.n2268 GND.n2267 9.457
R1560 GND.n2220 GND.n2219 9.457
R1561 GND.n2187 GND.n2186 9.457
R1562 GND.n2139 GND.n2138 9.457
R1563 GND.n2106 GND.n2105 9.457
R1564 GND.n2058 GND.n2057 9.457
R1565 GND.n2025 GND.n2024 9.457
R1566 GND.n1977 GND.n1976 9.457
R1567 GND.n1944 GND.n1943 9.457
R1568 GND.n3199 GND.n3198 9.457
R1569 GND.n3166 GND.n3165 9.457
R1570 GND.n3118 GND.n3117 9.457
R1571 GND.n3085 GND.n3084 9.457
R1572 GND.n3037 GND.n3036 9.457
R1573 GND.n3004 GND.n3003 9.457
R1574 GND.n2956 GND.n2955 9.457
R1575 GND.n2923 GND.n2922 9.457
R1576 GND.n2875 GND.n2874 9.457
R1577 GND.n2842 GND.n2841 9.457
R1578 GND.n2794 GND.n2793 9.457
R1579 GND.n2761 GND.n2760 9.457
R1580 GND.n2713 GND.n2712 9.457
R1581 GND.n2680 GND.n2679 9.457
R1582 GND.n2632 GND.n2631 9.457
R1583 GND.n2599 GND.n2598 9.457
R1584 GND.n3854 GND.n3853 9.457
R1585 GND.n3821 GND.n3820 9.457
R1586 GND.n3773 GND.n3772 9.457
R1587 GND.n3740 GND.n3739 9.457
R1588 GND.n3692 GND.n3691 9.457
R1589 GND.n3659 GND.n3658 9.457
R1590 GND.n3611 GND.n3610 9.457
R1591 GND.n3578 GND.n3577 9.457
R1592 GND.n3530 GND.n3529 9.457
R1593 GND.n3497 GND.n3496 9.457
R1594 GND.n3449 GND.n3448 9.457
R1595 GND.n3416 GND.n3415 9.457
R1596 GND.n3368 GND.n3367 9.457
R1597 GND.n3335 GND.n3334 9.457
R1598 GND.n3287 GND.n3286 9.457
R1599 GND.n3254 GND.n3253 9.457
R1600 GND.n4509 GND.n4508 9.457
R1601 GND.n4476 GND.n4475 9.457
R1602 GND.n4428 GND.n4427 9.457
R1603 GND.n4395 GND.n4394 9.457
R1604 GND.n4347 GND.n4346 9.457
R1605 GND.n4314 GND.n4313 9.457
R1606 GND.n4266 GND.n4265 9.457
R1607 GND.n4233 GND.n4232 9.457
R1608 GND.n4185 GND.n4184 9.457
R1609 GND.n4152 GND.n4151 9.457
R1610 GND.n4104 GND.n4103 9.457
R1611 GND.n4071 GND.n4070 9.457
R1612 GND.n4023 GND.n4022 9.457
R1613 GND.n3990 GND.n3989 9.457
R1614 GND.n3942 GND.n3941 9.457
R1615 GND.n3909 GND.n3908 9.457
R1616 GND.n5174 GND.n5173 9.457
R1617 GND.n5141 GND.n5140 9.457
R1618 GND.n5093 GND.n5092 9.457
R1619 GND.n5060 GND.n5059 9.457
R1620 GND.n5012 GND.n5011 9.457
R1621 GND.n4979 GND.n4978 9.457
R1622 GND.n4931 GND.n4930 9.457
R1623 GND.n4898 GND.n4897 9.457
R1624 GND.n4850 GND.n4849 9.457
R1625 GND.n4817 GND.n4816 9.457
R1626 GND.n4769 GND.n4768 9.457
R1627 GND.n4736 GND.n4735 9.457
R1628 GND.n4688 GND.n4687 9.457
R1629 GND.n4655 GND.n4654 9.457
R1630 GND.n4607 GND.n4606 9.457
R1631 GND.n4574 GND.n4573 9.457
R1632 GND.n86 GND.n85 9.3
R1633 GND.n88 GND.n87 9.3
R1634 GND.n67 GND.n66 9.3
R1635 GND.n65 GND.n64 9.3
R1636 GND.n75 GND.n74 9.3
R1637 GND.n74 GND.n73 9.3
R1638 GND.n84 GND.n83 9.3
R1639 GND.n83 GND.n82 9.3
R1640 GND.n57 GND.n56 9.3
R1641 GND.n56 GND.n55 9.3
R1642 GND.n46 GND.n45 9.3
R1643 GND.n27 GND.n26 9.3
R1644 GND.n25 GND.n24 9.3
R1645 GND.n35 GND.n34 9.3
R1646 GND.n34 GND.n33 9.3
R1647 GND.n44 GND.n43 9.3
R1648 GND.n43 GND.n42 9.3
R1649 GND.n48 GND.n47 9.3
R1650 GND.n17 GND.n16 9.3
R1651 GND.n16 GND.n15 9.3
R1652 GND.n258 GND.n257 9.3
R1653 GND.n239 GND.n238 9.3
R1654 GND.n237 GND.n236 9.3
R1655 GND.n260 GND.n259 9.3
R1656 GND.n247 GND.n246 9.3
R1657 GND.n246 GND.n245 9.3
R1658 GND.n256 GND.n255 9.3
R1659 GND.n255 GND.n254 9.3
R1660 GND.n235 GND.n234 9.3
R1661 GND.n218 GND.n217 9.3
R1662 GND.n199 GND.n198 9.3
R1663 GND.n197 GND.n196 9.3
R1664 GND.n207 GND.n206 9.3
R1665 GND.n206 GND.n205 9.3
R1666 GND.n216 GND.n215 9.3
R1667 GND.n215 GND.n214 9.3
R1668 GND.n220 GND.n219 9.3
R1669 GND.n189 GND.n188 9.3
R1670 GND.n188 GND.n187 9.3
R1671 GND.n177 GND.n176 9.3
R1672 GND.n158 GND.n157 9.3
R1673 GND.n156 GND.n155 9.3
R1674 GND.n179 GND.n178 9.3
R1675 GND.n166 GND.n165 9.3
R1676 GND.n165 GND.n164 9.3
R1677 GND.n175 GND.n174 9.3
R1678 GND.n174 GND.n173 9.3
R1679 GND.n154 GND.n153 9.3
R1680 GND.n137 GND.n136 9.3
R1681 GND.n118 GND.n117 9.3
R1682 GND.n116 GND.n115 9.3
R1683 GND.n126 GND.n125 9.3
R1684 GND.n125 GND.n124 9.3
R1685 GND.n135 GND.n134 9.3
R1686 GND.n134 GND.n133 9.3
R1687 GND.n139 GND.n138 9.3
R1688 GND.n108 GND.n107 9.3
R1689 GND.n107 GND.n106 9.3
R1690 GND.n593 GND.n592 9.3
R1691 GND.n574 GND.n573 9.3
R1692 GND.n572 GND.n571 9.3
R1693 GND.n595 GND.n594 9.3
R1694 GND.n582 GND.n581 9.3
R1695 GND.n581 GND.n580 9.3
R1696 GND.n591 GND.n590 9.3
R1697 GND.n590 GND.n589 9.3
R1698 GND.n570 GND.n569 9.3
R1699 GND.n553 GND.n552 9.3
R1700 GND.n534 GND.n533 9.3
R1701 GND.n532 GND.n531 9.3
R1702 GND.n542 GND.n541 9.3
R1703 GND.n541 GND.n540 9.3
R1704 GND.n551 GND.n550 9.3
R1705 GND.n550 GND.n549 9.3
R1706 GND.n555 GND.n554 9.3
R1707 GND.n524 GND.n523 9.3
R1708 GND.n523 GND.n522 9.3
R1709 GND.n512 GND.n511 9.3
R1710 GND.n493 GND.n492 9.3
R1711 GND.n491 GND.n490 9.3
R1712 GND.n514 GND.n513 9.3
R1713 GND.n501 GND.n500 9.3
R1714 GND.n500 GND.n499 9.3
R1715 GND.n510 GND.n509 9.3
R1716 GND.n509 GND.n508 9.3
R1717 GND.n489 GND.n488 9.3
R1718 GND.n472 GND.n471 9.3
R1719 GND.n453 GND.n452 9.3
R1720 GND.n451 GND.n450 9.3
R1721 GND.n461 GND.n460 9.3
R1722 GND.n460 GND.n459 9.3
R1723 GND.n470 GND.n469 9.3
R1724 GND.n469 GND.n468 9.3
R1725 GND.n474 GND.n473 9.3
R1726 GND.n443 GND.n442 9.3
R1727 GND.n442 GND.n441 9.3
R1728 GND.n431 GND.n430 9.3
R1729 GND.n412 GND.n411 9.3
R1730 GND.n410 GND.n409 9.3
R1731 GND.n433 GND.n432 9.3
R1732 GND.n420 GND.n419 9.3
R1733 GND.n419 GND.n418 9.3
R1734 GND.n429 GND.n428 9.3
R1735 GND.n428 GND.n427 9.3
R1736 GND.n408 GND.n407 9.3
R1737 GND.n391 GND.n390 9.3
R1738 GND.n372 GND.n371 9.3
R1739 GND.n370 GND.n369 9.3
R1740 GND.n380 GND.n379 9.3
R1741 GND.n379 GND.n378 9.3
R1742 GND.n389 GND.n388 9.3
R1743 GND.n388 GND.n387 9.3
R1744 GND.n393 GND.n392 9.3
R1745 GND.n362 GND.n361 9.3
R1746 GND.n361 GND.n360 9.3
R1747 GND.n350 GND.n349 9.3
R1748 GND.n331 GND.n330 9.3
R1749 GND.n329 GND.n328 9.3
R1750 GND.n352 GND.n351 9.3
R1751 GND.n339 GND.n338 9.3
R1752 GND.n338 GND.n337 9.3
R1753 GND.n348 GND.n347 9.3
R1754 GND.n347 GND.n346 9.3
R1755 GND.n327 GND.n326 9.3
R1756 GND.n310 GND.n309 9.3
R1757 GND.n291 GND.n290 9.3
R1758 GND.n289 GND.n288 9.3
R1759 GND.n299 GND.n298 9.3
R1760 GND.n298 GND.n297 9.3
R1761 GND.n308 GND.n307 9.3
R1762 GND.n307 GND.n306 9.3
R1763 GND.n312 GND.n311 9.3
R1764 GND.n281 GND.n280 9.3
R1765 GND.n280 GND.n279 9.3
R1766 GND.n1254 GND.n1253 9.3
R1767 GND.n1235 GND.n1234 9.3
R1768 GND.n1233 GND.n1232 9.3
R1769 GND.n1256 GND.n1255 9.3
R1770 GND.n1243 GND.n1242 9.3
R1771 GND.n1242 GND.n1241 9.3
R1772 GND.n1252 GND.n1251 9.3
R1773 GND.n1251 GND.n1250 9.3
R1774 GND.n1231 GND.n1230 9.3
R1775 GND.n1214 GND.n1213 9.3
R1776 GND.n1195 GND.n1194 9.3
R1777 GND.n1193 GND.n1192 9.3
R1778 GND.n1203 GND.n1202 9.3
R1779 GND.n1202 GND.n1201 9.3
R1780 GND.n1212 GND.n1211 9.3
R1781 GND.n1211 GND.n1210 9.3
R1782 GND.n1216 GND.n1215 9.3
R1783 GND.n1185 GND.n1184 9.3
R1784 GND.n1184 GND.n1183 9.3
R1785 GND.n1173 GND.n1172 9.3
R1786 GND.n1154 GND.n1153 9.3
R1787 GND.n1152 GND.n1151 9.3
R1788 GND.n1175 GND.n1174 9.3
R1789 GND.n1162 GND.n1161 9.3
R1790 GND.n1161 GND.n1160 9.3
R1791 GND.n1171 GND.n1170 9.3
R1792 GND.n1170 GND.n1169 9.3
R1793 GND.n1150 GND.n1149 9.3
R1794 GND.n1133 GND.n1132 9.3
R1795 GND.n1114 GND.n1113 9.3
R1796 GND.n1112 GND.n1111 9.3
R1797 GND.n1122 GND.n1121 9.3
R1798 GND.n1121 GND.n1120 9.3
R1799 GND.n1131 GND.n1130 9.3
R1800 GND.n1130 GND.n1129 9.3
R1801 GND.n1135 GND.n1134 9.3
R1802 GND.n1104 GND.n1103 9.3
R1803 GND.n1103 GND.n1102 9.3
R1804 GND.n1092 GND.n1091 9.3
R1805 GND.n1073 GND.n1072 9.3
R1806 GND.n1071 GND.n1070 9.3
R1807 GND.n1094 GND.n1093 9.3
R1808 GND.n1081 GND.n1080 9.3
R1809 GND.n1080 GND.n1079 9.3
R1810 GND.n1090 GND.n1089 9.3
R1811 GND.n1089 GND.n1088 9.3
R1812 GND.n1069 GND.n1068 9.3
R1813 GND.n1052 GND.n1051 9.3
R1814 GND.n1033 GND.n1032 9.3
R1815 GND.n1031 GND.n1030 9.3
R1816 GND.n1041 GND.n1040 9.3
R1817 GND.n1040 GND.n1039 9.3
R1818 GND.n1050 GND.n1049 9.3
R1819 GND.n1049 GND.n1048 9.3
R1820 GND.n1054 GND.n1053 9.3
R1821 GND.n1023 GND.n1022 9.3
R1822 GND.n1022 GND.n1021 9.3
R1823 GND.n1011 GND.n1010 9.3
R1824 GND.n992 GND.n991 9.3
R1825 GND.n990 GND.n989 9.3
R1826 GND.n1013 GND.n1012 9.3
R1827 GND.n1000 GND.n999 9.3
R1828 GND.n999 GND.n998 9.3
R1829 GND.n1009 GND.n1008 9.3
R1830 GND.n1008 GND.n1007 9.3
R1831 GND.n988 GND.n987 9.3
R1832 GND.n971 GND.n970 9.3
R1833 GND.n952 GND.n951 9.3
R1834 GND.n950 GND.n949 9.3
R1835 GND.n960 GND.n959 9.3
R1836 GND.n959 GND.n958 9.3
R1837 GND.n969 GND.n968 9.3
R1838 GND.n968 GND.n967 9.3
R1839 GND.n973 GND.n972 9.3
R1840 GND.n942 GND.n941 9.3
R1841 GND.n941 GND.n940 9.3
R1842 GND.n930 GND.n929 9.3
R1843 GND.n911 GND.n910 9.3
R1844 GND.n909 GND.n908 9.3
R1845 GND.n932 GND.n931 9.3
R1846 GND.n919 GND.n918 9.3
R1847 GND.n918 GND.n917 9.3
R1848 GND.n928 GND.n927 9.3
R1849 GND.n927 GND.n926 9.3
R1850 GND.n907 GND.n906 9.3
R1851 GND.n890 GND.n889 9.3
R1852 GND.n871 GND.n870 9.3
R1853 GND.n869 GND.n868 9.3
R1854 GND.n879 GND.n878 9.3
R1855 GND.n878 GND.n877 9.3
R1856 GND.n888 GND.n887 9.3
R1857 GND.n887 GND.n886 9.3
R1858 GND.n892 GND.n891 9.3
R1859 GND.n861 GND.n860 9.3
R1860 GND.n860 GND.n859 9.3
R1861 GND.n849 GND.n848 9.3
R1862 GND.n830 GND.n829 9.3
R1863 GND.n828 GND.n827 9.3
R1864 GND.n851 GND.n850 9.3
R1865 GND.n838 GND.n837 9.3
R1866 GND.n837 GND.n836 9.3
R1867 GND.n847 GND.n846 9.3
R1868 GND.n846 GND.n845 9.3
R1869 GND.n826 GND.n825 9.3
R1870 GND.n809 GND.n808 9.3
R1871 GND.n790 GND.n789 9.3
R1872 GND.n788 GND.n787 9.3
R1873 GND.n798 GND.n797 9.3
R1874 GND.n797 GND.n796 9.3
R1875 GND.n807 GND.n806 9.3
R1876 GND.n806 GND.n805 9.3
R1877 GND.n811 GND.n810 9.3
R1878 GND.n780 GND.n779 9.3
R1879 GND.n779 GND.n778 9.3
R1880 GND.n768 GND.n767 9.3
R1881 GND.n749 GND.n748 9.3
R1882 GND.n747 GND.n746 9.3
R1883 GND.n770 GND.n769 9.3
R1884 GND.n757 GND.n756 9.3
R1885 GND.n756 GND.n755 9.3
R1886 GND.n766 GND.n765 9.3
R1887 GND.n765 GND.n764 9.3
R1888 GND.n745 GND.n744 9.3
R1889 GND.n728 GND.n727 9.3
R1890 GND.n709 GND.n708 9.3
R1891 GND.n707 GND.n706 9.3
R1892 GND.n717 GND.n716 9.3
R1893 GND.n716 GND.n715 9.3
R1894 GND.n726 GND.n725 9.3
R1895 GND.n725 GND.n724 9.3
R1896 GND.n730 GND.n729 9.3
R1897 GND.n699 GND.n698 9.3
R1898 GND.n698 GND.n697 9.3
R1899 GND.n687 GND.n686 9.3
R1900 GND.n668 GND.n667 9.3
R1901 GND.n666 GND.n665 9.3
R1902 GND.n689 GND.n688 9.3
R1903 GND.n676 GND.n675 9.3
R1904 GND.n675 GND.n674 9.3
R1905 GND.n685 GND.n684 9.3
R1906 GND.n684 GND.n683 9.3
R1907 GND.n664 GND.n663 9.3
R1908 GND.n647 GND.n646 9.3
R1909 GND.n628 GND.n627 9.3
R1910 GND.n626 GND.n625 9.3
R1911 GND.n636 GND.n635 9.3
R1912 GND.n635 GND.n634 9.3
R1913 GND.n645 GND.n644 9.3
R1914 GND.n644 GND.n643 9.3
R1915 GND.n649 GND.n648 9.3
R1916 GND.n618 GND.n617 9.3
R1917 GND.n617 GND.n616 9.3
R1918 GND.n1909 GND.n1908 9.3
R1919 GND.n1890 GND.n1889 9.3
R1920 GND.n1888 GND.n1887 9.3
R1921 GND.n1911 GND.n1910 9.3
R1922 GND.n1898 GND.n1897 9.3
R1923 GND.n1897 GND.n1896 9.3
R1924 GND.n1907 GND.n1906 9.3
R1925 GND.n1906 GND.n1905 9.3
R1926 GND.n1886 GND.n1885 9.3
R1927 GND.n1869 GND.n1868 9.3
R1928 GND.n1850 GND.n1849 9.3
R1929 GND.n1848 GND.n1847 9.3
R1930 GND.n1858 GND.n1857 9.3
R1931 GND.n1857 GND.n1856 9.3
R1932 GND.n1867 GND.n1866 9.3
R1933 GND.n1866 GND.n1865 9.3
R1934 GND.n1871 GND.n1870 9.3
R1935 GND.n1840 GND.n1839 9.3
R1936 GND.n1839 GND.n1838 9.3
R1937 GND.n1828 GND.n1827 9.3
R1938 GND.n1809 GND.n1808 9.3
R1939 GND.n1807 GND.n1806 9.3
R1940 GND.n1830 GND.n1829 9.3
R1941 GND.n1817 GND.n1816 9.3
R1942 GND.n1816 GND.n1815 9.3
R1943 GND.n1826 GND.n1825 9.3
R1944 GND.n1825 GND.n1824 9.3
R1945 GND.n1805 GND.n1804 9.3
R1946 GND.n1788 GND.n1787 9.3
R1947 GND.n1769 GND.n1768 9.3
R1948 GND.n1767 GND.n1766 9.3
R1949 GND.n1777 GND.n1776 9.3
R1950 GND.n1776 GND.n1775 9.3
R1951 GND.n1786 GND.n1785 9.3
R1952 GND.n1785 GND.n1784 9.3
R1953 GND.n1790 GND.n1789 9.3
R1954 GND.n1759 GND.n1758 9.3
R1955 GND.n1758 GND.n1757 9.3
R1956 GND.n1747 GND.n1746 9.3
R1957 GND.n1728 GND.n1727 9.3
R1958 GND.n1726 GND.n1725 9.3
R1959 GND.n1749 GND.n1748 9.3
R1960 GND.n1736 GND.n1735 9.3
R1961 GND.n1735 GND.n1734 9.3
R1962 GND.n1745 GND.n1744 9.3
R1963 GND.n1744 GND.n1743 9.3
R1964 GND.n1724 GND.n1723 9.3
R1965 GND.n1707 GND.n1706 9.3
R1966 GND.n1688 GND.n1687 9.3
R1967 GND.n1686 GND.n1685 9.3
R1968 GND.n1696 GND.n1695 9.3
R1969 GND.n1695 GND.n1694 9.3
R1970 GND.n1705 GND.n1704 9.3
R1971 GND.n1704 GND.n1703 9.3
R1972 GND.n1709 GND.n1708 9.3
R1973 GND.n1678 GND.n1677 9.3
R1974 GND.n1677 GND.n1676 9.3
R1975 GND.n1666 GND.n1665 9.3
R1976 GND.n1647 GND.n1646 9.3
R1977 GND.n1645 GND.n1644 9.3
R1978 GND.n1668 GND.n1667 9.3
R1979 GND.n1655 GND.n1654 9.3
R1980 GND.n1654 GND.n1653 9.3
R1981 GND.n1664 GND.n1663 9.3
R1982 GND.n1663 GND.n1662 9.3
R1983 GND.n1643 GND.n1642 9.3
R1984 GND.n1626 GND.n1625 9.3
R1985 GND.n1607 GND.n1606 9.3
R1986 GND.n1605 GND.n1604 9.3
R1987 GND.n1615 GND.n1614 9.3
R1988 GND.n1614 GND.n1613 9.3
R1989 GND.n1624 GND.n1623 9.3
R1990 GND.n1623 GND.n1622 9.3
R1991 GND.n1628 GND.n1627 9.3
R1992 GND.n1597 GND.n1596 9.3
R1993 GND.n1596 GND.n1595 9.3
R1994 GND.n1585 GND.n1584 9.3
R1995 GND.n1566 GND.n1565 9.3
R1996 GND.n1564 GND.n1563 9.3
R1997 GND.n1587 GND.n1586 9.3
R1998 GND.n1574 GND.n1573 9.3
R1999 GND.n1573 GND.n1572 9.3
R2000 GND.n1583 GND.n1582 9.3
R2001 GND.n1582 GND.n1581 9.3
R2002 GND.n1562 GND.n1561 9.3
R2003 GND.n1545 GND.n1544 9.3
R2004 GND.n1526 GND.n1525 9.3
R2005 GND.n1524 GND.n1523 9.3
R2006 GND.n1534 GND.n1533 9.3
R2007 GND.n1533 GND.n1532 9.3
R2008 GND.n1543 GND.n1542 9.3
R2009 GND.n1542 GND.n1541 9.3
R2010 GND.n1547 GND.n1546 9.3
R2011 GND.n1516 GND.n1515 9.3
R2012 GND.n1515 GND.n1514 9.3
R2013 GND.n1504 GND.n1503 9.3
R2014 GND.n1485 GND.n1484 9.3
R2015 GND.n1483 GND.n1482 9.3
R2016 GND.n1506 GND.n1505 9.3
R2017 GND.n1493 GND.n1492 9.3
R2018 GND.n1492 GND.n1491 9.3
R2019 GND.n1502 GND.n1501 9.3
R2020 GND.n1501 GND.n1500 9.3
R2021 GND.n1481 GND.n1480 9.3
R2022 GND.n1464 GND.n1463 9.3
R2023 GND.n1445 GND.n1444 9.3
R2024 GND.n1443 GND.n1442 9.3
R2025 GND.n1453 GND.n1452 9.3
R2026 GND.n1452 GND.n1451 9.3
R2027 GND.n1462 GND.n1461 9.3
R2028 GND.n1461 GND.n1460 9.3
R2029 GND.n1466 GND.n1465 9.3
R2030 GND.n1435 GND.n1434 9.3
R2031 GND.n1434 GND.n1433 9.3
R2032 GND.n1423 GND.n1422 9.3
R2033 GND.n1404 GND.n1403 9.3
R2034 GND.n1402 GND.n1401 9.3
R2035 GND.n1425 GND.n1424 9.3
R2036 GND.n1412 GND.n1411 9.3
R2037 GND.n1411 GND.n1410 9.3
R2038 GND.n1421 GND.n1420 9.3
R2039 GND.n1420 GND.n1419 9.3
R2040 GND.n1400 GND.n1399 9.3
R2041 GND.n1383 GND.n1382 9.3
R2042 GND.n1364 GND.n1363 9.3
R2043 GND.n1362 GND.n1361 9.3
R2044 GND.n1372 GND.n1371 9.3
R2045 GND.n1371 GND.n1370 9.3
R2046 GND.n1381 GND.n1380 9.3
R2047 GND.n1380 GND.n1379 9.3
R2048 GND.n1385 GND.n1384 9.3
R2049 GND.n1354 GND.n1353 9.3
R2050 GND.n1353 GND.n1352 9.3
R2051 GND.n1342 GND.n1341 9.3
R2052 GND.n1323 GND.n1322 9.3
R2053 GND.n1321 GND.n1320 9.3
R2054 GND.n1344 GND.n1343 9.3
R2055 GND.n1331 GND.n1330 9.3
R2056 GND.n1330 GND.n1329 9.3
R2057 GND.n1340 GND.n1339 9.3
R2058 GND.n1339 GND.n1338 9.3
R2059 GND.n1319 GND.n1318 9.3
R2060 GND.n1302 GND.n1301 9.3
R2061 GND.n1283 GND.n1282 9.3
R2062 GND.n1281 GND.n1280 9.3
R2063 GND.n1291 GND.n1290 9.3
R2064 GND.n1290 GND.n1289 9.3
R2065 GND.n1300 GND.n1299 9.3
R2066 GND.n1299 GND.n1298 9.3
R2067 GND.n1304 GND.n1303 9.3
R2068 GND.n1273 GND.n1272 9.3
R2069 GND.n1272 GND.n1271 9.3
R2070 GND.n2574 GND.n2573 9.3
R2071 GND.n2555 GND.n2554 9.3
R2072 GND.n2553 GND.n2552 9.3
R2073 GND.n2576 GND.n2575 9.3
R2074 GND.n2563 GND.n2562 9.3
R2075 GND.n2562 GND.n2561 9.3
R2076 GND.n2572 GND.n2571 9.3
R2077 GND.n2571 GND.n2570 9.3
R2078 GND.n2551 GND.n2550 9.3
R2079 GND.n2534 GND.n2533 9.3
R2080 GND.n2515 GND.n2514 9.3
R2081 GND.n2513 GND.n2512 9.3
R2082 GND.n2523 GND.n2522 9.3
R2083 GND.n2522 GND.n2521 9.3
R2084 GND.n2532 GND.n2531 9.3
R2085 GND.n2531 GND.n2530 9.3
R2086 GND.n2536 GND.n2535 9.3
R2087 GND.n2505 GND.n2504 9.3
R2088 GND.n2504 GND.n2503 9.3
R2089 GND.n2493 GND.n2492 9.3
R2090 GND.n2474 GND.n2473 9.3
R2091 GND.n2472 GND.n2471 9.3
R2092 GND.n2495 GND.n2494 9.3
R2093 GND.n2482 GND.n2481 9.3
R2094 GND.n2481 GND.n2480 9.3
R2095 GND.n2491 GND.n2490 9.3
R2096 GND.n2490 GND.n2489 9.3
R2097 GND.n2470 GND.n2469 9.3
R2098 GND.n2453 GND.n2452 9.3
R2099 GND.n2434 GND.n2433 9.3
R2100 GND.n2432 GND.n2431 9.3
R2101 GND.n2442 GND.n2441 9.3
R2102 GND.n2441 GND.n2440 9.3
R2103 GND.n2451 GND.n2450 9.3
R2104 GND.n2450 GND.n2449 9.3
R2105 GND.n2455 GND.n2454 9.3
R2106 GND.n2424 GND.n2423 9.3
R2107 GND.n2423 GND.n2422 9.3
R2108 GND.n2412 GND.n2411 9.3
R2109 GND.n2393 GND.n2392 9.3
R2110 GND.n2391 GND.n2390 9.3
R2111 GND.n2414 GND.n2413 9.3
R2112 GND.n2401 GND.n2400 9.3
R2113 GND.n2400 GND.n2399 9.3
R2114 GND.n2410 GND.n2409 9.3
R2115 GND.n2409 GND.n2408 9.3
R2116 GND.n2389 GND.n2388 9.3
R2117 GND.n2372 GND.n2371 9.3
R2118 GND.n2353 GND.n2352 9.3
R2119 GND.n2351 GND.n2350 9.3
R2120 GND.n2361 GND.n2360 9.3
R2121 GND.n2360 GND.n2359 9.3
R2122 GND.n2370 GND.n2369 9.3
R2123 GND.n2369 GND.n2368 9.3
R2124 GND.n2374 GND.n2373 9.3
R2125 GND.n2343 GND.n2342 9.3
R2126 GND.n2342 GND.n2341 9.3
R2127 GND.n2331 GND.n2330 9.3
R2128 GND.n2312 GND.n2311 9.3
R2129 GND.n2310 GND.n2309 9.3
R2130 GND.n2333 GND.n2332 9.3
R2131 GND.n2320 GND.n2319 9.3
R2132 GND.n2319 GND.n2318 9.3
R2133 GND.n2329 GND.n2328 9.3
R2134 GND.n2328 GND.n2327 9.3
R2135 GND.n2308 GND.n2307 9.3
R2136 GND.n2291 GND.n2290 9.3
R2137 GND.n2272 GND.n2271 9.3
R2138 GND.n2270 GND.n2269 9.3
R2139 GND.n2280 GND.n2279 9.3
R2140 GND.n2279 GND.n2278 9.3
R2141 GND.n2289 GND.n2288 9.3
R2142 GND.n2288 GND.n2287 9.3
R2143 GND.n2293 GND.n2292 9.3
R2144 GND.n2262 GND.n2261 9.3
R2145 GND.n2261 GND.n2260 9.3
R2146 GND.n2250 GND.n2249 9.3
R2147 GND.n2231 GND.n2230 9.3
R2148 GND.n2229 GND.n2228 9.3
R2149 GND.n2252 GND.n2251 9.3
R2150 GND.n2239 GND.n2238 9.3
R2151 GND.n2238 GND.n2237 9.3
R2152 GND.n2248 GND.n2247 9.3
R2153 GND.n2247 GND.n2246 9.3
R2154 GND.n2227 GND.n2226 9.3
R2155 GND.n2210 GND.n2209 9.3
R2156 GND.n2191 GND.n2190 9.3
R2157 GND.n2189 GND.n2188 9.3
R2158 GND.n2199 GND.n2198 9.3
R2159 GND.n2198 GND.n2197 9.3
R2160 GND.n2208 GND.n2207 9.3
R2161 GND.n2207 GND.n2206 9.3
R2162 GND.n2212 GND.n2211 9.3
R2163 GND.n2181 GND.n2180 9.3
R2164 GND.n2180 GND.n2179 9.3
R2165 GND.n2169 GND.n2168 9.3
R2166 GND.n2150 GND.n2149 9.3
R2167 GND.n2148 GND.n2147 9.3
R2168 GND.n2171 GND.n2170 9.3
R2169 GND.n2158 GND.n2157 9.3
R2170 GND.n2157 GND.n2156 9.3
R2171 GND.n2167 GND.n2166 9.3
R2172 GND.n2166 GND.n2165 9.3
R2173 GND.n2146 GND.n2145 9.3
R2174 GND.n2129 GND.n2128 9.3
R2175 GND.n2110 GND.n2109 9.3
R2176 GND.n2108 GND.n2107 9.3
R2177 GND.n2118 GND.n2117 9.3
R2178 GND.n2117 GND.n2116 9.3
R2179 GND.n2127 GND.n2126 9.3
R2180 GND.n2126 GND.n2125 9.3
R2181 GND.n2131 GND.n2130 9.3
R2182 GND.n2100 GND.n2099 9.3
R2183 GND.n2099 GND.n2098 9.3
R2184 GND.n2088 GND.n2087 9.3
R2185 GND.n2069 GND.n2068 9.3
R2186 GND.n2067 GND.n2066 9.3
R2187 GND.n2090 GND.n2089 9.3
R2188 GND.n2077 GND.n2076 9.3
R2189 GND.n2076 GND.n2075 9.3
R2190 GND.n2086 GND.n2085 9.3
R2191 GND.n2085 GND.n2084 9.3
R2192 GND.n2065 GND.n2064 9.3
R2193 GND.n2048 GND.n2047 9.3
R2194 GND.n2029 GND.n2028 9.3
R2195 GND.n2027 GND.n2026 9.3
R2196 GND.n2037 GND.n2036 9.3
R2197 GND.n2036 GND.n2035 9.3
R2198 GND.n2046 GND.n2045 9.3
R2199 GND.n2045 GND.n2044 9.3
R2200 GND.n2050 GND.n2049 9.3
R2201 GND.n2019 GND.n2018 9.3
R2202 GND.n2018 GND.n2017 9.3
R2203 GND.n2007 GND.n2006 9.3
R2204 GND.n1988 GND.n1987 9.3
R2205 GND.n1986 GND.n1985 9.3
R2206 GND.n2009 GND.n2008 9.3
R2207 GND.n1996 GND.n1995 9.3
R2208 GND.n1995 GND.n1994 9.3
R2209 GND.n2005 GND.n2004 9.3
R2210 GND.n2004 GND.n2003 9.3
R2211 GND.n1984 GND.n1983 9.3
R2212 GND.n1967 GND.n1966 9.3
R2213 GND.n1948 GND.n1947 9.3
R2214 GND.n1946 GND.n1945 9.3
R2215 GND.n1956 GND.n1955 9.3
R2216 GND.n1955 GND.n1954 9.3
R2217 GND.n1965 GND.n1964 9.3
R2218 GND.n1964 GND.n1963 9.3
R2219 GND.n1969 GND.n1968 9.3
R2220 GND.n1938 GND.n1937 9.3
R2221 GND.n1937 GND.n1936 9.3
R2222 GND.n3229 GND.n3228 9.3
R2223 GND.n3210 GND.n3209 9.3
R2224 GND.n3208 GND.n3207 9.3
R2225 GND.n3231 GND.n3230 9.3
R2226 GND.n3218 GND.n3217 9.3
R2227 GND.n3217 GND.n3216 9.3
R2228 GND.n3227 GND.n3226 9.3
R2229 GND.n3226 GND.n3225 9.3
R2230 GND.n3206 GND.n3205 9.3
R2231 GND.n3189 GND.n3188 9.3
R2232 GND.n3170 GND.n3169 9.3
R2233 GND.n3168 GND.n3167 9.3
R2234 GND.n3178 GND.n3177 9.3
R2235 GND.n3177 GND.n3176 9.3
R2236 GND.n3187 GND.n3186 9.3
R2237 GND.n3186 GND.n3185 9.3
R2238 GND.n3191 GND.n3190 9.3
R2239 GND.n3160 GND.n3159 9.3
R2240 GND.n3159 GND.n3158 9.3
R2241 GND.n3148 GND.n3147 9.3
R2242 GND.n3129 GND.n3128 9.3
R2243 GND.n3127 GND.n3126 9.3
R2244 GND.n3150 GND.n3149 9.3
R2245 GND.n3137 GND.n3136 9.3
R2246 GND.n3136 GND.n3135 9.3
R2247 GND.n3146 GND.n3145 9.3
R2248 GND.n3145 GND.n3144 9.3
R2249 GND.n3125 GND.n3124 9.3
R2250 GND.n3108 GND.n3107 9.3
R2251 GND.n3089 GND.n3088 9.3
R2252 GND.n3087 GND.n3086 9.3
R2253 GND.n3097 GND.n3096 9.3
R2254 GND.n3096 GND.n3095 9.3
R2255 GND.n3106 GND.n3105 9.3
R2256 GND.n3105 GND.n3104 9.3
R2257 GND.n3110 GND.n3109 9.3
R2258 GND.n3079 GND.n3078 9.3
R2259 GND.n3078 GND.n3077 9.3
R2260 GND.n3067 GND.n3066 9.3
R2261 GND.n3048 GND.n3047 9.3
R2262 GND.n3046 GND.n3045 9.3
R2263 GND.n3069 GND.n3068 9.3
R2264 GND.n3056 GND.n3055 9.3
R2265 GND.n3055 GND.n3054 9.3
R2266 GND.n3065 GND.n3064 9.3
R2267 GND.n3064 GND.n3063 9.3
R2268 GND.n3044 GND.n3043 9.3
R2269 GND.n3027 GND.n3026 9.3
R2270 GND.n3008 GND.n3007 9.3
R2271 GND.n3006 GND.n3005 9.3
R2272 GND.n3016 GND.n3015 9.3
R2273 GND.n3015 GND.n3014 9.3
R2274 GND.n3025 GND.n3024 9.3
R2275 GND.n3024 GND.n3023 9.3
R2276 GND.n3029 GND.n3028 9.3
R2277 GND.n2998 GND.n2997 9.3
R2278 GND.n2997 GND.n2996 9.3
R2279 GND.n2986 GND.n2985 9.3
R2280 GND.n2967 GND.n2966 9.3
R2281 GND.n2965 GND.n2964 9.3
R2282 GND.n2988 GND.n2987 9.3
R2283 GND.n2975 GND.n2974 9.3
R2284 GND.n2974 GND.n2973 9.3
R2285 GND.n2984 GND.n2983 9.3
R2286 GND.n2983 GND.n2982 9.3
R2287 GND.n2963 GND.n2962 9.3
R2288 GND.n2946 GND.n2945 9.3
R2289 GND.n2927 GND.n2926 9.3
R2290 GND.n2925 GND.n2924 9.3
R2291 GND.n2935 GND.n2934 9.3
R2292 GND.n2934 GND.n2933 9.3
R2293 GND.n2944 GND.n2943 9.3
R2294 GND.n2943 GND.n2942 9.3
R2295 GND.n2948 GND.n2947 9.3
R2296 GND.n2917 GND.n2916 9.3
R2297 GND.n2916 GND.n2915 9.3
R2298 GND.n2905 GND.n2904 9.3
R2299 GND.n2886 GND.n2885 9.3
R2300 GND.n2884 GND.n2883 9.3
R2301 GND.n2907 GND.n2906 9.3
R2302 GND.n2894 GND.n2893 9.3
R2303 GND.n2893 GND.n2892 9.3
R2304 GND.n2903 GND.n2902 9.3
R2305 GND.n2902 GND.n2901 9.3
R2306 GND.n2882 GND.n2881 9.3
R2307 GND.n2865 GND.n2864 9.3
R2308 GND.n2846 GND.n2845 9.3
R2309 GND.n2844 GND.n2843 9.3
R2310 GND.n2854 GND.n2853 9.3
R2311 GND.n2853 GND.n2852 9.3
R2312 GND.n2863 GND.n2862 9.3
R2313 GND.n2862 GND.n2861 9.3
R2314 GND.n2867 GND.n2866 9.3
R2315 GND.n2836 GND.n2835 9.3
R2316 GND.n2835 GND.n2834 9.3
R2317 GND.n2824 GND.n2823 9.3
R2318 GND.n2805 GND.n2804 9.3
R2319 GND.n2803 GND.n2802 9.3
R2320 GND.n2826 GND.n2825 9.3
R2321 GND.n2813 GND.n2812 9.3
R2322 GND.n2812 GND.n2811 9.3
R2323 GND.n2822 GND.n2821 9.3
R2324 GND.n2821 GND.n2820 9.3
R2325 GND.n2801 GND.n2800 9.3
R2326 GND.n2784 GND.n2783 9.3
R2327 GND.n2765 GND.n2764 9.3
R2328 GND.n2763 GND.n2762 9.3
R2329 GND.n2773 GND.n2772 9.3
R2330 GND.n2772 GND.n2771 9.3
R2331 GND.n2782 GND.n2781 9.3
R2332 GND.n2781 GND.n2780 9.3
R2333 GND.n2786 GND.n2785 9.3
R2334 GND.n2755 GND.n2754 9.3
R2335 GND.n2754 GND.n2753 9.3
R2336 GND.n2743 GND.n2742 9.3
R2337 GND.n2724 GND.n2723 9.3
R2338 GND.n2722 GND.n2721 9.3
R2339 GND.n2745 GND.n2744 9.3
R2340 GND.n2732 GND.n2731 9.3
R2341 GND.n2731 GND.n2730 9.3
R2342 GND.n2741 GND.n2740 9.3
R2343 GND.n2740 GND.n2739 9.3
R2344 GND.n2720 GND.n2719 9.3
R2345 GND.n2703 GND.n2702 9.3
R2346 GND.n2684 GND.n2683 9.3
R2347 GND.n2682 GND.n2681 9.3
R2348 GND.n2692 GND.n2691 9.3
R2349 GND.n2691 GND.n2690 9.3
R2350 GND.n2701 GND.n2700 9.3
R2351 GND.n2700 GND.n2699 9.3
R2352 GND.n2705 GND.n2704 9.3
R2353 GND.n2674 GND.n2673 9.3
R2354 GND.n2673 GND.n2672 9.3
R2355 GND.n2662 GND.n2661 9.3
R2356 GND.n2643 GND.n2642 9.3
R2357 GND.n2641 GND.n2640 9.3
R2358 GND.n2664 GND.n2663 9.3
R2359 GND.n2651 GND.n2650 9.3
R2360 GND.n2650 GND.n2649 9.3
R2361 GND.n2660 GND.n2659 9.3
R2362 GND.n2659 GND.n2658 9.3
R2363 GND.n2639 GND.n2638 9.3
R2364 GND.n2622 GND.n2621 9.3
R2365 GND.n2603 GND.n2602 9.3
R2366 GND.n2601 GND.n2600 9.3
R2367 GND.n2611 GND.n2610 9.3
R2368 GND.n2610 GND.n2609 9.3
R2369 GND.n2620 GND.n2619 9.3
R2370 GND.n2619 GND.n2618 9.3
R2371 GND.n2624 GND.n2623 9.3
R2372 GND.n2593 GND.n2592 9.3
R2373 GND.n2592 GND.n2591 9.3
R2374 GND.n3884 GND.n3883 9.3
R2375 GND.n3865 GND.n3864 9.3
R2376 GND.n3863 GND.n3862 9.3
R2377 GND.n3886 GND.n3885 9.3
R2378 GND.n3873 GND.n3872 9.3
R2379 GND.n3872 GND.n3871 9.3
R2380 GND.n3882 GND.n3881 9.3
R2381 GND.n3881 GND.n3880 9.3
R2382 GND.n3861 GND.n3860 9.3
R2383 GND.n3844 GND.n3843 9.3
R2384 GND.n3825 GND.n3824 9.3
R2385 GND.n3823 GND.n3822 9.3
R2386 GND.n3833 GND.n3832 9.3
R2387 GND.n3832 GND.n3831 9.3
R2388 GND.n3842 GND.n3841 9.3
R2389 GND.n3841 GND.n3840 9.3
R2390 GND.n3846 GND.n3845 9.3
R2391 GND.n3815 GND.n3814 9.3
R2392 GND.n3814 GND.n3813 9.3
R2393 GND.n3803 GND.n3802 9.3
R2394 GND.n3784 GND.n3783 9.3
R2395 GND.n3782 GND.n3781 9.3
R2396 GND.n3805 GND.n3804 9.3
R2397 GND.n3792 GND.n3791 9.3
R2398 GND.n3791 GND.n3790 9.3
R2399 GND.n3801 GND.n3800 9.3
R2400 GND.n3800 GND.n3799 9.3
R2401 GND.n3780 GND.n3779 9.3
R2402 GND.n3763 GND.n3762 9.3
R2403 GND.n3744 GND.n3743 9.3
R2404 GND.n3742 GND.n3741 9.3
R2405 GND.n3752 GND.n3751 9.3
R2406 GND.n3751 GND.n3750 9.3
R2407 GND.n3761 GND.n3760 9.3
R2408 GND.n3760 GND.n3759 9.3
R2409 GND.n3765 GND.n3764 9.3
R2410 GND.n3734 GND.n3733 9.3
R2411 GND.n3733 GND.n3732 9.3
R2412 GND.n3722 GND.n3721 9.3
R2413 GND.n3703 GND.n3702 9.3
R2414 GND.n3701 GND.n3700 9.3
R2415 GND.n3724 GND.n3723 9.3
R2416 GND.n3711 GND.n3710 9.3
R2417 GND.n3710 GND.n3709 9.3
R2418 GND.n3720 GND.n3719 9.3
R2419 GND.n3719 GND.n3718 9.3
R2420 GND.n3699 GND.n3698 9.3
R2421 GND.n3682 GND.n3681 9.3
R2422 GND.n3663 GND.n3662 9.3
R2423 GND.n3661 GND.n3660 9.3
R2424 GND.n3671 GND.n3670 9.3
R2425 GND.n3670 GND.n3669 9.3
R2426 GND.n3680 GND.n3679 9.3
R2427 GND.n3679 GND.n3678 9.3
R2428 GND.n3684 GND.n3683 9.3
R2429 GND.n3653 GND.n3652 9.3
R2430 GND.n3652 GND.n3651 9.3
R2431 GND.n3641 GND.n3640 9.3
R2432 GND.n3622 GND.n3621 9.3
R2433 GND.n3620 GND.n3619 9.3
R2434 GND.n3643 GND.n3642 9.3
R2435 GND.n3630 GND.n3629 9.3
R2436 GND.n3629 GND.n3628 9.3
R2437 GND.n3639 GND.n3638 9.3
R2438 GND.n3638 GND.n3637 9.3
R2439 GND.n3618 GND.n3617 9.3
R2440 GND.n3601 GND.n3600 9.3
R2441 GND.n3582 GND.n3581 9.3
R2442 GND.n3580 GND.n3579 9.3
R2443 GND.n3590 GND.n3589 9.3
R2444 GND.n3589 GND.n3588 9.3
R2445 GND.n3599 GND.n3598 9.3
R2446 GND.n3598 GND.n3597 9.3
R2447 GND.n3603 GND.n3602 9.3
R2448 GND.n3572 GND.n3571 9.3
R2449 GND.n3571 GND.n3570 9.3
R2450 GND.n3560 GND.n3559 9.3
R2451 GND.n3541 GND.n3540 9.3
R2452 GND.n3539 GND.n3538 9.3
R2453 GND.n3562 GND.n3561 9.3
R2454 GND.n3549 GND.n3548 9.3
R2455 GND.n3548 GND.n3547 9.3
R2456 GND.n3558 GND.n3557 9.3
R2457 GND.n3557 GND.n3556 9.3
R2458 GND.n3537 GND.n3536 9.3
R2459 GND.n3520 GND.n3519 9.3
R2460 GND.n3501 GND.n3500 9.3
R2461 GND.n3499 GND.n3498 9.3
R2462 GND.n3509 GND.n3508 9.3
R2463 GND.n3508 GND.n3507 9.3
R2464 GND.n3518 GND.n3517 9.3
R2465 GND.n3517 GND.n3516 9.3
R2466 GND.n3522 GND.n3521 9.3
R2467 GND.n3491 GND.n3490 9.3
R2468 GND.n3490 GND.n3489 9.3
R2469 GND.n3479 GND.n3478 9.3
R2470 GND.n3460 GND.n3459 9.3
R2471 GND.n3458 GND.n3457 9.3
R2472 GND.n3481 GND.n3480 9.3
R2473 GND.n3468 GND.n3467 9.3
R2474 GND.n3467 GND.n3466 9.3
R2475 GND.n3477 GND.n3476 9.3
R2476 GND.n3476 GND.n3475 9.3
R2477 GND.n3456 GND.n3455 9.3
R2478 GND.n3439 GND.n3438 9.3
R2479 GND.n3420 GND.n3419 9.3
R2480 GND.n3418 GND.n3417 9.3
R2481 GND.n3428 GND.n3427 9.3
R2482 GND.n3427 GND.n3426 9.3
R2483 GND.n3437 GND.n3436 9.3
R2484 GND.n3436 GND.n3435 9.3
R2485 GND.n3441 GND.n3440 9.3
R2486 GND.n3410 GND.n3409 9.3
R2487 GND.n3409 GND.n3408 9.3
R2488 GND.n3398 GND.n3397 9.3
R2489 GND.n3379 GND.n3378 9.3
R2490 GND.n3377 GND.n3376 9.3
R2491 GND.n3400 GND.n3399 9.3
R2492 GND.n3387 GND.n3386 9.3
R2493 GND.n3386 GND.n3385 9.3
R2494 GND.n3396 GND.n3395 9.3
R2495 GND.n3395 GND.n3394 9.3
R2496 GND.n3375 GND.n3374 9.3
R2497 GND.n3358 GND.n3357 9.3
R2498 GND.n3339 GND.n3338 9.3
R2499 GND.n3337 GND.n3336 9.3
R2500 GND.n3347 GND.n3346 9.3
R2501 GND.n3346 GND.n3345 9.3
R2502 GND.n3356 GND.n3355 9.3
R2503 GND.n3355 GND.n3354 9.3
R2504 GND.n3360 GND.n3359 9.3
R2505 GND.n3329 GND.n3328 9.3
R2506 GND.n3328 GND.n3327 9.3
R2507 GND.n3317 GND.n3316 9.3
R2508 GND.n3298 GND.n3297 9.3
R2509 GND.n3296 GND.n3295 9.3
R2510 GND.n3319 GND.n3318 9.3
R2511 GND.n3306 GND.n3305 9.3
R2512 GND.n3305 GND.n3304 9.3
R2513 GND.n3315 GND.n3314 9.3
R2514 GND.n3314 GND.n3313 9.3
R2515 GND.n3294 GND.n3293 9.3
R2516 GND.n3277 GND.n3276 9.3
R2517 GND.n3258 GND.n3257 9.3
R2518 GND.n3256 GND.n3255 9.3
R2519 GND.n3266 GND.n3265 9.3
R2520 GND.n3265 GND.n3264 9.3
R2521 GND.n3275 GND.n3274 9.3
R2522 GND.n3274 GND.n3273 9.3
R2523 GND.n3279 GND.n3278 9.3
R2524 GND.n3248 GND.n3247 9.3
R2525 GND.n3247 GND.n3246 9.3
R2526 GND.n4539 GND.n4538 9.3
R2527 GND.n4520 GND.n4519 9.3
R2528 GND.n4518 GND.n4517 9.3
R2529 GND.n4541 GND.n4540 9.3
R2530 GND.n4528 GND.n4527 9.3
R2531 GND.n4527 GND.n4526 9.3
R2532 GND.n4537 GND.n4536 9.3
R2533 GND.n4536 GND.n4535 9.3
R2534 GND.n4516 GND.n4515 9.3
R2535 GND.n4499 GND.n4498 9.3
R2536 GND.n4480 GND.n4479 9.3
R2537 GND.n4478 GND.n4477 9.3
R2538 GND.n4488 GND.n4487 9.3
R2539 GND.n4487 GND.n4486 9.3
R2540 GND.n4497 GND.n4496 9.3
R2541 GND.n4496 GND.n4495 9.3
R2542 GND.n4501 GND.n4500 9.3
R2543 GND.n4470 GND.n4469 9.3
R2544 GND.n4469 GND.n4468 9.3
R2545 GND.n4458 GND.n4457 9.3
R2546 GND.n4439 GND.n4438 9.3
R2547 GND.n4437 GND.n4436 9.3
R2548 GND.n4460 GND.n4459 9.3
R2549 GND.n4447 GND.n4446 9.3
R2550 GND.n4446 GND.n4445 9.3
R2551 GND.n4456 GND.n4455 9.3
R2552 GND.n4455 GND.n4454 9.3
R2553 GND.n4435 GND.n4434 9.3
R2554 GND.n4418 GND.n4417 9.3
R2555 GND.n4399 GND.n4398 9.3
R2556 GND.n4397 GND.n4396 9.3
R2557 GND.n4407 GND.n4406 9.3
R2558 GND.n4406 GND.n4405 9.3
R2559 GND.n4416 GND.n4415 9.3
R2560 GND.n4415 GND.n4414 9.3
R2561 GND.n4420 GND.n4419 9.3
R2562 GND.n4389 GND.n4388 9.3
R2563 GND.n4388 GND.n4387 9.3
R2564 GND.n4377 GND.n4376 9.3
R2565 GND.n4358 GND.n4357 9.3
R2566 GND.n4356 GND.n4355 9.3
R2567 GND.n4379 GND.n4378 9.3
R2568 GND.n4366 GND.n4365 9.3
R2569 GND.n4365 GND.n4364 9.3
R2570 GND.n4375 GND.n4374 9.3
R2571 GND.n4374 GND.n4373 9.3
R2572 GND.n4354 GND.n4353 9.3
R2573 GND.n4337 GND.n4336 9.3
R2574 GND.n4318 GND.n4317 9.3
R2575 GND.n4316 GND.n4315 9.3
R2576 GND.n4326 GND.n4325 9.3
R2577 GND.n4325 GND.n4324 9.3
R2578 GND.n4335 GND.n4334 9.3
R2579 GND.n4334 GND.n4333 9.3
R2580 GND.n4339 GND.n4338 9.3
R2581 GND.n4308 GND.n4307 9.3
R2582 GND.n4307 GND.n4306 9.3
R2583 GND.n4296 GND.n4295 9.3
R2584 GND.n4277 GND.n4276 9.3
R2585 GND.n4275 GND.n4274 9.3
R2586 GND.n4298 GND.n4297 9.3
R2587 GND.n4285 GND.n4284 9.3
R2588 GND.n4284 GND.n4283 9.3
R2589 GND.n4294 GND.n4293 9.3
R2590 GND.n4293 GND.n4292 9.3
R2591 GND.n4273 GND.n4272 9.3
R2592 GND.n4256 GND.n4255 9.3
R2593 GND.n4237 GND.n4236 9.3
R2594 GND.n4235 GND.n4234 9.3
R2595 GND.n4245 GND.n4244 9.3
R2596 GND.n4244 GND.n4243 9.3
R2597 GND.n4254 GND.n4253 9.3
R2598 GND.n4253 GND.n4252 9.3
R2599 GND.n4258 GND.n4257 9.3
R2600 GND.n4227 GND.n4226 9.3
R2601 GND.n4226 GND.n4225 9.3
R2602 GND.n4215 GND.n4214 9.3
R2603 GND.n4196 GND.n4195 9.3
R2604 GND.n4194 GND.n4193 9.3
R2605 GND.n4217 GND.n4216 9.3
R2606 GND.n4204 GND.n4203 9.3
R2607 GND.n4203 GND.n4202 9.3
R2608 GND.n4213 GND.n4212 9.3
R2609 GND.n4212 GND.n4211 9.3
R2610 GND.n4192 GND.n4191 9.3
R2611 GND.n4175 GND.n4174 9.3
R2612 GND.n4156 GND.n4155 9.3
R2613 GND.n4154 GND.n4153 9.3
R2614 GND.n4164 GND.n4163 9.3
R2615 GND.n4163 GND.n4162 9.3
R2616 GND.n4173 GND.n4172 9.3
R2617 GND.n4172 GND.n4171 9.3
R2618 GND.n4177 GND.n4176 9.3
R2619 GND.n4146 GND.n4145 9.3
R2620 GND.n4145 GND.n4144 9.3
R2621 GND.n4134 GND.n4133 9.3
R2622 GND.n4115 GND.n4114 9.3
R2623 GND.n4113 GND.n4112 9.3
R2624 GND.n4136 GND.n4135 9.3
R2625 GND.n4123 GND.n4122 9.3
R2626 GND.n4122 GND.n4121 9.3
R2627 GND.n4132 GND.n4131 9.3
R2628 GND.n4131 GND.n4130 9.3
R2629 GND.n4111 GND.n4110 9.3
R2630 GND.n4094 GND.n4093 9.3
R2631 GND.n4075 GND.n4074 9.3
R2632 GND.n4073 GND.n4072 9.3
R2633 GND.n4083 GND.n4082 9.3
R2634 GND.n4082 GND.n4081 9.3
R2635 GND.n4092 GND.n4091 9.3
R2636 GND.n4091 GND.n4090 9.3
R2637 GND.n4096 GND.n4095 9.3
R2638 GND.n4065 GND.n4064 9.3
R2639 GND.n4064 GND.n4063 9.3
R2640 GND.n4053 GND.n4052 9.3
R2641 GND.n4034 GND.n4033 9.3
R2642 GND.n4032 GND.n4031 9.3
R2643 GND.n4055 GND.n4054 9.3
R2644 GND.n4042 GND.n4041 9.3
R2645 GND.n4041 GND.n4040 9.3
R2646 GND.n4051 GND.n4050 9.3
R2647 GND.n4050 GND.n4049 9.3
R2648 GND.n4030 GND.n4029 9.3
R2649 GND.n4013 GND.n4012 9.3
R2650 GND.n3994 GND.n3993 9.3
R2651 GND.n3992 GND.n3991 9.3
R2652 GND.n4002 GND.n4001 9.3
R2653 GND.n4001 GND.n4000 9.3
R2654 GND.n4011 GND.n4010 9.3
R2655 GND.n4010 GND.n4009 9.3
R2656 GND.n4015 GND.n4014 9.3
R2657 GND.n3984 GND.n3983 9.3
R2658 GND.n3983 GND.n3982 9.3
R2659 GND.n3972 GND.n3971 9.3
R2660 GND.n3953 GND.n3952 9.3
R2661 GND.n3951 GND.n3950 9.3
R2662 GND.n3974 GND.n3973 9.3
R2663 GND.n3961 GND.n3960 9.3
R2664 GND.n3960 GND.n3959 9.3
R2665 GND.n3970 GND.n3969 9.3
R2666 GND.n3969 GND.n3968 9.3
R2667 GND.n3949 GND.n3948 9.3
R2668 GND.n3932 GND.n3931 9.3
R2669 GND.n3913 GND.n3912 9.3
R2670 GND.n3911 GND.n3910 9.3
R2671 GND.n3921 GND.n3920 9.3
R2672 GND.n3920 GND.n3919 9.3
R2673 GND.n3930 GND.n3929 9.3
R2674 GND.n3929 GND.n3928 9.3
R2675 GND.n3934 GND.n3933 9.3
R2676 GND.n3903 GND.n3902 9.3
R2677 GND.n3902 GND.n3901 9.3
R2678 GND.n5204 GND.n5203 9.3
R2679 GND.n5185 GND.n5184 9.3
R2680 GND.n5183 GND.n5182 9.3
R2681 GND.n5206 GND.n5205 9.3
R2682 GND.n5193 GND.n5192 9.3
R2683 GND.n5192 GND.n5191 9.3
R2684 GND.n5202 GND.n5201 9.3
R2685 GND.n5201 GND.n5200 9.3
R2686 GND.n5181 GND.n5180 9.3
R2687 GND.n5164 GND.n5163 9.3
R2688 GND.n5145 GND.n5144 9.3
R2689 GND.n5143 GND.n5142 9.3
R2690 GND.n5153 GND.n5152 9.3
R2691 GND.n5152 GND.n5151 9.3
R2692 GND.n5162 GND.n5161 9.3
R2693 GND.n5161 GND.n5160 9.3
R2694 GND.n5166 GND.n5165 9.3
R2695 GND.n5135 GND.n5134 9.3
R2696 GND.n5134 GND.n5133 9.3
R2697 GND.n5123 GND.n5122 9.3
R2698 GND.n5104 GND.n5103 9.3
R2699 GND.n5102 GND.n5101 9.3
R2700 GND.n5125 GND.n5124 9.3
R2701 GND.n5112 GND.n5111 9.3
R2702 GND.n5111 GND.n5110 9.3
R2703 GND.n5121 GND.n5120 9.3
R2704 GND.n5120 GND.n5119 9.3
R2705 GND.n5100 GND.n5099 9.3
R2706 GND.n5083 GND.n5082 9.3
R2707 GND.n5064 GND.n5063 9.3
R2708 GND.n5062 GND.n5061 9.3
R2709 GND.n5072 GND.n5071 9.3
R2710 GND.n5071 GND.n5070 9.3
R2711 GND.n5081 GND.n5080 9.3
R2712 GND.n5080 GND.n5079 9.3
R2713 GND.n5085 GND.n5084 9.3
R2714 GND.n5054 GND.n5053 9.3
R2715 GND.n5053 GND.n5052 9.3
R2716 GND.n5042 GND.n5041 9.3
R2717 GND.n5023 GND.n5022 9.3
R2718 GND.n5021 GND.n5020 9.3
R2719 GND.n5044 GND.n5043 9.3
R2720 GND.n5031 GND.n5030 9.3
R2721 GND.n5030 GND.n5029 9.3
R2722 GND.n5040 GND.n5039 9.3
R2723 GND.n5039 GND.n5038 9.3
R2724 GND.n5019 GND.n5018 9.3
R2725 GND.n5002 GND.n5001 9.3
R2726 GND.n4983 GND.n4982 9.3
R2727 GND.n4981 GND.n4980 9.3
R2728 GND.n4991 GND.n4990 9.3
R2729 GND.n4990 GND.n4989 9.3
R2730 GND.n5000 GND.n4999 9.3
R2731 GND.n4999 GND.n4998 9.3
R2732 GND.n5004 GND.n5003 9.3
R2733 GND.n4973 GND.n4972 9.3
R2734 GND.n4972 GND.n4971 9.3
R2735 GND.n4961 GND.n4960 9.3
R2736 GND.n4942 GND.n4941 9.3
R2737 GND.n4940 GND.n4939 9.3
R2738 GND.n4963 GND.n4962 9.3
R2739 GND.n4950 GND.n4949 9.3
R2740 GND.n4949 GND.n4948 9.3
R2741 GND.n4959 GND.n4958 9.3
R2742 GND.n4958 GND.n4957 9.3
R2743 GND.n4938 GND.n4937 9.3
R2744 GND.n4921 GND.n4920 9.3
R2745 GND.n4902 GND.n4901 9.3
R2746 GND.n4900 GND.n4899 9.3
R2747 GND.n4910 GND.n4909 9.3
R2748 GND.n4909 GND.n4908 9.3
R2749 GND.n4919 GND.n4918 9.3
R2750 GND.n4918 GND.n4917 9.3
R2751 GND.n4923 GND.n4922 9.3
R2752 GND.n4892 GND.n4891 9.3
R2753 GND.n4891 GND.n4890 9.3
R2754 GND.n4880 GND.n4879 9.3
R2755 GND.n4861 GND.n4860 9.3
R2756 GND.n4859 GND.n4858 9.3
R2757 GND.n4882 GND.n4881 9.3
R2758 GND.n4869 GND.n4868 9.3
R2759 GND.n4868 GND.n4867 9.3
R2760 GND.n4878 GND.n4877 9.3
R2761 GND.n4877 GND.n4876 9.3
R2762 GND.n4857 GND.n4856 9.3
R2763 GND.n4840 GND.n4839 9.3
R2764 GND.n4821 GND.n4820 9.3
R2765 GND.n4819 GND.n4818 9.3
R2766 GND.n4829 GND.n4828 9.3
R2767 GND.n4828 GND.n4827 9.3
R2768 GND.n4838 GND.n4837 9.3
R2769 GND.n4837 GND.n4836 9.3
R2770 GND.n4842 GND.n4841 9.3
R2771 GND.n4811 GND.n4810 9.3
R2772 GND.n4810 GND.n4809 9.3
R2773 GND.n4799 GND.n4798 9.3
R2774 GND.n4780 GND.n4779 9.3
R2775 GND.n4778 GND.n4777 9.3
R2776 GND.n4801 GND.n4800 9.3
R2777 GND.n4788 GND.n4787 9.3
R2778 GND.n4787 GND.n4786 9.3
R2779 GND.n4797 GND.n4796 9.3
R2780 GND.n4796 GND.n4795 9.3
R2781 GND.n4776 GND.n4775 9.3
R2782 GND.n4759 GND.n4758 9.3
R2783 GND.n4740 GND.n4739 9.3
R2784 GND.n4738 GND.n4737 9.3
R2785 GND.n4748 GND.n4747 9.3
R2786 GND.n4747 GND.n4746 9.3
R2787 GND.n4757 GND.n4756 9.3
R2788 GND.n4756 GND.n4755 9.3
R2789 GND.n4761 GND.n4760 9.3
R2790 GND.n4730 GND.n4729 9.3
R2791 GND.n4729 GND.n4728 9.3
R2792 GND.n4718 GND.n4717 9.3
R2793 GND.n4699 GND.n4698 9.3
R2794 GND.n4697 GND.n4696 9.3
R2795 GND.n4720 GND.n4719 9.3
R2796 GND.n4707 GND.n4706 9.3
R2797 GND.n4706 GND.n4705 9.3
R2798 GND.n4716 GND.n4715 9.3
R2799 GND.n4715 GND.n4714 9.3
R2800 GND.n4695 GND.n4694 9.3
R2801 GND.n4678 GND.n4677 9.3
R2802 GND.n4659 GND.n4658 9.3
R2803 GND.n4657 GND.n4656 9.3
R2804 GND.n4667 GND.n4666 9.3
R2805 GND.n4666 GND.n4665 9.3
R2806 GND.n4676 GND.n4675 9.3
R2807 GND.n4675 GND.n4674 9.3
R2808 GND.n4680 GND.n4679 9.3
R2809 GND.n4649 GND.n4648 9.3
R2810 GND.n4648 GND.n4647 9.3
R2811 GND.n4637 GND.n4636 9.3
R2812 GND.n4618 GND.n4617 9.3
R2813 GND.n4616 GND.n4615 9.3
R2814 GND.n4639 GND.n4638 9.3
R2815 GND.n4626 GND.n4625 9.3
R2816 GND.n4625 GND.n4624 9.3
R2817 GND.n4635 GND.n4634 9.3
R2818 GND.n4634 GND.n4633 9.3
R2819 GND.n4614 GND.n4613 9.3
R2820 GND.n4597 GND.n4596 9.3
R2821 GND.n4578 GND.n4577 9.3
R2822 GND.n4576 GND.n4575 9.3
R2823 GND.n4586 GND.n4585 9.3
R2824 GND.n4585 GND.n4584 9.3
R2825 GND.n4595 GND.n4594 9.3
R2826 GND.n4594 GND.n4593 9.3
R2827 GND.n4599 GND.n4598 9.3
R2828 GND.n4568 GND.n4567 9.3
R2829 GND.n4567 GND.n4566 9.3
R2830 GND.n227 GND.n226 9.001
R2831 GND.n146 GND.n145 9.001
R2832 GND.n562 GND.n561 9.001
R2833 GND.n481 GND.n480 9.001
R2834 GND.n400 GND.n399 9.001
R2835 GND.n319 GND.n318 9.001
R2836 GND.n1223 GND.n1222 9.001
R2837 GND.n1142 GND.n1141 9.001
R2838 GND.n1061 GND.n1060 9.001
R2839 GND.n980 GND.n979 9.001
R2840 GND.n899 GND.n898 9.001
R2841 GND.n818 GND.n817 9.001
R2842 GND.n737 GND.n736 9.001
R2843 GND.n656 GND.n655 9.001
R2844 GND.n1878 GND.n1877 9.001
R2845 GND.n1797 GND.n1796 9.001
R2846 GND.n1716 GND.n1715 9.001
R2847 GND.n1635 GND.n1634 9.001
R2848 GND.n1554 GND.n1553 9.001
R2849 GND.n1473 GND.n1472 9.001
R2850 GND.n1392 GND.n1391 9.001
R2851 GND.n1311 GND.n1310 9.001
R2852 GND.n2543 GND.n2542 9.001
R2853 GND.n2462 GND.n2461 9.001
R2854 GND.n2381 GND.n2380 9.001
R2855 GND.n2300 GND.n2299 9.001
R2856 GND.n2219 GND.n2218 9.001
R2857 GND.n2138 GND.n2137 9.001
R2858 GND.n2057 GND.n2056 9.001
R2859 GND.n1976 GND.n1975 9.001
R2860 GND.n3198 GND.n3197 9.001
R2861 GND.n3117 GND.n3116 9.001
R2862 GND.n3036 GND.n3035 9.001
R2863 GND.n2955 GND.n2954 9.001
R2864 GND.n2874 GND.n2873 9.001
R2865 GND.n2793 GND.n2792 9.001
R2866 GND.n2712 GND.n2711 9.001
R2867 GND.n2631 GND.n2630 9.001
R2868 GND.n3853 GND.n3852 9.001
R2869 GND.n3772 GND.n3771 9.001
R2870 GND.n3691 GND.n3690 9.001
R2871 GND.n3610 GND.n3609 9.001
R2872 GND.n3529 GND.n3528 9.001
R2873 GND.n3448 GND.n3447 9.001
R2874 GND.n3367 GND.n3366 9.001
R2875 GND.n3286 GND.n3285 9.001
R2876 GND.n4508 GND.n4507 9.001
R2877 GND.n4427 GND.n4426 9.001
R2878 GND.n4346 GND.n4345 9.001
R2879 GND.n4265 GND.n4264 9.001
R2880 GND.n4184 GND.n4183 9.001
R2881 GND.n4103 GND.n4102 9.001
R2882 GND.n4022 GND.n4021 9.001
R2883 GND.n3941 GND.n3940 9.001
R2884 GND.n5173 GND.n5172 9.001
R2885 GND.n5092 GND.n5091 9.001
R2886 GND.n5011 GND.n5010 9.001
R2887 GND.n4930 GND.n4929 9.001
R2888 GND.n4849 GND.n4848 9.001
R2889 GND.n4768 GND.n4767 9.001
R2890 GND.n4687 GND.n4686 9.001
R2891 GND.n4606 GND.n4605 9.001
R2892 GND.n69 GND.n68 6.023
R2893 GND.n77 GND.n76 6.023
R2894 GND.n29 GND.n28 6.023
R2895 GND.n37 GND.n36 6.023
R2896 GND.n241 GND.n240 6.023
R2897 GND.n249 GND.n248 6.023
R2898 GND.n201 GND.n200 6.023
R2899 GND.n209 GND.n208 6.023
R2900 GND.n160 GND.n159 6.023
R2901 GND.n168 GND.n167 6.023
R2902 GND.n120 GND.n119 6.023
R2903 GND.n128 GND.n127 6.023
R2904 GND.n576 GND.n575 6.023
R2905 GND.n584 GND.n583 6.023
R2906 GND.n536 GND.n535 6.023
R2907 GND.n544 GND.n543 6.023
R2908 GND.n495 GND.n494 6.023
R2909 GND.n503 GND.n502 6.023
R2910 GND.n455 GND.n454 6.023
R2911 GND.n463 GND.n462 6.023
R2912 GND.n414 GND.n413 6.023
R2913 GND.n422 GND.n421 6.023
R2914 GND.n374 GND.n373 6.023
R2915 GND.n382 GND.n381 6.023
R2916 GND.n333 GND.n332 6.023
R2917 GND.n341 GND.n340 6.023
R2918 GND.n293 GND.n292 6.023
R2919 GND.n301 GND.n300 6.023
R2920 GND.n1237 GND.n1236 6.023
R2921 GND.n1245 GND.n1244 6.023
R2922 GND.n1197 GND.n1196 6.023
R2923 GND.n1205 GND.n1204 6.023
R2924 GND.n1156 GND.n1155 6.023
R2925 GND.n1164 GND.n1163 6.023
R2926 GND.n1116 GND.n1115 6.023
R2927 GND.n1124 GND.n1123 6.023
R2928 GND.n1075 GND.n1074 6.023
R2929 GND.n1083 GND.n1082 6.023
R2930 GND.n1035 GND.n1034 6.023
R2931 GND.n1043 GND.n1042 6.023
R2932 GND.n994 GND.n993 6.023
R2933 GND.n1002 GND.n1001 6.023
R2934 GND.n954 GND.n953 6.023
R2935 GND.n962 GND.n961 6.023
R2936 GND.n913 GND.n912 6.023
R2937 GND.n921 GND.n920 6.023
R2938 GND.n873 GND.n872 6.023
R2939 GND.n881 GND.n880 6.023
R2940 GND.n832 GND.n831 6.023
R2941 GND.n840 GND.n839 6.023
R2942 GND.n792 GND.n791 6.023
R2943 GND.n800 GND.n799 6.023
R2944 GND.n751 GND.n750 6.023
R2945 GND.n759 GND.n758 6.023
R2946 GND.n711 GND.n710 6.023
R2947 GND.n719 GND.n718 6.023
R2948 GND.n670 GND.n669 6.023
R2949 GND.n678 GND.n677 6.023
R2950 GND.n630 GND.n629 6.023
R2951 GND.n638 GND.n637 6.023
R2952 GND.n1892 GND.n1891 6.023
R2953 GND.n1900 GND.n1899 6.023
R2954 GND.n1852 GND.n1851 6.023
R2955 GND.n1860 GND.n1859 6.023
R2956 GND.n1811 GND.n1810 6.023
R2957 GND.n1819 GND.n1818 6.023
R2958 GND.n1771 GND.n1770 6.023
R2959 GND.n1779 GND.n1778 6.023
R2960 GND.n1730 GND.n1729 6.023
R2961 GND.n1738 GND.n1737 6.023
R2962 GND.n1690 GND.n1689 6.023
R2963 GND.n1698 GND.n1697 6.023
R2964 GND.n1649 GND.n1648 6.023
R2965 GND.n1657 GND.n1656 6.023
R2966 GND.n1609 GND.n1608 6.023
R2967 GND.n1617 GND.n1616 6.023
R2968 GND.n1568 GND.n1567 6.023
R2969 GND.n1576 GND.n1575 6.023
R2970 GND.n1528 GND.n1527 6.023
R2971 GND.n1536 GND.n1535 6.023
R2972 GND.n1487 GND.n1486 6.023
R2973 GND.n1495 GND.n1494 6.023
R2974 GND.n1447 GND.n1446 6.023
R2975 GND.n1455 GND.n1454 6.023
R2976 GND.n1406 GND.n1405 6.023
R2977 GND.n1414 GND.n1413 6.023
R2978 GND.n1366 GND.n1365 6.023
R2979 GND.n1374 GND.n1373 6.023
R2980 GND.n1325 GND.n1324 6.023
R2981 GND.n1333 GND.n1332 6.023
R2982 GND.n1285 GND.n1284 6.023
R2983 GND.n1293 GND.n1292 6.023
R2984 GND.n2557 GND.n2556 6.023
R2985 GND.n2565 GND.n2564 6.023
R2986 GND.n2517 GND.n2516 6.023
R2987 GND.n2525 GND.n2524 6.023
R2988 GND.n2476 GND.n2475 6.023
R2989 GND.n2484 GND.n2483 6.023
R2990 GND.n2436 GND.n2435 6.023
R2991 GND.n2444 GND.n2443 6.023
R2992 GND.n2395 GND.n2394 6.023
R2993 GND.n2403 GND.n2402 6.023
R2994 GND.n2355 GND.n2354 6.023
R2995 GND.n2363 GND.n2362 6.023
R2996 GND.n2314 GND.n2313 6.023
R2997 GND.n2322 GND.n2321 6.023
R2998 GND.n2274 GND.n2273 6.023
R2999 GND.n2282 GND.n2281 6.023
R3000 GND.n2233 GND.n2232 6.023
R3001 GND.n2241 GND.n2240 6.023
R3002 GND.n2193 GND.n2192 6.023
R3003 GND.n2201 GND.n2200 6.023
R3004 GND.n2152 GND.n2151 6.023
R3005 GND.n2160 GND.n2159 6.023
R3006 GND.n2112 GND.n2111 6.023
R3007 GND.n2120 GND.n2119 6.023
R3008 GND.n2071 GND.n2070 6.023
R3009 GND.n2079 GND.n2078 6.023
R3010 GND.n2031 GND.n2030 6.023
R3011 GND.n2039 GND.n2038 6.023
R3012 GND.n1990 GND.n1989 6.023
R3013 GND.n1998 GND.n1997 6.023
R3014 GND.n1950 GND.n1949 6.023
R3015 GND.n1958 GND.n1957 6.023
R3016 GND.n3212 GND.n3211 6.023
R3017 GND.n3220 GND.n3219 6.023
R3018 GND.n3172 GND.n3171 6.023
R3019 GND.n3180 GND.n3179 6.023
R3020 GND.n3131 GND.n3130 6.023
R3021 GND.n3139 GND.n3138 6.023
R3022 GND.n3091 GND.n3090 6.023
R3023 GND.n3099 GND.n3098 6.023
R3024 GND.n3050 GND.n3049 6.023
R3025 GND.n3058 GND.n3057 6.023
R3026 GND.n3010 GND.n3009 6.023
R3027 GND.n3018 GND.n3017 6.023
R3028 GND.n2969 GND.n2968 6.023
R3029 GND.n2977 GND.n2976 6.023
R3030 GND.n2929 GND.n2928 6.023
R3031 GND.n2937 GND.n2936 6.023
R3032 GND.n2888 GND.n2887 6.023
R3033 GND.n2896 GND.n2895 6.023
R3034 GND.n2848 GND.n2847 6.023
R3035 GND.n2856 GND.n2855 6.023
R3036 GND.n2807 GND.n2806 6.023
R3037 GND.n2815 GND.n2814 6.023
R3038 GND.n2767 GND.n2766 6.023
R3039 GND.n2775 GND.n2774 6.023
R3040 GND.n2726 GND.n2725 6.023
R3041 GND.n2734 GND.n2733 6.023
R3042 GND.n2686 GND.n2685 6.023
R3043 GND.n2694 GND.n2693 6.023
R3044 GND.n2645 GND.n2644 6.023
R3045 GND.n2653 GND.n2652 6.023
R3046 GND.n2605 GND.n2604 6.023
R3047 GND.n2613 GND.n2612 6.023
R3048 GND.n3867 GND.n3866 6.023
R3049 GND.n3875 GND.n3874 6.023
R3050 GND.n3827 GND.n3826 6.023
R3051 GND.n3835 GND.n3834 6.023
R3052 GND.n3786 GND.n3785 6.023
R3053 GND.n3794 GND.n3793 6.023
R3054 GND.n3746 GND.n3745 6.023
R3055 GND.n3754 GND.n3753 6.023
R3056 GND.n3705 GND.n3704 6.023
R3057 GND.n3713 GND.n3712 6.023
R3058 GND.n3665 GND.n3664 6.023
R3059 GND.n3673 GND.n3672 6.023
R3060 GND.n3624 GND.n3623 6.023
R3061 GND.n3632 GND.n3631 6.023
R3062 GND.n3584 GND.n3583 6.023
R3063 GND.n3592 GND.n3591 6.023
R3064 GND.n3543 GND.n3542 6.023
R3065 GND.n3551 GND.n3550 6.023
R3066 GND.n3503 GND.n3502 6.023
R3067 GND.n3511 GND.n3510 6.023
R3068 GND.n3462 GND.n3461 6.023
R3069 GND.n3470 GND.n3469 6.023
R3070 GND.n3422 GND.n3421 6.023
R3071 GND.n3430 GND.n3429 6.023
R3072 GND.n3381 GND.n3380 6.023
R3073 GND.n3389 GND.n3388 6.023
R3074 GND.n3341 GND.n3340 6.023
R3075 GND.n3349 GND.n3348 6.023
R3076 GND.n3300 GND.n3299 6.023
R3077 GND.n3308 GND.n3307 6.023
R3078 GND.n3260 GND.n3259 6.023
R3079 GND.n3268 GND.n3267 6.023
R3080 GND.n4522 GND.n4521 6.023
R3081 GND.n4530 GND.n4529 6.023
R3082 GND.n4482 GND.n4481 6.023
R3083 GND.n4490 GND.n4489 6.023
R3084 GND.n4441 GND.n4440 6.023
R3085 GND.n4449 GND.n4448 6.023
R3086 GND.n4401 GND.n4400 6.023
R3087 GND.n4409 GND.n4408 6.023
R3088 GND.n4360 GND.n4359 6.023
R3089 GND.n4368 GND.n4367 6.023
R3090 GND.n4320 GND.n4319 6.023
R3091 GND.n4328 GND.n4327 6.023
R3092 GND.n4279 GND.n4278 6.023
R3093 GND.n4287 GND.n4286 6.023
R3094 GND.n4239 GND.n4238 6.023
R3095 GND.n4247 GND.n4246 6.023
R3096 GND.n4198 GND.n4197 6.023
R3097 GND.n4206 GND.n4205 6.023
R3098 GND.n4158 GND.n4157 6.023
R3099 GND.n4166 GND.n4165 6.023
R3100 GND.n4117 GND.n4116 6.023
R3101 GND.n4125 GND.n4124 6.023
R3102 GND.n4077 GND.n4076 6.023
R3103 GND.n4085 GND.n4084 6.023
R3104 GND.n4036 GND.n4035 6.023
R3105 GND.n4044 GND.n4043 6.023
R3106 GND.n3996 GND.n3995 6.023
R3107 GND.n4004 GND.n4003 6.023
R3108 GND.n3955 GND.n3954 6.023
R3109 GND.n3963 GND.n3962 6.023
R3110 GND.n3915 GND.n3914 6.023
R3111 GND.n3923 GND.n3922 6.023
R3112 GND.n5187 GND.n5186 6.023
R3113 GND.n5195 GND.n5194 6.023
R3114 GND.n5147 GND.n5146 6.023
R3115 GND.n5155 GND.n5154 6.023
R3116 GND.n5106 GND.n5105 6.023
R3117 GND.n5114 GND.n5113 6.023
R3118 GND.n5066 GND.n5065 6.023
R3119 GND.n5074 GND.n5073 6.023
R3120 GND.n5025 GND.n5024 6.023
R3121 GND.n5033 GND.n5032 6.023
R3122 GND.n4985 GND.n4984 6.023
R3123 GND.n4993 GND.n4992 6.023
R3124 GND.n4944 GND.n4943 6.023
R3125 GND.n4952 GND.n4951 6.023
R3126 GND.n4904 GND.n4903 6.023
R3127 GND.n4912 GND.n4911 6.023
R3128 GND.n4863 GND.n4862 6.023
R3129 GND.n4871 GND.n4870 6.023
R3130 GND.n4823 GND.n4822 6.023
R3131 GND.n4831 GND.n4830 6.023
R3132 GND.n4782 GND.n4781 6.023
R3133 GND.n4790 GND.n4789 6.023
R3134 GND.n4742 GND.n4741 6.023
R3135 GND.n4750 GND.n4749 6.023
R3136 GND.n4701 GND.n4700 6.023
R3137 GND.n4709 GND.n4708 6.023
R3138 GND.n4661 GND.n4660 6.023
R3139 GND.n4669 GND.n4668 6.023
R3140 GND.n4620 GND.n4619 6.023
R3141 GND.n4628 GND.n4627 6.023
R3142 GND.n4580 GND.n4579 6.023
R3143 GND.n4588 GND.n4587 6.023
R3144 GND.n59 GND.n58 5.27
R3145 GND.n51 GND.n50 5.27
R3146 GND.n19 GND.n18 5.27
R3147 GND.n11 GND.n10 5.27
R3148 GND.n230 GND.n229 5.27
R3149 GND.n223 GND.n222 5.27
R3150 GND.n191 GND.n190 5.27
R3151 GND.n183 GND.n182 5.27
R3152 GND.n149 GND.n148 5.27
R3153 GND.n142 GND.n141 5.27
R3154 GND.n110 GND.n109 5.27
R3155 GND.n102 GND.n101 5.27
R3156 GND.n565 GND.n564 5.27
R3157 GND.n558 GND.n557 5.27
R3158 GND.n526 GND.n525 5.27
R3159 GND.n518 GND.n517 5.27
R3160 GND.n484 GND.n483 5.27
R3161 GND.n477 GND.n476 5.27
R3162 GND.n445 GND.n444 5.27
R3163 GND.n437 GND.n436 5.27
R3164 GND.n403 GND.n402 5.27
R3165 GND.n396 GND.n395 5.27
R3166 GND.n364 GND.n363 5.27
R3167 GND.n356 GND.n355 5.27
R3168 GND.n322 GND.n321 5.27
R3169 GND.n315 GND.n314 5.27
R3170 GND.n283 GND.n282 5.27
R3171 GND.n275 GND.n274 5.27
R3172 GND.n1226 GND.n1225 5.27
R3173 GND.n1219 GND.n1218 5.27
R3174 GND.n1187 GND.n1186 5.27
R3175 GND.n1179 GND.n1178 5.27
R3176 GND.n1145 GND.n1144 5.27
R3177 GND.n1138 GND.n1137 5.27
R3178 GND.n1106 GND.n1105 5.27
R3179 GND.n1098 GND.n1097 5.27
R3180 GND.n1064 GND.n1063 5.27
R3181 GND.n1057 GND.n1056 5.27
R3182 GND.n1025 GND.n1024 5.27
R3183 GND.n1017 GND.n1016 5.27
R3184 GND.n983 GND.n982 5.27
R3185 GND.n976 GND.n975 5.27
R3186 GND.n944 GND.n943 5.27
R3187 GND.n936 GND.n935 5.27
R3188 GND.n902 GND.n901 5.27
R3189 GND.n895 GND.n894 5.27
R3190 GND.n863 GND.n862 5.27
R3191 GND.n855 GND.n854 5.27
R3192 GND.n821 GND.n820 5.27
R3193 GND.n814 GND.n813 5.27
R3194 GND.n782 GND.n781 5.27
R3195 GND.n774 GND.n773 5.27
R3196 GND.n740 GND.n739 5.27
R3197 GND.n733 GND.n732 5.27
R3198 GND.n701 GND.n700 5.27
R3199 GND.n693 GND.n692 5.27
R3200 GND.n659 GND.n658 5.27
R3201 GND.n652 GND.n651 5.27
R3202 GND.n620 GND.n619 5.27
R3203 GND.n612 GND.n611 5.27
R3204 GND.n1881 GND.n1880 5.27
R3205 GND.n1874 GND.n1873 5.27
R3206 GND.n1842 GND.n1841 5.27
R3207 GND.n1834 GND.n1833 5.27
R3208 GND.n1800 GND.n1799 5.27
R3209 GND.n1793 GND.n1792 5.27
R3210 GND.n1761 GND.n1760 5.27
R3211 GND.n1753 GND.n1752 5.27
R3212 GND.n1719 GND.n1718 5.27
R3213 GND.n1712 GND.n1711 5.27
R3214 GND.n1680 GND.n1679 5.27
R3215 GND.n1672 GND.n1671 5.27
R3216 GND.n1638 GND.n1637 5.27
R3217 GND.n1631 GND.n1630 5.27
R3218 GND.n1599 GND.n1598 5.27
R3219 GND.n1591 GND.n1590 5.27
R3220 GND.n1557 GND.n1556 5.27
R3221 GND.n1550 GND.n1549 5.27
R3222 GND.n1518 GND.n1517 5.27
R3223 GND.n1510 GND.n1509 5.27
R3224 GND.n1476 GND.n1475 5.27
R3225 GND.n1469 GND.n1468 5.27
R3226 GND.n1437 GND.n1436 5.27
R3227 GND.n1429 GND.n1428 5.27
R3228 GND.n1395 GND.n1394 5.27
R3229 GND.n1388 GND.n1387 5.27
R3230 GND.n1356 GND.n1355 5.27
R3231 GND.n1348 GND.n1347 5.27
R3232 GND.n1314 GND.n1313 5.27
R3233 GND.n1307 GND.n1306 5.27
R3234 GND.n1275 GND.n1274 5.27
R3235 GND.n1267 GND.n1266 5.27
R3236 GND.n2546 GND.n2545 5.27
R3237 GND.n2539 GND.n2538 5.27
R3238 GND.n2507 GND.n2506 5.27
R3239 GND.n2499 GND.n2498 5.27
R3240 GND.n2465 GND.n2464 5.27
R3241 GND.n2458 GND.n2457 5.27
R3242 GND.n2426 GND.n2425 5.27
R3243 GND.n2418 GND.n2417 5.27
R3244 GND.n2384 GND.n2383 5.27
R3245 GND.n2377 GND.n2376 5.27
R3246 GND.n2345 GND.n2344 5.27
R3247 GND.n2337 GND.n2336 5.27
R3248 GND.n2303 GND.n2302 5.27
R3249 GND.n2296 GND.n2295 5.27
R3250 GND.n2264 GND.n2263 5.27
R3251 GND.n2256 GND.n2255 5.27
R3252 GND.n2222 GND.n2221 5.27
R3253 GND.n2215 GND.n2214 5.27
R3254 GND.n2183 GND.n2182 5.27
R3255 GND.n2175 GND.n2174 5.27
R3256 GND.n2141 GND.n2140 5.27
R3257 GND.n2134 GND.n2133 5.27
R3258 GND.n2102 GND.n2101 5.27
R3259 GND.n2094 GND.n2093 5.27
R3260 GND.n2060 GND.n2059 5.27
R3261 GND.n2053 GND.n2052 5.27
R3262 GND.n2021 GND.n2020 5.27
R3263 GND.n2013 GND.n2012 5.27
R3264 GND.n1979 GND.n1978 5.27
R3265 GND.n1972 GND.n1971 5.27
R3266 GND.n1940 GND.n1939 5.27
R3267 GND.n1932 GND.n1931 5.27
R3268 GND.n3201 GND.n3200 5.27
R3269 GND.n3194 GND.n3193 5.27
R3270 GND.n3162 GND.n3161 5.27
R3271 GND.n3154 GND.n3153 5.27
R3272 GND.n3120 GND.n3119 5.27
R3273 GND.n3113 GND.n3112 5.27
R3274 GND.n3081 GND.n3080 5.27
R3275 GND.n3073 GND.n3072 5.27
R3276 GND.n3039 GND.n3038 5.27
R3277 GND.n3032 GND.n3031 5.27
R3278 GND.n3000 GND.n2999 5.27
R3279 GND.n2992 GND.n2991 5.27
R3280 GND.n2958 GND.n2957 5.27
R3281 GND.n2951 GND.n2950 5.27
R3282 GND.n2919 GND.n2918 5.27
R3283 GND.n2911 GND.n2910 5.27
R3284 GND.n2877 GND.n2876 5.27
R3285 GND.n2870 GND.n2869 5.27
R3286 GND.n2838 GND.n2837 5.27
R3287 GND.n2830 GND.n2829 5.27
R3288 GND.n2796 GND.n2795 5.27
R3289 GND.n2789 GND.n2788 5.27
R3290 GND.n2757 GND.n2756 5.27
R3291 GND.n2749 GND.n2748 5.27
R3292 GND.n2715 GND.n2714 5.27
R3293 GND.n2708 GND.n2707 5.27
R3294 GND.n2676 GND.n2675 5.27
R3295 GND.n2668 GND.n2667 5.27
R3296 GND.n2634 GND.n2633 5.27
R3297 GND.n2627 GND.n2626 5.27
R3298 GND.n2595 GND.n2594 5.27
R3299 GND.n2587 GND.n2586 5.27
R3300 GND.n3856 GND.n3855 5.27
R3301 GND.n3849 GND.n3848 5.27
R3302 GND.n3817 GND.n3816 5.27
R3303 GND.n3809 GND.n3808 5.27
R3304 GND.n3775 GND.n3774 5.27
R3305 GND.n3768 GND.n3767 5.27
R3306 GND.n3736 GND.n3735 5.27
R3307 GND.n3728 GND.n3727 5.27
R3308 GND.n3694 GND.n3693 5.27
R3309 GND.n3687 GND.n3686 5.27
R3310 GND.n3655 GND.n3654 5.27
R3311 GND.n3647 GND.n3646 5.27
R3312 GND.n3613 GND.n3612 5.27
R3313 GND.n3606 GND.n3605 5.27
R3314 GND.n3574 GND.n3573 5.27
R3315 GND.n3566 GND.n3565 5.27
R3316 GND.n3532 GND.n3531 5.27
R3317 GND.n3525 GND.n3524 5.27
R3318 GND.n3493 GND.n3492 5.27
R3319 GND.n3485 GND.n3484 5.27
R3320 GND.n3451 GND.n3450 5.27
R3321 GND.n3444 GND.n3443 5.27
R3322 GND.n3412 GND.n3411 5.27
R3323 GND.n3404 GND.n3403 5.27
R3324 GND.n3370 GND.n3369 5.27
R3325 GND.n3363 GND.n3362 5.27
R3326 GND.n3331 GND.n3330 5.27
R3327 GND.n3323 GND.n3322 5.27
R3328 GND.n3289 GND.n3288 5.27
R3329 GND.n3282 GND.n3281 5.27
R3330 GND.n3250 GND.n3249 5.27
R3331 GND.n3242 GND.n3241 5.27
R3332 GND.n4511 GND.n4510 5.27
R3333 GND.n4504 GND.n4503 5.27
R3334 GND.n4472 GND.n4471 5.27
R3335 GND.n4464 GND.n4463 5.27
R3336 GND.n4430 GND.n4429 5.27
R3337 GND.n4423 GND.n4422 5.27
R3338 GND.n4391 GND.n4390 5.27
R3339 GND.n4383 GND.n4382 5.27
R3340 GND.n4349 GND.n4348 5.27
R3341 GND.n4342 GND.n4341 5.27
R3342 GND.n4310 GND.n4309 5.27
R3343 GND.n4302 GND.n4301 5.27
R3344 GND.n4268 GND.n4267 5.27
R3345 GND.n4261 GND.n4260 5.27
R3346 GND.n4229 GND.n4228 5.27
R3347 GND.n4221 GND.n4220 5.27
R3348 GND.n4187 GND.n4186 5.27
R3349 GND.n4180 GND.n4179 5.27
R3350 GND.n4148 GND.n4147 5.27
R3351 GND.n4140 GND.n4139 5.27
R3352 GND.n4106 GND.n4105 5.27
R3353 GND.n4099 GND.n4098 5.27
R3354 GND.n4067 GND.n4066 5.27
R3355 GND.n4059 GND.n4058 5.27
R3356 GND.n4025 GND.n4024 5.27
R3357 GND.n4018 GND.n4017 5.27
R3358 GND.n3986 GND.n3985 5.27
R3359 GND.n3978 GND.n3977 5.27
R3360 GND.n3944 GND.n3943 5.27
R3361 GND.n3937 GND.n3936 5.27
R3362 GND.n3905 GND.n3904 5.27
R3363 GND.n3897 GND.n3896 5.27
R3364 GND.n5176 GND.n5175 5.27
R3365 GND.n5169 GND.n5168 5.27
R3366 GND.n5137 GND.n5136 5.27
R3367 GND.n5129 GND.n5128 5.27
R3368 GND.n5095 GND.n5094 5.27
R3369 GND.n5088 GND.n5087 5.27
R3370 GND.n5056 GND.n5055 5.27
R3371 GND.n5048 GND.n5047 5.27
R3372 GND.n5014 GND.n5013 5.27
R3373 GND.n5007 GND.n5006 5.27
R3374 GND.n4975 GND.n4974 5.27
R3375 GND.n4967 GND.n4966 5.27
R3376 GND.n4933 GND.n4932 5.27
R3377 GND.n4926 GND.n4925 5.27
R3378 GND.n4894 GND.n4893 5.27
R3379 GND.n4886 GND.n4885 5.27
R3380 GND.n4852 GND.n4851 5.27
R3381 GND.n4845 GND.n4844 5.27
R3382 GND.n4813 GND.n4812 5.27
R3383 GND.n4805 GND.n4804 5.27
R3384 GND.n4771 GND.n4770 5.27
R3385 GND.n4764 GND.n4763 5.27
R3386 GND.n4732 GND.n4731 5.27
R3387 GND.n4724 GND.n4723 5.27
R3388 GND.n4690 GND.n4689 5.27
R3389 GND.n4683 GND.n4682 5.27
R3390 GND.n4651 GND.n4650 5.27
R3391 GND.n4643 GND.n4642 5.27
R3392 GND.n4609 GND.n4608 5.27
R3393 GND.n4602 GND.n4601 5.27
R3394 GND.n4570 GND.n4569 5.27
R3395 GND.n4562 GND.n4561 5.27
R3396 GND.n65 GND.n63 4.048
R3397 GND.n25 GND.n23 4.048
R3398 GND.n197 GND.n195 4.048
R3399 GND.n116 GND.n114 4.048
R3400 GND.n532 GND.n530 4.048
R3401 GND.n451 GND.n449 4.048
R3402 GND.n370 GND.n368 4.048
R3403 GND.n289 GND.n287 4.048
R3404 GND.n1193 GND.n1191 4.048
R3405 GND.n1112 GND.n1110 4.048
R3406 GND.n1031 GND.n1029 4.048
R3407 GND.n950 GND.n948 4.048
R3408 GND.n869 GND.n867 4.048
R3409 GND.n788 GND.n786 4.048
R3410 GND.n707 GND.n705 4.048
R3411 GND.n626 GND.n624 4.048
R3412 GND.n1848 GND.n1846 4.048
R3413 GND.n1767 GND.n1765 4.048
R3414 GND.n1686 GND.n1684 4.048
R3415 GND.n1605 GND.n1603 4.048
R3416 GND.n1524 GND.n1522 4.048
R3417 GND.n1443 GND.n1441 4.048
R3418 GND.n1362 GND.n1360 4.048
R3419 GND.n1281 GND.n1279 4.048
R3420 GND.n2513 GND.n2511 4.048
R3421 GND.n2432 GND.n2430 4.048
R3422 GND.n2351 GND.n2349 4.048
R3423 GND.n2270 GND.n2268 4.048
R3424 GND.n2189 GND.n2187 4.048
R3425 GND.n2108 GND.n2106 4.048
R3426 GND.n2027 GND.n2025 4.048
R3427 GND.n1946 GND.n1944 4.048
R3428 GND.n3168 GND.n3166 4.048
R3429 GND.n3087 GND.n3085 4.048
R3430 GND.n3006 GND.n3004 4.048
R3431 GND.n2925 GND.n2923 4.048
R3432 GND.n2844 GND.n2842 4.048
R3433 GND.n2763 GND.n2761 4.048
R3434 GND.n2682 GND.n2680 4.048
R3435 GND.n2601 GND.n2599 4.048
R3436 GND.n3823 GND.n3821 4.048
R3437 GND.n3742 GND.n3740 4.048
R3438 GND.n3661 GND.n3659 4.048
R3439 GND.n3580 GND.n3578 4.048
R3440 GND.n3499 GND.n3497 4.048
R3441 GND.n3418 GND.n3416 4.048
R3442 GND.n3337 GND.n3335 4.048
R3443 GND.n3256 GND.n3254 4.048
R3444 GND.n4478 GND.n4476 4.048
R3445 GND.n4397 GND.n4395 4.048
R3446 GND.n4316 GND.n4314 4.048
R3447 GND.n4235 GND.n4233 4.048
R3448 GND.n4154 GND.n4152 4.048
R3449 GND.n4073 GND.n4071 4.048
R3450 GND.n3992 GND.n3990 4.048
R3451 GND.n3911 GND.n3909 4.048
R3452 GND.n5143 GND.n5141 4.048
R3453 GND.n5062 GND.n5060 4.048
R3454 GND.n4981 GND.n4979 4.048
R3455 GND.n4900 GND.n4898 4.048
R3456 GND.n4819 GND.n4817 4.048
R3457 GND.n4738 GND.n4736 4.048
R3458 GND.n4657 GND.n4655 4.048
R3459 GND.n4576 GND.n4574 4.048
R3460 GND.n237 GND.n235 4.047
R3461 GND.n156 GND.n154 4.047
R3462 GND.n572 GND.n570 4.047
R3463 GND.n491 GND.n489 4.047
R3464 GND.n410 GND.n408 4.047
R3465 GND.n329 GND.n327 4.047
R3466 GND.n1233 GND.n1231 4.047
R3467 GND.n1152 GND.n1150 4.047
R3468 GND.n1071 GND.n1069 4.047
R3469 GND.n990 GND.n988 4.047
R3470 GND.n909 GND.n907 4.047
R3471 GND.n828 GND.n826 4.047
R3472 GND.n747 GND.n745 4.047
R3473 GND.n666 GND.n664 4.047
R3474 GND.n1888 GND.n1886 4.047
R3475 GND.n1807 GND.n1805 4.047
R3476 GND.n1726 GND.n1724 4.047
R3477 GND.n1645 GND.n1643 4.047
R3478 GND.n1564 GND.n1562 4.047
R3479 GND.n1483 GND.n1481 4.047
R3480 GND.n1402 GND.n1400 4.047
R3481 GND.n1321 GND.n1319 4.047
R3482 GND.n2553 GND.n2551 4.047
R3483 GND.n2472 GND.n2470 4.047
R3484 GND.n2391 GND.n2389 4.047
R3485 GND.n2310 GND.n2308 4.047
R3486 GND.n2229 GND.n2227 4.047
R3487 GND.n2148 GND.n2146 4.047
R3488 GND.n2067 GND.n2065 4.047
R3489 GND.n1986 GND.n1984 4.047
R3490 GND.n3208 GND.n3206 4.047
R3491 GND.n3127 GND.n3125 4.047
R3492 GND.n3046 GND.n3044 4.047
R3493 GND.n2965 GND.n2963 4.047
R3494 GND.n2884 GND.n2882 4.047
R3495 GND.n2803 GND.n2801 4.047
R3496 GND.n2722 GND.n2720 4.047
R3497 GND.n2641 GND.n2639 4.047
R3498 GND.n3863 GND.n3861 4.047
R3499 GND.n3782 GND.n3780 4.047
R3500 GND.n3701 GND.n3699 4.047
R3501 GND.n3620 GND.n3618 4.047
R3502 GND.n3539 GND.n3537 4.047
R3503 GND.n3458 GND.n3456 4.047
R3504 GND.n3377 GND.n3375 4.047
R3505 GND.n3296 GND.n3294 4.047
R3506 GND.n4518 GND.n4516 4.047
R3507 GND.n4437 GND.n4435 4.047
R3508 GND.n4356 GND.n4354 4.047
R3509 GND.n4275 GND.n4273 4.047
R3510 GND.n4194 GND.n4192 4.047
R3511 GND.n4113 GND.n4111 4.047
R3512 GND.n4032 GND.n4030 4.047
R3513 GND.n3951 GND.n3949 4.047
R3514 GND.n5183 GND.n5181 4.047
R3515 GND.n5102 GND.n5100 4.047
R3516 GND.n5021 GND.n5019 4.047
R3517 GND.n4940 GND.n4938 4.047
R3518 GND.n4859 GND.n4857 4.047
R3519 GND.n4778 GND.n4776 4.047
R3520 GND.n4697 GND.n4695 4.047
R3521 GND.n4616 GND.n4614 4.047
R3522 GND.n89 GND.n57 3.924
R3523 GND.n49 GND.n17 3.924
R3524 GND.n261 GND.n228 3.924
R3525 GND.n221 GND.n189 3.924
R3526 GND.n180 GND.n147 3.924
R3527 GND.n140 GND.n108 3.924
R3528 GND.n596 GND.n563 3.924
R3529 GND.n556 GND.n524 3.924
R3530 GND.n515 GND.n482 3.924
R3531 GND.n475 GND.n443 3.924
R3532 GND.n434 GND.n401 3.924
R3533 GND.n394 GND.n362 3.924
R3534 GND.n353 GND.n320 3.924
R3535 GND.n313 GND.n281 3.924
R3536 GND.n1257 GND.n1224 3.924
R3537 GND.n1217 GND.n1185 3.924
R3538 GND.n1176 GND.n1143 3.924
R3539 GND.n1136 GND.n1104 3.924
R3540 GND.n1095 GND.n1062 3.924
R3541 GND.n1055 GND.n1023 3.924
R3542 GND.n1014 GND.n981 3.924
R3543 GND.n974 GND.n942 3.924
R3544 GND.n933 GND.n900 3.924
R3545 GND.n893 GND.n861 3.924
R3546 GND.n852 GND.n819 3.924
R3547 GND.n812 GND.n780 3.924
R3548 GND.n771 GND.n738 3.924
R3549 GND.n731 GND.n699 3.924
R3550 GND.n690 GND.n657 3.924
R3551 GND.n650 GND.n618 3.924
R3552 GND.n1912 GND.n1879 3.924
R3553 GND.n1872 GND.n1840 3.924
R3554 GND.n1831 GND.n1798 3.924
R3555 GND.n1791 GND.n1759 3.924
R3556 GND.n1750 GND.n1717 3.924
R3557 GND.n1710 GND.n1678 3.924
R3558 GND.n1669 GND.n1636 3.924
R3559 GND.n1629 GND.n1597 3.924
R3560 GND.n1588 GND.n1555 3.924
R3561 GND.n1548 GND.n1516 3.924
R3562 GND.n1507 GND.n1474 3.924
R3563 GND.n1467 GND.n1435 3.924
R3564 GND.n1426 GND.n1393 3.924
R3565 GND.n1386 GND.n1354 3.924
R3566 GND.n1345 GND.n1312 3.924
R3567 GND.n1305 GND.n1273 3.924
R3568 GND.n2577 GND.n2544 3.924
R3569 GND.n2537 GND.n2505 3.924
R3570 GND.n2496 GND.n2463 3.924
R3571 GND.n2456 GND.n2424 3.924
R3572 GND.n2415 GND.n2382 3.924
R3573 GND.n2375 GND.n2343 3.924
R3574 GND.n2334 GND.n2301 3.924
R3575 GND.n2294 GND.n2262 3.924
R3576 GND.n2253 GND.n2220 3.924
R3577 GND.n2213 GND.n2181 3.924
R3578 GND.n2172 GND.n2139 3.924
R3579 GND.n2132 GND.n2100 3.924
R3580 GND.n2091 GND.n2058 3.924
R3581 GND.n2051 GND.n2019 3.924
R3582 GND.n2010 GND.n1977 3.924
R3583 GND.n1970 GND.n1938 3.924
R3584 GND.n3232 GND.n3199 3.924
R3585 GND.n3192 GND.n3160 3.924
R3586 GND.n3151 GND.n3118 3.924
R3587 GND.n3111 GND.n3079 3.924
R3588 GND.n3070 GND.n3037 3.924
R3589 GND.n3030 GND.n2998 3.924
R3590 GND.n2989 GND.n2956 3.924
R3591 GND.n2949 GND.n2917 3.924
R3592 GND.n2908 GND.n2875 3.924
R3593 GND.n2868 GND.n2836 3.924
R3594 GND.n2827 GND.n2794 3.924
R3595 GND.n2787 GND.n2755 3.924
R3596 GND.n2746 GND.n2713 3.924
R3597 GND.n2706 GND.n2674 3.924
R3598 GND.n2665 GND.n2632 3.924
R3599 GND.n2625 GND.n2593 3.924
R3600 GND.n3887 GND.n3854 3.924
R3601 GND.n3847 GND.n3815 3.924
R3602 GND.n3806 GND.n3773 3.924
R3603 GND.n3766 GND.n3734 3.924
R3604 GND.n3725 GND.n3692 3.924
R3605 GND.n3685 GND.n3653 3.924
R3606 GND.n3644 GND.n3611 3.924
R3607 GND.n3604 GND.n3572 3.924
R3608 GND.n3563 GND.n3530 3.924
R3609 GND.n3523 GND.n3491 3.924
R3610 GND.n3482 GND.n3449 3.924
R3611 GND.n3442 GND.n3410 3.924
R3612 GND.n3401 GND.n3368 3.924
R3613 GND.n3361 GND.n3329 3.924
R3614 GND.n3320 GND.n3287 3.924
R3615 GND.n3280 GND.n3248 3.924
R3616 GND.n4542 GND.n4509 3.924
R3617 GND.n4502 GND.n4470 3.924
R3618 GND.n4461 GND.n4428 3.924
R3619 GND.n4421 GND.n4389 3.924
R3620 GND.n4380 GND.n4347 3.924
R3621 GND.n4340 GND.n4308 3.924
R3622 GND.n4299 GND.n4266 3.924
R3623 GND.n4259 GND.n4227 3.924
R3624 GND.n4218 GND.n4185 3.924
R3625 GND.n4178 GND.n4146 3.924
R3626 GND.n4137 GND.n4104 3.924
R3627 GND.n4097 GND.n4065 3.924
R3628 GND.n4056 GND.n4023 3.924
R3629 GND.n4016 GND.n3984 3.924
R3630 GND.n3975 GND.n3942 3.924
R3631 GND.n3935 GND.n3903 3.924
R3632 GND.n5207 GND.n5174 3.924
R3633 GND.n5167 GND.n5135 3.924
R3634 GND.n5126 GND.n5093 3.924
R3635 GND.n5086 GND.n5054 3.924
R3636 GND.n5045 GND.n5012 3.924
R3637 GND.n5005 GND.n4973 3.924
R3638 GND.n4964 GND.n4931 3.924
R3639 GND.n4924 GND.n4892 3.924
R3640 GND.n4883 GND.n4850 3.924
R3641 GND.n4843 GND.n4811 3.924
R3642 GND.n4802 GND.n4769 3.924
R3643 GND.n4762 GND.n4730 3.924
R3644 GND.n4721 GND.n4688 3.924
R3645 GND.n4681 GND.n4649 3.924
R3646 GND.n4640 GND.n4607 3.924
R3647 GND.n4600 GND.n4568 3.924
R3648 GND.n254 GND.n252 3.396
R3649 GND.n173 GND.n171 3.396
R3650 GND.n589 GND.n587 3.396
R3651 GND.n508 GND.n506 3.396
R3652 GND.n427 GND.n425 3.396
R3653 GND.n346 GND.n344 3.396
R3654 GND.n1250 GND.n1248 3.396
R3655 GND.n1169 GND.n1167 3.396
R3656 GND.n1088 GND.n1086 3.396
R3657 GND.n1007 GND.n1005 3.396
R3658 GND.n926 GND.n924 3.396
R3659 GND.n845 GND.n843 3.396
R3660 GND.n764 GND.n762 3.396
R3661 GND.n683 GND.n681 3.396
R3662 GND.n1905 GND.n1903 3.396
R3663 GND.n1824 GND.n1822 3.396
R3664 GND.n1743 GND.n1741 3.396
R3665 GND.n1662 GND.n1660 3.396
R3666 GND.n1581 GND.n1579 3.396
R3667 GND.n1500 GND.n1498 3.396
R3668 GND.n1419 GND.n1417 3.396
R3669 GND.n1338 GND.n1336 3.396
R3670 GND.n2570 GND.n2568 3.396
R3671 GND.n2489 GND.n2487 3.396
R3672 GND.n2408 GND.n2406 3.396
R3673 GND.n2327 GND.n2325 3.396
R3674 GND.n2246 GND.n2244 3.396
R3675 GND.n2165 GND.n2163 3.396
R3676 GND.n2084 GND.n2082 3.396
R3677 GND.n2003 GND.n2001 3.396
R3678 GND.n3225 GND.n3223 3.396
R3679 GND.n3144 GND.n3142 3.396
R3680 GND.n3063 GND.n3061 3.396
R3681 GND.n2982 GND.n2980 3.396
R3682 GND.n2901 GND.n2899 3.396
R3683 GND.n2820 GND.n2818 3.396
R3684 GND.n2739 GND.n2737 3.396
R3685 GND.n2658 GND.n2656 3.396
R3686 GND.n3880 GND.n3878 3.396
R3687 GND.n3799 GND.n3797 3.396
R3688 GND.n3718 GND.n3716 3.396
R3689 GND.n3637 GND.n3635 3.396
R3690 GND.n3556 GND.n3554 3.396
R3691 GND.n3475 GND.n3473 3.396
R3692 GND.n3394 GND.n3392 3.396
R3693 GND.n3313 GND.n3311 3.396
R3694 GND.n4535 GND.n4533 3.396
R3695 GND.n4454 GND.n4452 3.396
R3696 GND.n4373 GND.n4371 3.396
R3697 GND.n4292 GND.n4290 3.396
R3698 GND.n4211 GND.n4209 3.396
R3699 GND.n4130 GND.n4128 3.396
R3700 GND.n4049 GND.n4047 3.396
R3701 GND.n3968 GND.n3966 3.396
R3702 GND.n5200 GND.n5198 3.396
R3703 GND.n5119 GND.n5117 3.396
R3704 GND.n5038 GND.n5036 3.396
R3705 GND.n4957 GND.n4955 3.396
R3706 GND.n4876 GND.n4874 3.396
R3707 GND.n4795 GND.n4793 3.396
R3708 GND.n4714 GND.n4712 3.396
R3709 GND.n4633 GND.n4631 3.396
R3710 GND.n81 GND.n80 3.324
R3711 GND.n72 GND.n71 3.324
R3712 GND.n41 GND.n40 3.324
R3713 GND.n32 GND.n31 3.324
R3714 GND.n244 GND.n243 3.324
R3715 GND.n213 GND.n212 3.324
R3716 GND.n204 GND.n203 3.324
R3717 GND.n163 GND.n162 3.324
R3718 GND.n132 GND.n131 3.324
R3719 GND.n123 GND.n122 3.324
R3720 GND.n579 GND.n578 3.324
R3721 GND.n548 GND.n547 3.324
R3722 GND.n539 GND.n538 3.324
R3723 GND.n498 GND.n497 3.324
R3724 GND.n467 GND.n466 3.324
R3725 GND.n458 GND.n457 3.324
R3726 GND.n417 GND.n416 3.324
R3727 GND.n386 GND.n385 3.324
R3728 GND.n377 GND.n376 3.324
R3729 GND.n336 GND.n335 3.324
R3730 GND.n305 GND.n304 3.324
R3731 GND.n296 GND.n295 3.324
R3732 GND.n1240 GND.n1239 3.324
R3733 GND.n1209 GND.n1208 3.324
R3734 GND.n1200 GND.n1199 3.324
R3735 GND.n1159 GND.n1158 3.324
R3736 GND.n1128 GND.n1127 3.324
R3737 GND.n1119 GND.n1118 3.324
R3738 GND.n1078 GND.n1077 3.324
R3739 GND.n1047 GND.n1046 3.324
R3740 GND.n1038 GND.n1037 3.324
R3741 GND.n997 GND.n996 3.324
R3742 GND.n966 GND.n965 3.324
R3743 GND.n957 GND.n956 3.324
R3744 GND.n916 GND.n915 3.324
R3745 GND.n885 GND.n884 3.324
R3746 GND.n876 GND.n875 3.324
R3747 GND.n835 GND.n834 3.324
R3748 GND.n804 GND.n803 3.324
R3749 GND.n795 GND.n794 3.324
R3750 GND.n754 GND.n753 3.324
R3751 GND.n723 GND.n722 3.324
R3752 GND.n714 GND.n713 3.324
R3753 GND.n673 GND.n672 3.324
R3754 GND.n642 GND.n641 3.324
R3755 GND.n633 GND.n632 3.324
R3756 GND.n1895 GND.n1894 3.324
R3757 GND.n1864 GND.n1863 3.324
R3758 GND.n1855 GND.n1854 3.324
R3759 GND.n1814 GND.n1813 3.324
R3760 GND.n1783 GND.n1782 3.324
R3761 GND.n1774 GND.n1773 3.324
R3762 GND.n1733 GND.n1732 3.324
R3763 GND.n1702 GND.n1701 3.324
R3764 GND.n1693 GND.n1692 3.324
R3765 GND.n1652 GND.n1651 3.324
R3766 GND.n1621 GND.n1620 3.324
R3767 GND.n1612 GND.n1611 3.324
R3768 GND.n1571 GND.n1570 3.324
R3769 GND.n1540 GND.n1539 3.324
R3770 GND.n1531 GND.n1530 3.324
R3771 GND.n1490 GND.n1489 3.324
R3772 GND.n1459 GND.n1458 3.324
R3773 GND.n1450 GND.n1449 3.324
R3774 GND.n1409 GND.n1408 3.324
R3775 GND.n1378 GND.n1377 3.324
R3776 GND.n1369 GND.n1368 3.324
R3777 GND.n1328 GND.n1327 3.324
R3778 GND.n1297 GND.n1296 3.324
R3779 GND.n1288 GND.n1287 3.324
R3780 GND.n2560 GND.n2559 3.324
R3781 GND.n2529 GND.n2528 3.324
R3782 GND.n2520 GND.n2519 3.324
R3783 GND.n2479 GND.n2478 3.324
R3784 GND.n2448 GND.n2447 3.324
R3785 GND.n2439 GND.n2438 3.324
R3786 GND.n2398 GND.n2397 3.324
R3787 GND.n2367 GND.n2366 3.324
R3788 GND.n2358 GND.n2357 3.324
R3789 GND.n2317 GND.n2316 3.324
R3790 GND.n2286 GND.n2285 3.324
R3791 GND.n2277 GND.n2276 3.324
R3792 GND.n2236 GND.n2235 3.324
R3793 GND.n2205 GND.n2204 3.324
R3794 GND.n2196 GND.n2195 3.324
R3795 GND.n2155 GND.n2154 3.324
R3796 GND.n2124 GND.n2123 3.324
R3797 GND.n2115 GND.n2114 3.324
R3798 GND.n2074 GND.n2073 3.324
R3799 GND.n2043 GND.n2042 3.324
R3800 GND.n2034 GND.n2033 3.324
R3801 GND.n1993 GND.n1992 3.324
R3802 GND.n1962 GND.n1961 3.324
R3803 GND.n1953 GND.n1952 3.324
R3804 GND.n3215 GND.n3214 3.324
R3805 GND.n3184 GND.n3183 3.324
R3806 GND.n3175 GND.n3174 3.324
R3807 GND.n3134 GND.n3133 3.324
R3808 GND.n3103 GND.n3102 3.324
R3809 GND.n3094 GND.n3093 3.324
R3810 GND.n3053 GND.n3052 3.324
R3811 GND.n3022 GND.n3021 3.324
R3812 GND.n3013 GND.n3012 3.324
R3813 GND.n2972 GND.n2971 3.324
R3814 GND.n2941 GND.n2940 3.324
R3815 GND.n2932 GND.n2931 3.324
R3816 GND.n2891 GND.n2890 3.324
R3817 GND.n2860 GND.n2859 3.324
R3818 GND.n2851 GND.n2850 3.324
R3819 GND.n2810 GND.n2809 3.324
R3820 GND.n2779 GND.n2778 3.324
R3821 GND.n2770 GND.n2769 3.324
R3822 GND.n2729 GND.n2728 3.324
R3823 GND.n2698 GND.n2697 3.324
R3824 GND.n2689 GND.n2688 3.324
R3825 GND.n2648 GND.n2647 3.324
R3826 GND.n2617 GND.n2616 3.324
R3827 GND.n2608 GND.n2607 3.324
R3828 GND.n3870 GND.n3869 3.324
R3829 GND.n3839 GND.n3838 3.324
R3830 GND.n3830 GND.n3829 3.324
R3831 GND.n3789 GND.n3788 3.324
R3832 GND.n3758 GND.n3757 3.324
R3833 GND.n3749 GND.n3748 3.324
R3834 GND.n3708 GND.n3707 3.324
R3835 GND.n3677 GND.n3676 3.324
R3836 GND.n3668 GND.n3667 3.324
R3837 GND.n3627 GND.n3626 3.324
R3838 GND.n3596 GND.n3595 3.324
R3839 GND.n3587 GND.n3586 3.324
R3840 GND.n3546 GND.n3545 3.324
R3841 GND.n3515 GND.n3514 3.324
R3842 GND.n3506 GND.n3505 3.324
R3843 GND.n3465 GND.n3464 3.324
R3844 GND.n3434 GND.n3433 3.324
R3845 GND.n3425 GND.n3424 3.324
R3846 GND.n3384 GND.n3383 3.324
R3847 GND.n3353 GND.n3352 3.324
R3848 GND.n3344 GND.n3343 3.324
R3849 GND.n3303 GND.n3302 3.324
R3850 GND.n3272 GND.n3271 3.324
R3851 GND.n3263 GND.n3262 3.324
R3852 GND.n4525 GND.n4524 3.324
R3853 GND.n4494 GND.n4493 3.324
R3854 GND.n4485 GND.n4484 3.324
R3855 GND.n4444 GND.n4443 3.324
R3856 GND.n4413 GND.n4412 3.324
R3857 GND.n4404 GND.n4403 3.324
R3858 GND.n4363 GND.n4362 3.324
R3859 GND.n4332 GND.n4331 3.324
R3860 GND.n4323 GND.n4322 3.324
R3861 GND.n4282 GND.n4281 3.324
R3862 GND.n4251 GND.n4250 3.324
R3863 GND.n4242 GND.n4241 3.324
R3864 GND.n4201 GND.n4200 3.324
R3865 GND.n4170 GND.n4169 3.324
R3866 GND.n4161 GND.n4160 3.324
R3867 GND.n4120 GND.n4119 3.324
R3868 GND.n4089 GND.n4088 3.324
R3869 GND.n4080 GND.n4079 3.324
R3870 GND.n4039 GND.n4038 3.324
R3871 GND.n4008 GND.n4007 3.324
R3872 GND.n3999 GND.n3998 3.324
R3873 GND.n3958 GND.n3957 3.324
R3874 GND.n3927 GND.n3926 3.324
R3875 GND.n3918 GND.n3917 3.324
R3876 GND.n5190 GND.n5189 3.324
R3877 GND.n5159 GND.n5158 3.324
R3878 GND.n5150 GND.n5149 3.324
R3879 GND.n5109 GND.n5108 3.324
R3880 GND.n5078 GND.n5077 3.324
R3881 GND.n5069 GND.n5068 3.324
R3882 GND.n5028 GND.n5027 3.324
R3883 GND.n4997 GND.n4996 3.324
R3884 GND.n4988 GND.n4987 3.324
R3885 GND.n4947 GND.n4946 3.324
R3886 GND.n4916 GND.n4915 3.324
R3887 GND.n4907 GND.n4906 3.324
R3888 GND.n4866 GND.n4865 3.324
R3889 GND.n4835 GND.n4834 3.324
R3890 GND.n4826 GND.n4825 3.324
R3891 GND.n4785 GND.n4784 3.324
R3892 GND.n4754 GND.n4753 3.324
R3893 GND.n4745 GND.n4744 3.324
R3894 GND.n4704 GND.n4703 3.324
R3895 GND.n4673 GND.n4672 3.324
R3896 GND.n4664 GND.n4663 3.324
R3897 GND.n4623 GND.n4622 3.324
R3898 GND.n4592 GND.n4591 3.324
R3899 GND.n4583 GND.n4582 3.324
R3900 GND.n3 GND.n2 2.461
R3901 GND.n94 GND.n93 2.461
R3902 GND.n267 GND.n266 2.461
R3903 GND.n604 GND.n603 2.461
R3904 GND.n1924 GND.n1923 2.461
R3905 GND.n4554 GND.n4553 2.461
R3906 GND.n5230 GND.n9 2.272
R3907 GND.n5228 GND.n100 2.272
R3908 GND.n5226 GND.n273 2.272
R3909 GND.n5224 GND.n610 2.272
R3910 GND.n5221 GND.n1930 2.272
R3911 GND.n5216 GND.n4560 2.272
R3912 GND.n254 GND.n253 2.163
R3913 GND.n173 GND.n172 2.163
R3914 GND.n589 GND.n588 2.163
R3915 GND.n508 GND.n507 2.163
R3916 GND.n427 GND.n426 2.163
R3917 GND.n346 GND.n345 2.163
R3918 GND.n1250 GND.n1249 2.163
R3919 GND.n1169 GND.n1168 2.163
R3920 GND.n1088 GND.n1087 2.163
R3921 GND.n1007 GND.n1006 2.163
R3922 GND.n926 GND.n925 2.163
R3923 GND.n845 GND.n844 2.163
R3924 GND.n764 GND.n763 2.163
R3925 GND.n683 GND.n682 2.163
R3926 GND.n1905 GND.n1904 2.163
R3927 GND.n1824 GND.n1823 2.163
R3928 GND.n1743 GND.n1742 2.163
R3929 GND.n1662 GND.n1661 2.163
R3930 GND.n1581 GND.n1580 2.163
R3931 GND.n1500 GND.n1499 2.163
R3932 GND.n1419 GND.n1418 2.163
R3933 GND.n1338 GND.n1337 2.163
R3934 GND.n2570 GND.n2569 2.163
R3935 GND.n2489 GND.n2488 2.163
R3936 GND.n2408 GND.n2407 2.163
R3937 GND.n2327 GND.n2326 2.163
R3938 GND.n2246 GND.n2245 2.163
R3939 GND.n2165 GND.n2164 2.163
R3940 GND.n2084 GND.n2083 2.163
R3941 GND.n2003 GND.n2002 2.163
R3942 GND.n3225 GND.n3224 2.163
R3943 GND.n3144 GND.n3143 2.163
R3944 GND.n3063 GND.n3062 2.163
R3945 GND.n2982 GND.n2981 2.163
R3946 GND.n2901 GND.n2900 2.163
R3947 GND.n2820 GND.n2819 2.163
R3948 GND.n2739 GND.n2738 2.163
R3949 GND.n2658 GND.n2657 2.163
R3950 GND.n3880 GND.n3879 2.163
R3951 GND.n3799 GND.n3798 2.163
R3952 GND.n3718 GND.n3717 2.163
R3953 GND.n3637 GND.n3636 2.163
R3954 GND.n3556 GND.n3555 2.163
R3955 GND.n3475 GND.n3474 2.163
R3956 GND.n3394 GND.n3393 2.163
R3957 GND.n3313 GND.n3312 2.163
R3958 GND.n4535 GND.n4534 2.163
R3959 GND.n4454 GND.n4453 2.163
R3960 GND.n4373 GND.n4372 2.163
R3961 GND.n4292 GND.n4291 2.163
R3962 GND.n4211 GND.n4210 2.163
R3963 GND.n4130 GND.n4129 2.163
R3964 GND.n4049 GND.n4048 2.163
R3965 GND.n3968 GND.n3967 2.163
R3966 GND.n5200 GND.n5199 2.163
R3967 GND.n5119 GND.n5118 2.163
R3968 GND.n5038 GND.n5037 2.163
R3969 GND.n4957 GND.n4956 2.163
R3970 GND.n4876 GND.n4875 2.163
R3971 GND.n4795 GND.n4794 2.163
R3972 GND.n4714 GND.n4713 2.163
R3973 GND.n4633 GND.n4632 2.163
R3974 GND.n263 GND.n262 1.378
R3975 GND.n598 GND.n597 1.378
R3976 GND.n1259 GND.n1258 1.378
R3977 GND.n1914 GND.n1913 1.378
R3978 GND.n2579 GND.n2578 1.378
R3979 GND.n3234 GND.n3233 1.378
R3980 GND.n3889 GND.n3888 1.378
R3981 GND.n4544 GND.n4543 1.378
R3982 GND.n5209 GND.n5208 1.378
R3983 GND.n5229 GND.n90 1.206
R3984 GND.n63 GND.n59 1.129
R3985 GND.n57 GND.n51 1.129
R3986 GND.n23 GND.n19 1.129
R3987 GND.n17 GND.n11 1.129
R3988 GND.n235 GND.n230 1.129
R3989 GND.n228 GND.n223 1.129
R3990 GND.n195 GND.n191 1.129
R3991 GND.n189 GND.n183 1.129
R3992 GND.n154 GND.n149 1.129
R3993 GND.n147 GND.n142 1.129
R3994 GND.n114 GND.n110 1.129
R3995 GND.n108 GND.n102 1.129
R3996 GND.n570 GND.n565 1.129
R3997 GND.n563 GND.n558 1.129
R3998 GND.n530 GND.n526 1.129
R3999 GND.n524 GND.n518 1.129
R4000 GND.n489 GND.n484 1.129
R4001 GND.n482 GND.n477 1.129
R4002 GND.n449 GND.n445 1.129
R4003 GND.n443 GND.n437 1.129
R4004 GND.n408 GND.n403 1.129
R4005 GND.n401 GND.n396 1.129
R4006 GND.n368 GND.n364 1.129
R4007 GND.n362 GND.n356 1.129
R4008 GND.n327 GND.n322 1.129
R4009 GND.n320 GND.n315 1.129
R4010 GND.n287 GND.n283 1.129
R4011 GND.n281 GND.n275 1.129
R4012 GND.n1231 GND.n1226 1.129
R4013 GND.n1224 GND.n1219 1.129
R4014 GND.n1191 GND.n1187 1.129
R4015 GND.n1185 GND.n1179 1.129
R4016 GND.n1150 GND.n1145 1.129
R4017 GND.n1143 GND.n1138 1.129
R4018 GND.n1110 GND.n1106 1.129
R4019 GND.n1104 GND.n1098 1.129
R4020 GND.n1069 GND.n1064 1.129
R4021 GND.n1062 GND.n1057 1.129
R4022 GND.n1029 GND.n1025 1.129
R4023 GND.n1023 GND.n1017 1.129
R4024 GND.n988 GND.n983 1.129
R4025 GND.n981 GND.n976 1.129
R4026 GND.n948 GND.n944 1.129
R4027 GND.n942 GND.n936 1.129
R4028 GND.n907 GND.n902 1.129
R4029 GND.n900 GND.n895 1.129
R4030 GND.n867 GND.n863 1.129
R4031 GND.n861 GND.n855 1.129
R4032 GND.n826 GND.n821 1.129
R4033 GND.n819 GND.n814 1.129
R4034 GND.n786 GND.n782 1.129
R4035 GND.n780 GND.n774 1.129
R4036 GND.n745 GND.n740 1.129
R4037 GND.n738 GND.n733 1.129
R4038 GND.n705 GND.n701 1.129
R4039 GND.n699 GND.n693 1.129
R4040 GND.n664 GND.n659 1.129
R4041 GND.n657 GND.n652 1.129
R4042 GND.n624 GND.n620 1.129
R4043 GND.n618 GND.n612 1.129
R4044 GND.n1886 GND.n1881 1.129
R4045 GND.n1879 GND.n1874 1.129
R4046 GND.n1846 GND.n1842 1.129
R4047 GND.n1840 GND.n1834 1.129
R4048 GND.n1805 GND.n1800 1.129
R4049 GND.n1798 GND.n1793 1.129
R4050 GND.n1765 GND.n1761 1.129
R4051 GND.n1759 GND.n1753 1.129
R4052 GND.n1724 GND.n1719 1.129
R4053 GND.n1717 GND.n1712 1.129
R4054 GND.n1684 GND.n1680 1.129
R4055 GND.n1678 GND.n1672 1.129
R4056 GND.n1643 GND.n1638 1.129
R4057 GND.n1636 GND.n1631 1.129
R4058 GND.n1603 GND.n1599 1.129
R4059 GND.n1597 GND.n1591 1.129
R4060 GND.n1562 GND.n1557 1.129
R4061 GND.n1555 GND.n1550 1.129
R4062 GND.n1522 GND.n1518 1.129
R4063 GND.n1516 GND.n1510 1.129
R4064 GND.n1481 GND.n1476 1.129
R4065 GND.n1474 GND.n1469 1.129
R4066 GND.n1441 GND.n1437 1.129
R4067 GND.n1435 GND.n1429 1.129
R4068 GND.n1400 GND.n1395 1.129
R4069 GND.n1393 GND.n1388 1.129
R4070 GND.n1360 GND.n1356 1.129
R4071 GND.n1354 GND.n1348 1.129
R4072 GND.n1319 GND.n1314 1.129
R4073 GND.n1312 GND.n1307 1.129
R4074 GND.n1279 GND.n1275 1.129
R4075 GND.n1273 GND.n1267 1.129
R4076 GND.n2551 GND.n2546 1.129
R4077 GND.n2544 GND.n2539 1.129
R4078 GND.n2511 GND.n2507 1.129
R4079 GND.n2505 GND.n2499 1.129
R4080 GND.n2470 GND.n2465 1.129
R4081 GND.n2463 GND.n2458 1.129
R4082 GND.n2430 GND.n2426 1.129
R4083 GND.n2424 GND.n2418 1.129
R4084 GND.n2389 GND.n2384 1.129
R4085 GND.n2382 GND.n2377 1.129
R4086 GND.n2349 GND.n2345 1.129
R4087 GND.n2343 GND.n2337 1.129
R4088 GND.n2308 GND.n2303 1.129
R4089 GND.n2301 GND.n2296 1.129
R4090 GND.n2268 GND.n2264 1.129
R4091 GND.n2262 GND.n2256 1.129
R4092 GND.n2227 GND.n2222 1.129
R4093 GND.n2220 GND.n2215 1.129
R4094 GND.n2187 GND.n2183 1.129
R4095 GND.n2181 GND.n2175 1.129
R4096 GND.n2146 GND.n2141 1.129
R4097 GND.n2139 GND.n2134 1.129
R4098 GND.n2106 GND.n2102 1.129
R4099 GND.n2100 GND.n2094 1.129
R4100 GND.n2065 GND.n2060 1.129
R4101 GND.n2058 GND.n2053 1.129
R4102 GND.n2025 GND.n2021 1.129
R4103 GND.n2019 GND.n2013 1.129
R4104 GND.n1984 GND.n1979 1.129
R4105 GND.n1977 GND.n1972 1.129
R4106 GND.n1944 GND.n1940 1.129
R4107 GND.n1938 GND.n1932 1.129
R4108 GND.n3206 GND.n3201 1.129
R4109 GND.n3199 GND.n3194 1.129
R4110 GND.n3166 GND.n3162 1.129
R4111 GND.n3160 GND.n3154 1.129
R4112 GND.n3125 GND.n3120 1.129
R4113 GND.n3118 GND.n3113 1.129
R4114 GND.n3085 GND.n3081 1.129
R4115 GND.n3079 GND.n3073 1.129
R4116 GND.n3044 GND.n3039 1.129
R4117 GND.n3037 GND.n3032 1.129
R4118 GND.n3004 GND.n3000 1.129
R4119 GND.n2998 GND.n2992 1.129
R4120 GND.n2963 GND.n2958 1.129
R4121 GND.n2956 GND.n2951 1.129
R4122 GND.n2923 GND.n2919 1.129
R4123 GND.n2917 GND.n2911 1.129
R4124 GND.n2882 GND.n2877 1.129
R4125 GND.n2875 GND.n2870 1.129
R4126 GND.n2842 GND.n2838 1.129
R4127 GND.n2836 GND.n2830 1.129
R4128 GND.n2801 GND.n2796 1.129
R4129 GND.n2794 GND.n2789 1.129
R4130 GND.n2761 GND.n2757 1.129
R4131 GND.n2755 GND.n2749 1.129
R4132 GND.n2720 GND.n2715 1.129
R4133 GND.n2713 GND.n2708 1.129
R4134 GND.n2680 GND.n2676 1.129
R4135 GND.n2674 GND.n2668 1.129
R4136 GND.n2639 GND.n2634 1.129
R4137 GND.n2632 GND.n2627 1.129
R4138 GND.n2599 GND.n2595 1.129
R4139 GND.n2593 GND.n2587 1.129
R4140 GND.n3861 GND.n3856 1.129
R4141 GND.n3854 GND.n3849 1.129
R4142 GND.n3821 GND.n3817 1.129
R4143 GND.n3815 GND.n3809 1.129
R4144 GND.n3780 GND.n3775 1.129
R4145 GND.n3773 GND.n3768 1.129
R4146 GND.n3740 GND.n3736 1.129
R4147 GND.n3734 GND.n3728 1.129
R4148 GND.n3699 GND.n3694 1.129
R4149 GND.n3692 GND.n3687 1.129
R4150 GND.n3659 GND.n3655 1.129
R4151 GND.n3653 GND.n3647 1.129
R4152 GND.n3618 GND.n3613 1.129
R4153 GND.n3611 GND.n3606 1.129
R4154 GND.n3578 GND.n3574 1.129
R4155 GND.n3572 GND.n3566 1.129
R4156 GND.n3537 GND.n3532 1.129
R4157 GND.n3530 GND.n3525 1.129
R4158 GND.n3497 GND.n3493 1.129
R4159 GND.n3491 GND.n3485 1.129
R4160 GND.n3456 GND.n3451 1.129
R4161 GND.n3449 GND.n3444 1.129
R4162 GND.n3416 GND.n3412 1.129
R4163 GND.n3410 GND.n3404 1.129
R4164 GND.n3375 GND.n3370 1.129
R4165 GND.n3368 GND.n3363 1.129
R4166 GND.n3335 GND.n3331 1.129
R4167 GND.n3329 GND.n3323 1.129
R4168 GND.n3294 GND.n3289 1.129
R4169 GND.n3287 GND.n3282 1.129
R4170 GND.n3254 GND.n3250 1.129
R4171 GND.n3248 GND.n3242 1.129
R4172 GND.n4516 GND.n4511 1.129
R4173 GND.n4509 GND.n4504 1.129
R4174 GND.n4476 GND.n4472 1.129
R4175 GND.n4470 GND.n4464 1.129
R4176 GND.n4435 GND.n4430 1.129
R4177 GND.n4428 GND.n4423 1.129
R4178 GND.n4395 GND.n4391 1.129
R4179 GND.n4389 GND.n4383 1.129
R4180 GND.n4354 GND.n4349 1.129
R4181 GND.n4347 GND.n4342 1.129
R4182 GND.n4314 GND.n4310 1.129
R4183 GND.n4308 GND.n4302 1.129
R4184 GND.n4273 GND.n4268 1.129
R4185 GND.n4266 GND.n4261 1.129
R4186 GND.n4233 GND.n4229 1.129
R4187 GND.n4227 GND.n4221 1.129
R4188 GND.n4192 GND.n4187 1.129
R4189 GND.n4185 GND.n4180 1.129
R4190 GND.n4152 GND.n4148 1.129
R4191 GND.n4146 GND.n4140 1.129
R4192 GND.n4111 GND.n4106 1.129
R4193 GND.n4104 GND.n4099 1.129
R4194 GND.n4071 GND.n4067 1.129
R4195 GND.n4065 GND.n4059 1.129
R4196 GND.n4030 GND.n4025 1.129
R4197 GND.n4023 GND.n4018 1.129
R4198 GND.n3990 GND.n3986 1.129
R4199 GND.n3984 GND.n3978 1.129
R4200 GND.n3949 GND.n3944 1.129
R4201 GND.n3942 GND.n3937 1.129
R4202 GND.n3909 GND.n3905 1.129
R4203 GND.n3903 GND.n3897 1.129
R4204 GND.n5181 GND.n5176 1.129
R4205 GND.n5174 GND.n5169 1.129
R4206 GND.n5141 GND.n5137 1.129
R4207 GND.n5135 GND.n5129 1.129
R4208 GND.n5100 GND.n5095 1.129
R4209 GND.n5093 GND.n5088 1.129
R4210 GND.n5060 GND.n5056 1.129
R4211 GND.n5054 GND.n5048 1.129
R4212 GND.n5019 GND.n5014 1.129
R4213 GND.n5012 GND.n5007 1.129
R4214 GND.n4979 GND.n4975 1.129
R4215 GND.n4973 GND.n4967 1.129
R4216 GND.n4938 GND.n4933 1.129
R4217 GND.n4931 GND.n4926 1.129
R4218 GND.n4898 GND.n4894 1.129
R4219 GND.n4892 GND.n4886 1.129
R4220 GND.n4857 GND.n4852 1.129
R4221 GND.n4850 GND.n4845 1.129
R4222 GND.n4817 GND.n4813 1.129
R4223 GND.n4811 GND.n4805 1.129
R4224 GND.n4776 GND.n4771 1.129
R4225 GND.n4769 GND.n4764 1.129
R4226 GND.n4736 GND.n4732 1.129
R4227 GND.n4730 GND.n4724 1.129
R4228 GND.n4695 GND.n4690 1.129
R4229 GND.n4688 GND.n4683 1.129
R4230 GND.n4655 GND.n4651 1.129
R4231 GND.n4649 GND.n4643 1.129
R4232 GND.n4614 GND.n4609 1.129
R4233 GND.n4607 GND.n4602 1.129
R4234 GND.n4574 GND.n4570 1.129
R4235 GND.n4568 GND.n4562 1.129
R4236 GND GND.n5230 1.031
R4237 GND.n90 GND.n89 0.919
R4238 GND.n90 GND.n49 0.919
R4239 GND.n262 GND.n261 0.919
R4240 GND.n262 GND.n221 0.919
R4241 GND.n181 GND.n180 0.919
R4242 GND.n181 GND.n140 0.919
R4243 GND.n597 GND.n596 0.919
R4244 GND.n597 GND.n556 0.919
R4245 GND.n516 GND.n515 0.919
R4246 GND.n516 GND.n475 0.919
R4247 GND.n435 GND.n434 0.919
R4248 GND.n435 GND.n394 0.919
R4249 GND.n354 GND.n353 0.919
R4250 GND.n354 GND.n313 0.919
R4251 GND.n1258 GND.n1257 0.919
R4252 GND.n1258 GND.n1217 0.919
R4253 GND.n1177 GND.n1176 0.919
R4254 GND.n1177 GND.n1136 0.919
R4255 GND.n1096 GND.n1095 0.919
R4256 GND.n1096 GND.n1055 0.919
R4257 GND.n1015 GND.n1014 0.919
R4258 GND.n1015 GND.n974 0.919
R4259 GND.n934 GND.n933 0.919
R4260 GND.n934 GND.n893 0.919
R4261 GND.n853 GND.n852 0.919
R4262 GND.n853 GND.n812 0.919
R4263 GND.n772 GND.n771 0.919
R4264 GND.n772 GND.n731 0.919
R4265 GND.n691 GND.n690 0.919
R4266 GND.n691 GND.n650 0.919
R4267 GND.n1913 GND.n1912 0.919
R4268 GND.n1913 GND.n1872 0.919
R4269 GND.n1832 GND.n1831 0.919
R4270 GND.n1832 GND.n1791 0.919
R4271 GND.n1751 GND.n1750 0.919
R4272 GND.n1751 GND.n1710 0.919
R4273 GND.n1670 GND.n1669 0.919
R4274 GND.n1670 GND.n1629 0.919
R4275 GND.n1589 GND.n1588 0.919
R4276 GND.n1589 GND.n1548 0.919
R4277 GND.n1508 GND.n1507 0.919
R4278 GND.n1508 GND.n1467 0.919
R4279 GND.n1427 GND.n1426 0.919
R4280 GND.n1427 GND.n1386 0.919
R4281 GND.n1346 GND.n1345 0.919
R4282 GND.n1346 GND.n1305 0.919
R4283 GND.n2578 GND.n2577 0.919
R4284 GND.n2578 GND.n2537 0.919
R4285 GND.n2497 GND.n2496 0.919
R4286 GND.n2497 GND.n2456 0.919
R4287 GND.n2416 GND.n2415 0.919
R4288 GND.n2416 GND.n2375 0.919
R4289 GND.n2335 GND.n2334 0.919
R4290 GND.n2335 GND.n2294 0.919
R4291 GND.n2254 GND.n2253 0.919
R4292 GND.n2254 GND.n2213 0.919
R4293 GND.n2173 GND.n2172 0.919
R4294 GND.n2173 GND.n2132 0.919
R4295 GND.n2092 GND.n2091 0.919
R4296 GND.n2092 GND.n2051 0.919
R4297 GND.n2011 GND.n2010 0.919
R4298 GND.n2011 GND.n1970 0.919
R4299 GND.n3233 GND.n3232 0.919
R4300 GND.n3233 GND.n3192 0.919
R4301 GND.n3152 GND.n3151 0.919
R4302 GND.n3152 GND.n3111 0.919
R4303 GND.n3071 GND.n3070 0.919
R4304 GND.n3071 GND.n3030 0.919
R4305 GND.n2990 GND.n2989 0.919
R4306 GND.n2990 GND.n2949 0.919
R4307 GND.n2909 GND.n2908 0.919
R4308 GND.n2909 GND.n2868 0.919
R4309 GND.n2828 GND.n2827 0.919
R4310 GND.n2828 GND.n2787 0.919
R4311 GND.n2747 GND.n2746 0.919
R4312 GND.n2747 GND.n2706 0.919
R4313 GND.n2666 GND.n2665 0.919
R4314 GND.n2666 GND.n2625 0.919
R4315 GND.n3888 GND.n3887 0.919
R4316 GND.n3888 GND.n3847 0.919
R4317 GND.n3807 GND.n3806 0.919
R4318 GND.n3807 GND.n3766 0.919
R4319 GND.n3726 GND.n3725 0.919
R4320 GND.n3726 GND.n3685 0.919
R4321 GND.n3645 GND.n3644 0.919
R4322 GND.n3645 GND.n3604 0.919
R4323 GND.n3564 GND.n3563 0.919
R4324 GND.n3564 GND.n3523 0.919
R4325 GND.n3483 GND.n3482 0.919
R4326 GND.n3483 GND.n3442 0.919
R4327 GND.n3402 GND.n3401 0.919
R4328 GND.n3402 GND.n3361 0.919
R4329 GND.n3321 GND.n3320 0.919
R4330 GND.n3321 GND.n3280 0.919
R4331 GND.n4543 GND.n4542 0.919
R4332 GND.n4543 GND.n4502 0.919
R4333 GND.n4462 GND.n4461 0.919
R4334 GND.n4462 GND.n4421 0.919
R4335 GND.n4381 GND.n4380 0.919
R4336 GND.n4381 GND.n4340 0.919
R4337 GND.n4300 GND.n4299 0.919
R4338 GND.n4300 GND.n4259 0.919
R4339 GND.n4219 GND.n4218 0.919
R4340 GND.n4219 GND.n4178 0.919
R4341 GND.n4138 GND.n4137 0.919
R4342 GND.n4138 GND.n4097 0.919
R4343 GND.n4057 GND.n4056 0.919
R4344 GND.n4057 GND.n4016 0.919
R4345 GND.n3976 GND.n3975 0.919
R4346 GND.n3976 GND.n3935 0.919
R4347 GND.n5208 GND.n5207 0.919
R4348 GND.n5208 GND.n5167 0.919
R4349 GND.n5127 GND.n5126 0.919
R4350 GND.n5127 GND.n5086 0.919
R4351 GND.n5046 GND.n5045 0.919
R4352 GND.n5046 GND.n5005 0.919
R4353 GND.n4965 GND.n4964 0.919
R4354 GND.n4965 GND.n4924 0.919
R4355 GND.n4884 GND.n4883 0.919
R4356 GND.n4884 GND.n4843 0.919
R4357 GND.n4803 GND.n4802 0.919
R4358 GND.n4803 GND.n4762 0.919
R4359 GND.n4722 GND.n4721 0.919
R4360 GND.n4722 GND.n4681 0.919
R4361 GND.n4641 GND.n4640 0.919
R4362 GND.n4641 GND.n4600 0.919
R4363 GND.n263 GND.n181 0.803
R4364 GND.n598 GND.n516 0.803
R4365 GND.n599 GND.n435 0.803
R4366 GND.n600 GND.n354 0.803
R4367 GND.n1259 GND.n1177 0.803
R4368 GND.n1260 GND.n1096 0.803
R4369 GND.n1261 GND.n1015 0.803
R4370 GND.n1262 GND.n934 0.803
R4371 GND.n1263 GND.n853 0.803
R4372 GND.n1264 GND.n772 0.803
R4373 GND.n1265 GND.n691 0.803
R4374 GND.n1914 GND.n1832 0.803
R4375 GND.n1915 GND.n1751 0.803
R4376 GND.n1916 GND.n1670 0.803
R4377 GND.n1917 GND.n1589 0.803
R4378 GND.n1918 GND.n1508 0.803
R4379 GND.n1919 GND.n1427 0.803
R4380 GND.n1920 GND.n1346 0.803
R4381 GND.n2579 GND.n2497 0.803
R4382 GND.n2580 GND.n2416 0.803
R4383 GND.n2581 GND.n2335 0.803
R4384 GND.n2582 GND.n2254 0.803
R4385 GND.n2583 GND.n2173 0.803
R4386 GND.n2584 GND.n2092 0.803
R4387 GND.n2585 GND.n2011 0.803
R4388 GND.n3234 GND.n3152 0.803
R4389 GND.n3235 GND.n3071 0.803
R4390 GND.n3236 GND.n2990 0.803
R4391 GND.n3237 GND.n2909 0.803
R4392 GND.n3238 GND.n2828 0.803
R4393 GND.n3239 GND.n2747 0.803
R4394 GND.n3240 GND.n2666 0.803
R4395 GND.n3889 GND.n3807 0.803
R4396 GND.n3890 GND.n3726 0.803
R4397 GND.n3891 GND.n3645 0.803
R4398 GND.n3892 GND.n3564 0.803
R4399 GND.n3893 GND.n3483 0.803
R4400 GND.n3894 GND.n3402 0.803
R4401 GND.n3895 GND.n3321 0.803
R4402 GND.n4544 GND.n4462 0.803
R4403 GND.n4545 GND.n4381 0.803
R4404 GND.n4546 GND.n4300 0.803
R4405 GND.n4547 GND.n4219 0.803
R4406 GND.n4548 GND.n4138 0.803
R4407 GND.n4549 GND.n4057 0.803
R4408 GND.n4550 GND.n3976 0.803
R4409 GND.n5209 GND.n5127 0.803
R4410 GND.n5210 GND.n5046 0.803
R4411 GND.n5211 GND.n4965 0.803
R4412 GND.n5212 GND.n4884 0.803
R4413 GND.n5213 GND.n4803 0.803
R4414 GND.n5214 GND.n4722 0.803
R4415 GND.n5215 GND.n4641 0.803
R4416 GND.n3 GND.n1 0.656
R4417 GND.n94 GND.n92 0.656
R4418 GND.n267 GND.n265 0.656
R4419 GND.n604 GND.n602 0.656
R4420 GND.n1924 GND.n1922 0.656
R4421 GND.n4554 GND.n4552 0.656
R4422 GND.n5223 GND.n5222 0.614
R4423 GND.n5220 GND.n5219 0.614
R4424 GND.n5219 GND.n5218 0.614
R4425 GND.n5218 GND.n5217 0.614
R4426 GND.n5216 GND.n5215 0.611
R4427 GND.n599 GND.n598 0.575
R4428 GND.n600 GND.n599 0.575
R4429 GND.n1260 GND.n1259 0.575
R4430 GND.n1261 GND.n1260 0.575
R4431 GND.n1262 GND.n1261 0.575
R4432 GND.n1263 GND.n1262 0.575
R4433 GND.n1264 GND.n1263 0.575
R4434 GND.n1265 GND.n1264 0.575
R4435 GND.n1915 GND.n1914 0.575
R4436 GND.n1916 GND.n1915 0.575
R4437 GND.n1917 GND.n1916 0.575
R4438 GND.n1918 GND.n1917 0.575
R4439 GND.n1919 GND.n1918 0.575
R4440 GND.n1920 GND.n1919 0.575
R4441 GND.n2580 GND.n2579 0.575
R4442 GND.n2581 GND.n2580 0.575
R4443 GND.n2582 GND.n2581 0.575
R4444 GND.n2583 GND.n2582 0.575
R4445 GND.n2584 GND.n2583 0.575
R4446 GND.n2585 GND.n2584 0.575
R4447 GND.n3235 GND.n3234 0.575
R4448 GND.n3236 GND.n3235 0.575
R4449 GND.n3237 GND.n3236 0.575
R4450 GND.n3238 GND.n3237 0.575
R4451 GND.n3239 GND.n3238 0.575
R4452 GND.n3240 GND.n3239 0.575
R4453 GND.n3890 GND.n3889 0.575
R4454 GND.n3891 GND.n3890 0.575
R4455 GND.n3892 GND.n3891 0.575
R4456 GND.n3893 GND.n3892 0.575
R4457 GND.n3894 GND.n3893 0.575
R4458 GND.n3895 GND.n3894 0.575
R4459 GND.n4545 GND.n4544 0.575
R4460 GND.n4546 GND.n4545 0.575
R4461 GND.n4547 GND.n4546 0.575
R4462 GND.n4548 GND.n4547 0.575
R4463 GND.n4549 GND.n4548 0.575
R4464 GND.n4550 GND.n4549 0.575
R4465 GND.n5210 GND.n5209 0.575
R4466 GND.n5211 GND.n5210 0.575
R4467 GND.n5212 GND.n5211 0.575
R4468 GND.n5213 GND.n5212 0.575
R4469 GND.n5214 GND.n5213 0.575
R4470 GND.n5215 GND.n5214 0.575
R4471 GND.n5229 GND.n5228 0.406
R4472 GND.n5227 GND.n5226 0.406
R4473 GND.n5225 GND.n5224 0.406
R4474 GND.n5222 GND.n5221 0.406
R4475 GND.n5217 GND.n5216 0.406
R4476 GND.n5227 GND.n263 0.403
R4477 GND.n5225 GND.n600 0.403
R4478 GND.n5223 GND.n1265 0.403
R4479 GND.n5222 GND.n1920 0.403
R4480 GND.n5220 GND.n2585 0.403
R4481 GND.n5219 GND.n3240 0.403
R4482 GND.n5218 GND.n3895 0.403
R4483 GND.n5217 GND.n4550 0.403
R4484 GND.n74 GND.n69 0.376
R4485 GND.n83 GND.n77 0.376
R4486 GND.n34 GND.n29 0.376
R4487 GND.n43 GND.n37 0.376
R4488 GND.n246 GND.n241 0.376
R4489 GND.n255 GND.n249 0.376
R4490 GND.n206 GND.n201 0.376
R4491 GND.n215 GND.n209 0.376
R4492 GND.n165 GND.n160 0.376
R4493 GND.n174 GND.n168 0.376
R4494 GND.n125 GND.n120 0.376
R4495 GND.n134 GND.n128 0.376
R4496 GND.n581 GND.n576 0.376
R4497 GND.n590 GND.n584 0.376
R4498 GND.n541 GND.n536 0.376
R4499 GND.n550 GND.n544 0.376
R4500 GND.n500 GND.n495 0.376
R4501 GND.n509 GND.n503 0.376
R4502 GND.n460 GND.n455 0.376
R4503 GND.n469 GND.n463 0.376
R4504 GND.n419 GND.n414 0.376
R4505 GND.n428 GND.n422 0.376
R4506 GND.n379 GND.n374 0.376
R4507 GND.n388 GND.n382 0.376
R4508 GND.n338 GND.n333 0.376
R4509 GND.n347 GND.n341 0.376
R4510 GND.n298 GND.n293 0.376
R4511 GND.n307 GND.n301 0.376
R4512 GND.n1242 GND.n1237 0.376
R4513 GND.n1251 GND.n1245 0.376
R4514 GND.n1202 GND.n1197 0.376
R4515 GND.n1211 GND.n1205 0.376
R4516 GND.n1161 GND.n1156 0.376
R4517 GND.n1170 GND.n1164 0.376
R4518 GND.n1121 GND.n1116 0.376
R4519 GND.n1130 GND.n1124 0.376
R4520 GND.n1080 GND.n1075 0.376
R4521 GND.n1089 GND.n1083 0.376
R4522 GND.n1040 GND.n1035 0.376
R4523 GND.n1049 GND.n1043 0.376
R4524 GND.n999 GND.n994 0.376
R4525 GND.n1008 GND.n1002 0.376
R4526 GND.n959 GND.n954 0.376
R4527 GND.n968 GND.n962 0.376
R4528 GND.n918 GND.n913 0.376
R4529 GND.n927 GND.n921 0.376
R4530 GND.n878 GND.n873 0.376
R4531 GND.n887 GND.n881 0.376
R4532 GND.n837 GND.n832 0.376
R4533 GND.n846 GND.n840 0.376
R4534 GND.n797 GND.n792 0.376
R4535 GND.n806 GND.n800 0.376
R4536 GND.n756 GND.n751 0.376
R4537 GND.n765 GND.n759 0.376
R4538 GND.n716 GND.n711 0.376
R4539 GND.n725 GND.n719 0.376
R4540 GND.n675 GND.n670 0.376
R4541 GND.n684 GND.n678 0.376
R4542 GND.n635 GND.n630 0.376
R4543 GND.n644 GND.n638 0.376
R4544 GND.n1897 GND.n1892 0.376
R4545 GND.n1906 GND.n1900 0.376
R4546 GND.n1857 GND.n1852 0.376
R4547 GND.n1866 GND.n1860 0.376
R4548 GND.n1816 GND.n1811 0.376
R4549 GND.n1825 GND.n1819 0.376
R4550 GND.n1776 GND.n1771 0.376
R4551 GND.n1785 GND.n1779 0.376
R4552 GND.n1735 GND.n1730 0.376
R4553 GND.n1744 GND.n1738 0.376
R4554 GND.n1695 GND.n1690 0.376
R4555 GND.n1704 GND.n1698 0.376
R4556 GND.n1654 GND.n1649 0.376
R4557 GND.n1663 GND.n1657 0.376
R4558 GND.n1614 GND.n1609 0.376
R4559 GND.n1623 GND.n1617 0.376
R4560 GND.n1573 GND.n1568 0.376
R4561 GND.n1582 GND.n1576 0.376
R4562 GND.n1533 GND.n1528 0.376
R4563 GND.n1542 GND.n1536 0.376
R4564 GND.n1492 GND.n1487 0.376
R4565 GND.n1501 GND.n1495 0.376
R4566 GND.n1452 GND.n1447 0.376
R4567 GND.n1461 GND.n1455 0.376
R4568 GND.n1411 GND.n1406 0.376
R4569 GND.n1420 GND.n1414 0.376
R4570 GND.n1371 GND.n1366 0.376
R4571 GND.n1380 GND.n1374 0.376
R4572 GND.n1330 GND.n1325 0.376
R4573 GND.n1339 GND.n1333 0.376
R4574 GND.n1290 GND.n1285 0.376
R4575 GND.n1299 GND.n1293 0.376
R4576 GND.n2562 GND.n2557 0.376
R4577 GND.n2571 GND.n2565 0.376
R4578 GND.n2522 GND.n2517 0.376
R4579 GND.n2531 GND.n2525 0.376
R4580 GND.n2481 GND.n2476 0.376
R4581 GND.n2490 GND.n2484 0.376
R4582 GND.n2441 GND.n2436 0.376
R4583 GND.n2450 GND.n2444 0.376
R4584 GND.n2400 GND.n2395 0.376
R4585 GND.n2409 GND.n2403 0.376
R4586 GND.n2360 GND.n2355 0.376
R4587 GND.n2369 GND.n2363 0.376
R4588 GND.n2319 GND.n2314 0.376
R4589 GND.n2328 GND.n2322 0.376
R4590 GND.n2279 GND.n2274 0.376
R4591 GND.n2288 GND.n2282 0.376
R4592 GND.n2238 GND.n2233 0.376
R4593 GND.n2247 GND.n2241 0.376
R4594 GND.n2198 GND.n2193 0.376
R4595 GND.n2207 GND.n2201 0.376
R4596 GND.n2157 GND.n2152 0.376
R4597 GND.n2166 GND.n2160 0.376
R4598 GND.n2117 GND.n2112 0.376
R4599 GND.n2126 GND.n2120 0.376
R4600 GND.n2076 GND.n2071 0.376
R4601 GND.n2085 GND.n2079 0.376
R4602 GND.n2036 GND.n2031 0.376
R4603 GND.n2045 GND.n2039 0.376
R4604 GND.n1995 GND.n1990 0.376
R4605 GND.n2004 GND.n1998 0.376
R4606 GND.n1955 GND.n1950 0.376
R4607 GND.n1964 GND.n1958 0.376
R4608 GND.n3217 GND.n3212 0.376
R4609 GND.n3226 GND.n3220 0.376
R4610 GND.n3177 GND.n3172 0.376
R4611 GND.n3186 GND.n3180 0.376
R4612 GND.n3136 GND.n3131 0.376
R4613 GND.n3145 GND.n3139 0.376
R4614 GND.n3096 GND.n3091 0.376
R4615 GND.n3105 GND.n3099 0.376
R4616 GND.n3055 GND.n3050 0.376
R4617 GND.n3064 GND.n3058 0.376
R4618 GND.n3015 GND.n3010 0.376
R4619 GND.n3024 GND.n3018 0.376
R4620 GND.n2974 GND.n2969 0.376
R4621 GND.n2983 GND.n2977 0.376
R4622 GND.n2934 GND.n2929 0.376
R4623 GND.n2943 GND.n2937 0.376
R4624 GND.n2893 GND.n2888 0.376
R4625 GND.n2902 GND.n2896 0.376
R4626 GND.n2853 GND.n2848 0.376
R4627 GND.n2862 GND.n2856 0.376
R4628 GND.n2812 GND.n2807 0.376
R4629 GND.n2821 GND.n2815 0.376
R4630 GND.n2772 GND.n2767 0.376
R4631 GND.n2781 GND.n2775 0.376
R4632 GND.n2731 GND.n2726 0.376
R4633 GND.n2740 GND.n2734 0.376
R4634 GND.n2691 GND.n2686 0.376
R4635 GND.n2700 GND.n2694 0.376
R4636 GND.n2650 GND.n2645 0.376
R4637 GND.n2659 GND.n2653 0.376
R4638 GND.n2610 GND.n2605 0.376
R4639 GND.n2619 GND.n2613 0.376
R4640 GND.n3872 GND.n3867 0.376
R4641 GND.n3881 GND.n3875 0.376
R4642 GND.n3832 GND.n3827 0.376
R4643 GND.n3841 GND.n3835 0.376
R4644 GND.n3791 GND.n3786 0.376
R4645 GND.n3800 GND.n3794 0.376
R4646 GND.n3751 GND.n3746 0.376
R4647 GND.n3760 GND.n3754 0.376
R4648 GND.n3710 GND.n3705 0.376
R4649 GND.n3719 GND.n3713 0.376
R4650 GND.n3670 GND.n3665 0.376
R4651 GND.n3679 GND.n3673 0.376
R4652 GND.n3629 GND.n3624 0.376
R4653 GND.n3638 GND.n3632 0.376
R4654 GND.n3589 GND.n3584 0.376
R4655 GND.n3598 GND.n3592 0.376
R4656 GND.n3548 GND.n3543 0.376
R4657 GND.n3557 GND.n3551 0.376
R4658 GND.n3508 GND.n3503 0.376
R4659 GND.n3517 GND.n3511 0.376
R4660 GND.n3467 GND.n3462 0.376
R4661 GND.n3476 GND.n3470 0.376
R4662 GND.n3427 GND.n3422 0.376
R4663 GND.n3436 GND.n3430 0.376
R4664 GND.n3386 GND.n3381 0.376
R4665 GND.n3395 GND.n3389 0.376
R4666 GND.n3346 GND.n3341 0.376
R4667 GND.n3355 GND.n3349 0.376
R4668 GND.n3305 GND.n3300 0.376
R4669 GND.n3314 GND.n3308 0.376
R4670 GND.n3265 GND.n3260 0.376
R4671 GND.n3274 GND.n3268 0.376
R4672 GND.n4527 GND.n4522 0.376
R4673 GND.n4536 GND.n4530 0.376
R4674 GND.n4487 GND.n4482 0.376
R4675 GND.n4496 GND.n4490 0.376
R4676 GND.n4446 GND.n4441 0.376
R4677 GND.n4455 GND.n4449 0.376
R4678 GND.n4406 GND.n4401 0.376
R4679 GND.n4415 GND.n4409 0.376
R4680 GND.n4365 GND.n4360 0.376
R4681 GND.n4374 GND.n4368 0.376
R4682 GND.n4325 GND.n4320 0.376
R4683 GND.n4334 GND.n4328 0.376
R4684 GND.n4284 GND.n4279 0.376
R4685 GND.n4293 GND.n4287 0.376
R4686 GND.n4244 GND.n4239 0.376
R4687 GND.n4253 GND.n4247 0.376
R4688 GND.n4203 GND.n4198 0.376
R4689 GND.n4212 GND.n4206 0.376
R4690 GND.n4163 GND.n4158 0.376
R4691 GND.n4172 GND.n4166 0.376
R4692 GND.n4122 GND.n4117 0.376
R4693 GND.n4131 GND.n4125 0.376
R4694 GND.n4082 GND.n4077 0.376
R4695 GND.n4091 GND.n4085 0.376
R4696 GND.n4041 GND.n4036 0.376
R4697 GND.n4050 GND.n4044 0.376
R4698 GND.n4001 GND.n3996 0.376
R4699 GND.n4010 GND.n4004 0.376
R4700 GND.n3960 GND.n3955 0.376
R4701 GND.n3969 GND.n3963 0.376
R4702 GND.n3920 GND.n3915 0.376
R4703 GND.n3929 GND.n3923 0.376
R4704 GND.n5192 GND.n5187 0.376
R4705 GND.n5201 GND.n5195 0.376
R4706 GND.n5152 GND.n5147 0.376
R4707 GND.n5161 GND.n5155 0.376
R4708 GND.n5111 GND.n5106 0.376
R4709 GND.n5120 GND.n5114 0.376
R4710 GND.n5071 GND.n5066 0.376
R4711 GND.n5080 GND.n5074 0.376
R4712 GND.n5030 GND.n5025 0.376
R4713 GND.n5039 GND.n5033 0.376
R4714 GND.n4990 GND.n4985 0.376
R4715 GND.n4999 GND.n4993 0.376
R4716 GND.n4949 GND.n4944 0.376
R4717 GND.n4958 GND.n4952 0.376
R4718 GND.n4909 GND.n4904 0.376
R4719 GND.n4918 GND.n4912 0.376
R4720 GND.n4868 GND.n4863 0.376
R4721 GND.n4877 GND.n4871 0.376
R4722 GND.n4828 GND.n4823 0.376
R4723 GND.n4837 GND.n4831 0.376
R4724 GND.n4787 GND.n4782 0.376
R4725 GND.n4796 GND.n4790 0.376
R4726 GND.n4747 GND.n4742 0.376
R4727 GND.n4756 GND.n4750 0.376
R4728 GND.n4706 GND.n4701 0.376
R4729 GND.n4715 GND.n4709 0.376
R4730 GND.n4666 GND.n4661 0.376
R4731 GND.n4675 GND.n4669 0.376
R4732 GND.n4625 GND.n4620 0.376
R4733 GND.n4634 GND.n4628 0.376
R4734 GND.n4585 GND.n4580 0.376
R4735 GND.n4594 GND.n4588 0.376
R4736 GND.n5230 GND.n5229 0.208
R4737 GND.n5228 GND.n5227 0.208
R4738 GND.n5226 GND.n5225 0.208
R4739 GND.n5224 GND.n5223 0.208
R4740 GND.n5221 GND.n5220 0.208
R4741 GND.n4 GND.n3 0.152
R4742 GND.n95 GND.n94 0.152
R4743 GND.n268 GND.n267 0.152
R4744 GND.n605 GND.n604 0.152
R4745 GND.n1925 GND.n1924 0.152
R4746 GND.n4555 GND.n4554 0.152
R4747 GND.n84 GND.n75 0.15
R4748 GND.n44 GND.n35 0.15
R4749 GND.n256 GND.n247 0.15
R4750 GND.n216 GND.n207 0.15
R4751 GND.n175 GND.n166 0.15
R4752 GND.n135 GND.n126 0.15
R4753 GND.n591 GND.n582 0.15
R4754 GND.n551 GND.n542 0.15
R4755 GND.n510 GND.n501 0.15
R4756 GND.n470 GND.n461 0.15
R4757 GND.n429 GND.n420 0.15
R4758 GND.n389 GND.n380 0.15
R4759 GND.n348 GND.n339 0.15
R4760 GND.n308 GND.n299 0.15
R4761 GND.n1252 GND.n1243 0.15
R4762 GND.n1212 GND.n1203 0.15
R4763 GND.n1171 GND.n1162 0.15
R4764 GND.n1131 GND.n1122 0.15
R4765 GND.n1090 GND.n1081 0.15
R4766 GND.n1050 GND.n1041 0.15
R4767 GND.n1009 GND.n1000 0.15
R4768 GND.n969 GND.n960 0.15
R4769 GND.n928 GND.n919 0.15
R4770 GND.n888 GND.n879 0.15
R4771 GND.n847 GND.n838 0.15
R4772 GND.n807 GND.n798 0.15
R4773 GND.n766 GND.n757 0.15
R4774 GND.n726 GND.n717 0.15
R4775 GND.n685 GND.n676 0.15
R4776 GND.n645 GND.n636 0.15
R4777 GND.n1907 GND.n1898 0.15
R4778 GND.n1867 GND.n1858 0.15
R4779 GND.n1826 GND.n1817 0.15
R4780 GND.n1786 GND.n1777 0.15
R4781 GND.n1745 GND.n1736 0.15
R4782 GND.n1705 GND.n1696 0.15
R4783 GND.n1664 GND.n1655 0.15
R4784 GND.n1624 GND.n1615 0.15
R4785 GND.n1583 GND.n1574 0.15
R4786 GND.n1543 GND.n1534 0.15
R4787 GND.n1502 GND.n1493 0.15
R4788 GND.n1462 GND.n1453 0.15
R4789 GND.n1421 GND.n1412 0.15
R4790 GND.n1381 GND.n1372 0.15
R4791 GND.n1340 GND.n1331 0.15
R4792 GND.n1300 GND.n1291 0.15
R4793 GND.n2572 GND.n2563 0.15
R4794 GND.n2532 GND.n2523 0.15
R4795 GND.n2491 GND.n2482 0.15
R4796 GND.n2451 GND.n2442 0.15
R4797 GND.n2410 GND.n2401 0.15
R4798 GND.n2370 GND.n2361 0.15
R4799 GND.n2329 GND.n2320 0.15
R4800 GND.n2289 GND.n2280 0.15
R4801 GND.n2248 GND.n2239 0.15
R4802 GND.n2208 GND.n2199 0.15
R4803 GND.n2167 GND.n2158 0.15
R4804 GND.n2127 GND.n2118 0.15
R4805 GND.n2086 GND.n2077 0.15
R4806 GND.n2046 GND.n2037 0.15
R4807 GND.n2005 GND.n1996 0.15
R4808 GND.n1965 GND.n1956 0.15
R4809 GND.n3227 GND.n3218 0.15
R4810 GND.n3187 GND.n3178 0.15
R4811 GND.n3146 GND.n3137 0.15
R4812 GND.n3106 GND.n3097 0.15
R4813 GND.n3065 GND.n3056 0.15
R4814 GND.n3025 GND.n3016 0.15
R4815 GND.n2984 GND.n2975 0.15
R4816 GND.n2944 GND.n2935 0.15
R4817 GND.n2903 GND.n2894 0.15
R4818 GND.n2863 GND.n2854 0.15
R4819 GND.n2822 GND.n2813 0.15
R4820 GND.n2782 GND.n2773 0.15
R4821 GND.n2741 GND.n2732 0.15
R4822 GND.n2701 GND.n2692 0.15
R4823 GND.n2660 GND.n2651 0.15
R4824 GND.n2620 GND.n2611 0.15
R4825 GND.n3882 GND.n3873 0.15
R4826 GND.n3842 GND.n3833 0.15
R4827 GND.n3801 GND.n3792 0.15
R4828 GND.n3761 GND.n3752 0.15
R4829 GND.n3720 GND.n3711 0.15
R4830 GND.n3680 GND.n3671 0.15
R4831 GND.n3639 GND.n3630 0.15
R4832 GND.n3599 GND.n3590 0.15
R4833 GND.n3558 GND.n3549 0.15
R4834 GND.n3518 GND.n3509 0.15
R4835 GND.n3477 GND.n3468 0.15
R4836 GND.n3437 GND.n3428 0.15
R4837 GND.n3396 GND.n3387 0.15
R4838 GND.n3356 GND.n3347 0.15
R4839 GND.n3315 GND.n3306 0.15
R4840 GND.n3275 GND.n3266 0.15
R4841 GND.n4537 GND.n4528 0.15
R4842 GND.n4497 GND.n4488 0.15
R4843 GND.n4456 GND.n4447 0.15
R4844 GND.n4416 GND.n4407 0.15
R4845 GND.n4375 GND.n4366 0.15
R4846 GND.n4335 GND.n4326 0.15
R4847 GND.n4294 GND.n4285 0.15
R4848 GND.n4254 GND.n4245 0.15
R4849 GND.n4213 GND.n4204 0.15
R4850 GND.n4173 GND.n4164 0.15
R4851 GND.n4132 GND.n4123 0.15
R4852 GND.n4092 GND.n4083 0.15
R4853 GND.n4051 GND.n4042 0.15
R4854 GND.n4011 GND.n4002 0.15
R4855 GND.n3970 GND.n3961 0.15
R4856 GND.n3930 GND.n3921 0.15
R4857 GND.n5202 GND.n5193 0.15
R4858 GND.n5162 GND.n5153 0.15
R4859 GND.n5121 GND.n5112 0.15
R4860 GND.n5081 GND.n5072 0.15
R4861 GND.n5040 GND.n5031 0.15
R4862 GND.n5000 GND.n4991 0.15
R4863 GND.n4959 GND.n4950 0.15
R4864 GND.n4919 GND.n4910 0.15
R4865 GND.n4878 GND.n4869 0.15
R4866 GND.n4838 GND.n4829 0.15
R4867 GND.n4797 GND.n4788 0.15
R4868 GND.n4757 GND.n4748 0.15
R4869 GND.n4716 GND.n4707 0.15
R4870 GND.n4676 GND.n4667 0.15
R4871 GND.n4635 GND.n4626 0.15
R4872 GND.n4595 GND.n4586 0.15
R4873 GND.n89 GND.n88 0.125
R4874 GND.n49 GND.n48 0.125
R4875 GND.n261 GND.n260 0.125
R4876 GND.n221 GND.n220 0.125
R4877 GND.n180 GND.n179 0.125
R4878 GND.n140 GND.n139 0.125
R4879 GND.n596 GND.n595 0.125
R4880 GND.n556 GND.n555 0.125
R4881 GND.n515 GND.n514 0.125
R4882 GND.n475 GND.n474 0.125
R4883 GND.n434 GND.n433 0.125
R4884 GND.n394 GND.n393 0.125
R4885 GND.n353 GND.n352 0.125
R4886 GND.n313 GND.n312 0.125
R4887 GND.n1257 GND.n1256 0.125
R4888 GND.n1217 GND.n1216 0.125
R4889 GND.n1176 GND.n1175 0.125
R4890 GND.n1136 GND.n1135 0.125
R4891 GND.n1095 GND.n1094 0.125
R4892 GND.n1055 GND.n1054 0.125
R4893 GND.n1014 GND.n1013 0.125
R4894 GND.n974 GND.n973 0.125
R4895 GND.n933 GND.n932 0.125
R4896 GND.n893 GND.n892 0.125
R4897 GND.n852 GND.n851 0.125
R4898 GND.n812 GND.n811 0.125
R4899 GND.n771 GND.n770 0.125
R4900 GND.n731 GND.n730 0.125
R4901 GND.n690 GND.n689 0.125
R4902 GND.n650 GND.n649 0.125
R4903 GND.n1912 GND.n1911 0.125
R4904 GND.n1872 GND.n1871 0.125
R4905 GND.n1831 GND.n1830 0.125
R4906 GND.n1791 GND.n1790 0.125
R4907 GND.n1750 GND.n1749 0.125
R4908 GND.n1710 GND.n1709 0.125
R4909 GND.n1669 GND.n1668 0.125
R4910 GND.n1629 GND.n1628 0.125
R4911 GND.n1588 GND.n1587 0.125
R4912 GND.n1548 GND.n1547 0.125
R4913 GND.n1507 GND.n1506 0.125
R4914 GND.n1467 GND.n1466 0.125
R4915 GND.n1426 GND.n1425 0.125
R4916 GND.n1386 GND.n1385 0.125
R4917 GND.n1345 GND.n1344 0.125
R4918 GND.n1305 GND.n1304 0.125
R4919 GND.n2577 GND.n2576 0.125
R4920 GND.n2537 GND.n2536 0.125
R4921 GND.n2496 GND.n2495 0.125
R4922 GND.n2456 GND.n2455 0.125
R4923 GND.n2415 GND.n2414 0.125
R4924 GND.n2375 GND.n2374 0.125
R4925 GND.n2334 GND.n2333 0.125
R4926 GND.n2294 GND.n2293 0.125
R4927 GND.n2253 GND.n2252 0.125
R4928 GND.n2213 GND.n2212 0.125
R4929 GND.n2172 GND.n2171 0.125
R4930 GND.n2132 GND.n2131 0.125
R4931 GND.n2091 GND.n2090 0.125
R4932 GND.n2051 GND.n2050 0.125
R4933 GND.n2010 GND.n2009 0.125
R4934 GND.n1970 GND.n1969 0.125
R4935 GND.n3232 GND.n3231 0.125
R4936 GND.n3192 GND.n3191 0.125
R4937 GND.n3151 GND.n3150 0.125
R4938 GND.n3111 GND.n3110 0.125
R4939 GND.n3070 GND.n3069 0.125
R4940 GND.n3030 GND.n3029 0.125
R4941 GND.n2989 GND.n2988 0.125
R4942 GND.n2949 GND.n2948 0.125
R4943 GND.n2908 GND.n2907 0.125
R4944 GND.n2868 GND.n2867 0.125
R4945 GND.n2827 GND.n2826 0.125
R4946 GND.n2787 GND.n2786 0.125
R4947 GND.n2746 GND.n2745 0.125
R4948 GND.n2706 GND.n2705 0.125
R4949 GND.n2665 GND.n2664 0.125
R4950 GND.n2625 GND.n2624 0.125
R4951 GND.n3887 GND.n3886 0.125
R4952 GND.n3847 GND.n3846 0.125
R4953 GND.n3806 GND.n3805 0.125
R4954 GND.n3766 GND.n3765 0.125
R4955 GND.n3725 GND.n3724 0.125
R4956 GND.n3685 GND.n3684 0.125
R4957 GND.n3644 GND.n3643 0.125
R4958 GND.n3604 GND.n3603 0.125
R4959 GND.n3563 GND.n3562 0.125
R4960 GND.n3523 GND.n3522 0.125
R4961 GND.n3482 GND.n3481 0.125
R4962 GND.n3442 GND.n3441 0.125
R4963 GND.n3401 GND.n3400 0.125
R4964 GND.n3361 GND.n3360 0.125
R4965 GND.n3320 GND.n3319 0.125
R4966 GND.n3280 GND.n3279 0.125
R4967 GND.n4542 GND.n4541 0.125
R4968 GND.n4502 GND.n4501 0.125
R4969 GND.n4461 GND.n4460 0.125
R4970 GND.n4421 GND.n4420 0.125
R4971 GND.n4380 GND.n4379 0.125
R4972 GND.n4340 GND.n4339 0.125
R4973 GND.n4299 GND.n4298 0.125
R4974 GND.n4259 GND.n4258 0.125
R4975 GND.n4218 GND.n4217 0.125
R4976 GND.n4178 GND.n4177 0.125
R4977 GND.n4137 GND.n4136 0.125
R4978 GND.n4097 GND.n4096 0.125
R4979 GND.n4056 GND.n4055 0.125
R4980 GND.n4016 GND.n4015 0.125
R4981 GND.n3975 GND.n3974 0.125
R4982 GND.n3935 GND.n3934 0.125
R4983 GND.n5207 GND.n5206 0.125
R4984 GND.n5167 GND.n5166 0.125
R4985 GND.n5126 GND.n5125 0.125
R4986 GND.n5086 GND.n5085 0.125
R4987 GND.n5045 GND.n5044 0.125
R4988 GND.n5005 GND.n5004 0.125
R4989 GND.n4964 GND.n4963 0.125
R4990 GND.n4924 GND.n4923 0.125
R4991 GND.n4883 GND.n4882 0.125
R4992 GND.n4843 GND.n4842 0.125
R4993 GND.n4802 GND.n4801 0.125
R4994 GND.n4762 GND.n4761 0.125
R4995 GND.n4721 GND.n4720 0.125
R4996 GND.n4681 GND.n4680 0.125
R4997 GND.n4640 GND.n4639 0.125
R4998 GND.n4600 GND.n4599 0.125
R4999 GND.n5 GND.n4 0.103
R5000 GND.n96 GND.n95 0.103
R5001 GND.n269 GND.n268 0.103
R5002 GND.n606 GND.n605 0.103
R5003 GND.n1926 GND.n1925 0.103
R5004 GND.n4556 GND.n4555 0.103
R5005 GND.n73 GND.n72 0.053
R5006 GND.n82 GND.n81 0.053
R5007 GND.n33 GND.n32 0.053
R5008 GND.n42 GND.n41 0.053
R5009 GND.n245 GND.n244 0.053
R5010 GND.n205 GND.n204 0.053
R5011 GND.n214 GND.n213 0.053
R5012 GND.n164 GND.n163 0.053
R5013 GND.n124 GND.n123 0.053
R5014 GND.n133 GND.n132 0.053
R5015 GND.n580 GND.n579 0.053
R5016 GND.n540 GND.n539 0.053
R5017 GND.n549 GND.n548 0.053
R5018 GND.n499 GND.n498 0.053
R5019 GND.n459 GND.n458 0.053
R5020 GND.n468 GND.n467 0.053
R5021 GND.n418 GND.n417 0.053
R5022 GND.n378 GND.n377 0.053
R5023 GND.n387 GND.n386 0.053
R5024 GND.n337 GND.n336 0.053
R5025 GND.n297 GND.n296 0.053
R5026 GND.n306 GND.n305 0.053
R5027 GND.n1241 GND.n1240 0.053
R5028 GND.n1201 GND.n1200 0.053
R5029 GND.n1210 GND.n1209 0.053
R5030 GND.n1160 GND.n1159 0.053
R5031 GND.n1120 GND.n1119 0.053
R5032 GND.n1129 GND.n1128 0.053
R5033 GND.n1079 GND.n1078 0.053
R5034 GND.n1039 GND.n1038 0.053
R5035 GND.n1048 GND.n1047 0.053
R5036 GND.n998 GND.n997 0.053
R5037 GND.n958 GND.n957 0.053
R5038 GND.n967 GND.n966 0.053
R5039 GND.n917 GND.n916 0.053
R5040 GND.n877 GND.n876 0.053
R5041 GND.n886 GND.n885 0.053
R5042 GND.n836 GND.n835 0.053
R5043 GND.n796 GND.n795 0.053
R5044 GND.n805 GND.n804 0.053
R5045 GND.n755 GND.n754 0.053
R5046 GND.n715 GND.n714 0.053
R5047 GND.n724 GND.n723 0.053
R5048 GND.n674 GND.n673 0.053
R5049 GND.n634 GND.n633 0.053
R5050 GND.n643 GND.n642 0.053
R5051 GND.n1896 GND.n1895 0.053
R5052 GND.n1856 GND.n1855 0.053
R5053 GND.n1865 GND.n1864 0.053
R5054 GND.n1815 GND.n1814 0.053
R5055 GND.n1775 GND.n1774 0.053
R5056 GND.n1784 GND.n1783 0.053
R5057 GND.n1734 GND.n1733 0.053
R5058 GND.n1694 GND.n1693 0.053
R5059 GND.n1703 GND.n1702 0.053
R5060 GND.n1653 GND.n1652 0.053
R5061 GND.n1613 GND.n1612 0.053
R5062 GND.n1622 GND.n1621 0.053
R5063 GND.n1572 GND.n1571 0.053
R5064 GND.n1532 GND.n1531 0.053
R5065 GND.n1541 GND.n1540 0.053
R5066 GND.n1491 GND.n1490 0.053
R5067 GND.n1451 GND.n1450 0.053
R5068 GND.n1460 GND.n1459 0.053
R5069 GND.n1410 GND.n1409 0.053
R5070 GND.n1370 GND.n1369 0.053
R5071 GND.n1379 GND.n1378 0.053
R5072 GND.n1329 GND.n1328 0.053
R5073 GND.n1289 GND.n1288 0.053
R5074 GND.n1298 GND.n1297 0.053
R5075 GND.n2561 GND.n2560 0.053
R5076 GND.n2521 GND.n2520 0.053
R5077 GND.n2530 GND.n2529 0.053
R5078 GND.n2480 GND.n2479 0.053
R5079 GND.n2440 GND.n2439 0.053
R5080 GND.n2449 GND.n2448 0.053
R5081 GND.n2399 GND.n2398 0.053
R5082 GND.n2359 GND.n2358 0.053
R5083 GND.n2368 GND.n2367 0.053
R5084 GND.n2318 GND.n2317 0.053
R5085 GND.n2278 GND.n2277 0.053
R5086 GND.n2287 GND.n2286 0.053
R5087 GND.n2237 GND.n2236 0.053
R5088 GND.n2197 GND.n2196 0.053
R5089 GND.n2206 GND.n2205 0.053
R5090 GND.n2156 GND.n2155 0.053
R5091 GND.n2116 GND.n2115 0.053
R5092 GND.n2125 GND.n2124 0.053
R5093 GND.n2075 GND.n2074 0.053
R5094 GND.n2035 GND.n2034 0.053
R5095 GND.n2044 GND.n2043 0.053
R5096 GND.n1994 GND.n1993 0.053
R5097 GND.n1954 GND.n1953 0.053
R5098 GND.n1963 GND.n1962 0.053
R5099 GND.n3216 GND.n3215 0.053
R5100 GND.n3176 GND.n3175 0.053
R5101 GND.n3185 GND.n3184 0.053
R5102 GND.n3135 GND.n3134 0.053
R5103 GND.n3095 GND.n3094 0.053
R5104 GND.n3104 GND.n3103 0.053
R5105 GND.n3054 GND.n3053 0.053
R5106 GND.n3014 GND.n3013 0.053
R5107 GND.n3023 GND.n3022 0.053
R5108 GND.n2973 GND.n2972 0.053
R5109 GND.n2933 GND.n2932 0.053
R5110 GND.n2942 GND.n2941 0.053
R5111 GND.n2892 GND.n2891 0.053
R5112 GND.n2852 GND.n2851 0.053
R5113 GND.n2861 GND.n2860 0.053
R5114 GND.n2811 GND.n2810 0.053
R5115 GND.n2771 GND.n2770 0.053
R5116 GND.n2780 GND.n2779 0.053
R5117 GND.n2730 GND.n2729 0.053
R5118 GND.n2690 GND.n2689 0.053
R5119 GND.n2699 GND.n2698 0.053
R5120 GND.n2649 GND.n2648 0.053
R5121 GND.n2609 GND.n2608 0.053
R5122 GND.n2618 GND.n2617 0.053
R5123 GND.n3871 GND.n3870 0.053
R5124 GND.n3831 GND.n3830 0.053
R5125 GND.n3840 GND.n3839 0.053
R5126 GND.n3790 GND.n3789 0.053
R5127 GND.n3750 GND.n3749 0.053
R5128 GND.n3759 GND.n3758 0.053
R5129 GND.n3709 GND.n3708 0.053
R5130 GND.n3669 GND.n3668 0.053
R5131 GND.n3678 GND.n3677 0.053
R5132 GND.n3628 GND.n3627 0.053
R5133 GND.n3588 GND.n3587 0.053
R5134 GND.n3597 GND.n3596 0.053
R5135 GND.n3547 GND.n3546 0.053
R5136 GND.n3507 GND.n3506 0.053
R5137 GND.n3516 GND.n3515 0.053
R5138 GND.n3466 GND.n3465 0.053
R5139 GND.n3426 GND.n3425 0.053
R5140 GND.n3435 GND.n3434 0.053
R5141 GND.n3385 GND.n3384 0.053
R5142 GND.n3345 GND.n3344 0.053
R5143 GND.n3354 GND.n3353 0.053
R5144 GND.n3304 GND.n3303 0.053
R5145 GND.n3264 GND.n3263 0.053
R5146 GND.n3273 GND.n3272 0.053
R5147 GND.n4526 GND.n4525 0.053
R5148 GND.n4486 GND.n4485 0.053
R5149 GND.n4495 GND.n4494 0.053
R5150 GND.n4445 GND.n4444 0.053
R5151 GND.n4405 GND.n4404 0.053
R5152 GND.n4414 GND.n4413 0.053
R5153 GND.n4364 GND.n4363 0.053
R5154 GND.n4324 GND.n4323 0.053
R5155 GND.n4333 GND.n4332 0.053
R5156 GND.n4283 GND.n4282 0.053
R5157 GND.n4243 GND.n4242 0.053
R5158 GND.n4252 GND.n4251 0.053
R5159 GND.n4202 GND.n4201 0.053
R5160 GND.n4162 GND.n4161 0.053
R5161 GND.n4171 GND.n4170 0.053
R5162 GND.n4121 GND.n4120 0.053
R5163 GND.n4081 GND.n4080 0.053
R5164 GND.n4090 GND.n4089 0.053
R5165 GND.n4040 GND.n4039 0.053
R5166 GND.n4000 GND.n3999 0.053
R5167 GND.n4009 GND.n4008 0.053
R5168 GND.n3959 GND.n3958 0.053
R5169 GND.n3919 GND.n3918 0.053
R5170 GND.n3928 GND.n3927 0.053
R5171 GND.n5191 GND.n5190 0.053
R5172 GND.n5151 GND.n5150 0.053
R5173 GND.n5160 GND.n5159 0.053
R5174 GND.n5110 GND.n5109 0.053
R5175 GND.n5070 GND.n5069 0.053
R5176 GND.n5079 GND.n5078 0.053
R5177 GND.n5029 GND.n5028 0.053
R5178 GND.n4989 GND.n4988 0.053
R5179 GND.n4998 GND.n4997 0.053
R5180 GND.n4948 GND.n4947 0.053
R5181 GND.n4908 GND.n4907 0.053
R5182 GND.n4917 GND.n4916 0.053
R5183 GND.n4867 GND.n4866 0.053
R5184 GND.n4827 GND.n4826 0.053
R5185 GND.n4836 GND.n4835 0.053
R5186 GND.n4786 GND.n4785 0.053
R5187 GND.n4746 GND.n4745 0.053
R5188 GND.n4755 GND.n4754 0.053
R5189 GND.n4705 GND.n4704 0.053
R5190 GND.n4665 GND.n4664 0.053
R5191 GND.n4674 GND.n4673 0.053
R5192 GND.n4624 GND.n4623 0.053
R5193 GND.n4584 GND.n4583 0.053
R5194 GND.n4593 GND.n4592 0.053
R5195 GND.n6 GND.n5 0.049
R5196 GND.n97 GND.n96 0.049
R5197 GND.n270 GND.n269 0.049
R5198 GND.n607 GND.n606 0.049
R5199 GND.n1927 GND.n1926 0.049
R5200 GND.n4557 GND.n4556 0.049
R5201 GND.n67 GND.n65 0.034
R5202 GND.n88 GND.n86 0.034
R5203 GND.n27 GND.n25 0.034
R5204 GND.n48 GND.n46 0.034
R5205 GND.n239 GND.n237 0.034
R5206 GND.n260 GND.n258 0.034
R5207 GND.n199 GND.n197 0.034
R5208 GND.n220 GND.n218 0.034
R5209 GND.n158 GND.n156 0.034
R5210 GND.n179 GND.n177 0.034
R5211 GND.n118 GND.n116 0.034
R5212 GND.n139 GND.n137 0.034
R5213 GND.n574 GND.n572 0.034
R5214 GND.n595 GND.n593 0.034
R5215 GND.n534 GND.n532 0.034
R5216 GND.n555 GND.n553 0.034
R5217 GND.n493 GND.n491 0.034
R5218 GND.n514 GND.n512 0.034
R5219 GND.n453 GND.n451 0.034
R5220 GND.n474 GND.n472 0.034
R5221 GND.n412 GND.n410 0.034
R5222 GND.n433 GND.n431 0.034
R5223 GND.n372 GND.n370 0.034
R5224 GND.n393 GND.n391 0.034
R5225 GND.n331 GND.n329 0.034
R5226 GND.n352 GND.n350 0.034
R5227 GND.n291 GND.n289 0.034
R5228 GND.n312 GND.n310 0.034
R5229 GND.n1235 GND.n1233 0.034
R5230 GND.n1256 GND.n1254 0.034
R5231 GND.n1195 GND.n1193 0.034
R5232 GND.n1216 GND.n1214 0.034
R5233 GND.n1154 GND.n1152 0.034
R5234 GND.n1175 GND.n1173 0.034
R5235 GND.n1114 GND.n1112 0.034
R5236 GND.n1135 GND.n1133 0.034
R5237 GND.n1073 GND.n1071 0.034
R5238 GND.n1094 GND.n1092 0.034
R5239 GND.n1033 GND.n1031 0.034
R5240 GND.n1054 GND.n1052 0.034
R5241 GND.n992 GND.n990 0.034
R5242 GND.n1013 GND.n1011 0.034
R5243 GND.n952 GND.n950 0.034
R5244 GND.n973 GND.n971 0.034
R5245 GND.n911 GND.n909 0.034
R5246 GND.n932 GND.n930 0.034
R5247 GND.n871 GND.n869 0.034
R5248 GND.n892 GND.n890 0.034
R5249 GND.n830 GND.n828 0.034
R5250 GND.n851 GND.n849 0.034
R5251 GND.n790 GND.n788 0.034
R5252 GND.n811 GND.n809 0.034
R5253 GND.n749 GND.n747 0.034
R5254 GND.n770 GND.n768 0.034
R5255 GND.n709 GND.n707 0.034
R5256 GND.n730 GND.n728 0.034
R5257 GND.n668 GND.n666 0.034
R5258 GND.n689 GND.n687 0.034
R5259 GND.n628 GND.n626 0.034
R5260 GND.n649 GND.n647 0.034
R5261 GND.n1890 GND.n1888 0.034
R5262 GND.n1911 GND.n1909 0.034
R5263 GND.n1850 GND.n1848 0.034
R5264 GND.n1871 GND.n1869 0.034
R5265 GND.n1809 GND.n1807 0.034
R5266 GND.n1830 GND.n1828 0.034
R5267 GND.n1769 GND.n1767 0.034
R5268 GND.n1790 GND.n1788 0.034
R5269 GND.n1728 GND.n1726 0.034
R5270 GND.n1749 GND.n1747 0.034
R5271 GND.n1688 GND.n1686 0.034
R5272 GND.n1709 GND.n1707 0.034
R5273 GND.n1647 GND.n1645 0.034
R5274 GND.n1668 GND.n1666 0.034
R5275 GND.n1607 GND.n1605 0.034
R5276 GND.n1628 GND.n1626 0.034
R5277 GND.n1566 GND.n1564 0.034
R5278 GND.n1587 GND.n1585 0.034
R5279 GND.n1526 GND.n1524 0.034
R5280 GND.n1547 GND.n1545 0.034
R5281 GND.n1485 GND.n1483 0.034
R5282 GND.n1506 GND.n1504 0.034
R5283 GND.n1445 GND.n1443 0.034
R5284 GND.n1466 GND.n1464 0.034
R5285 GND.n1404 GND.n1402 0.034
R5286 GND.n1425 GND.n1423 0.034
R5287 GND.n1364 GND.n1362 0.034
R5288 GND.n1385 GND.n1383 0.034
R5289 GND.n1323 GND.n1321 0.034
R5290 GND.n1344 GND.n1342 0.034
R5291 GND.n1283 GND.n1281 0.034
R5292 GND.n1304 GND.n1302 0.034
R5293 GND.n2555 GND.n2553 0.034
R5294 GND.n2576 GND.n2574 0.034
R5295 GND.n2515 GND.n2513 0.034
R5296 GND.n2536 GND.n2534 0.034
R5297 GND.n2474 GND.n2472 0.034
R5298 GND.n2495 GND.n2493 0.034
R5299 GND.n2434 GND.n2432 0.034
R5300 GND.n2455 GND.n2453 0.034
R5301 GND.n2393 GND.n2391 0.034
R5302 GND.n2414 GND.n2412 0.034
R5303 GND.n2353 GND.n2351 0.034
R5304 GND.n2374 GND.n2372 0.034
R5305 GND.n2312 GND.n2310 0.034
R5306 GND.n2333 GND.n2331 0.034
R5307 GND.n2272 GND.n2270 0.034
R5308 GND.n2293 GND.n2291 0.034
R5309 GND.n2231 GND.n2229 0.034
R5310 GND.n2252 GND.n2250 0.034
R5311 GND.n2191 GND.n2189 0.034
R5312 GND.n2212 GND.n2210 0.034
R5313 GND.n2150 GND.n2148 0.034
R5314 GND.n2171 GND.n2169 0.034
R5315 GND.n2110 GND.n2108 0.034
R5316 GND.n2131 GND.n2129 0.034
R5317 GND.n2069 GND.n2067 0.034
R5318 GND.n2090 GND.n2088 0.034
R5319 GND.n2029 GND.n2027 0.034
R5320 GND.n2050 GND.n2048 0.034
R5321 GND.n1988 GND.n1986 0.034
R5322 GND.n2009 GND.n2007 0.034
R5323 GND.n1948 GND.n1946 0.034
R5324 GND.n1969 GND.n1967 0.034
R5325 GND.n3210 GND.n3208 0.034
R5326 GND.n3231 GND.n3229 0.034
R5327 GND.n3170 GND.n3168 0.034
R5328 GND.n3191 GND.n3189 0.034
R5329 GND.n3129 GND.n3127 0.034
R5330 GND.n3150 GND.n3148 0.034
R5331 GND.n3089 GND.n3087 0.034
R5332 GND.n3110 GND.n3108 0.034
R5333 GND.n3048 GND.n3046 0.034
R5334 GND.n3069 GND.n3067 0.034
R5335 GND.n3008 GND.n3006 0.034
R5336 GND.n3029 GND.n3027 0.034
R5337 GND.n2967 GND.n2965 0.034
R5338 GND.n2988 GND.n2986 0.034
R5339 GND.n2927 GND.n2925 0.034
R5340 GND.n2948 GND.n2946 0.034
R5341 GND.n2886 GND.n2884 0.034
R5342 GND.n2907 GND.n2905 0.034
R5343 GND.n2846 GND.n2844 0.034
R5344 GND.n2867 GND.n2865 0.034
R5345 GND.n2805 GND.n2803 0.034
R5346 GND.n2826 GND.n2824 0.034
R5347 GND.n2765 GND.n2763 0.034
R5348 GND.n2786 GND.n2784 0.034
R5349 GND.n2724 GND.n2722 0.034
R5350 GND.n2745 GND.n2743 0.034
R5351 GND.n2684 GND.n2682 0.034
R5352 GND.n2705 GND.n2703 0.034
R5353 GND.n2643 GND.n2641 0.034
R5354 GND.n2664 GND.n2662 0.034
R5355 GND.n2603 GND.n2601 0.034
R5356 GND.n2624 GND.n2622 0.034
R5357 GND.n3865 GND.n3863 0.034
R5358 GND.n3886 GND.n3884 0.034
R5359 GND.n3825 GND.n3823 0.034
R5360 GND.n3846 GND.n3844 0.034
R5361 GND.n3784 GND.n3782 0.034
R5362 GND.n3805 GND.n3803 0.034
R5363 GND.n3744 GND.n3742 0.034
R5364 GND.n3765 GND.n3763 0.034
R5365 GND.n3703 GND.n3701 0.034
R5366 GND.n3724 GND.n3722 0.034
R5367 GND.n3663 GND.n3661 0.034
R5368 GND.n3684 GND.n3682 0.034
R5369 GND.n3622 GND.n3620 0.034
R5370 GND.n3643 GND.n3641 0.034
R5371 GND.n3582 GND.n3580 0.034
R5372 GND.n3603 GND.n3601 0.034
R5373 GND.n3541 GND.n3539 0.034
R5374 GND.n3562 GND.n3560 0.034
R5375 GND.n3501 GND.n3499 0.034
R5376 GND.n3522 GND.n3520 0.034
R5377 GND.n3460 GND.n3458 0.034
R5378 GND.n3481 GND.n3479 0.034
R5379 GND.n3420 GND.n3418 0.034
R5380 GND.n3441 GND.n3439 0.034
R5381 GND.n3379 GND.n3377 0.034
R5382 GND.n3400 GND.n3398 0.034
R5383 GND.n3339 GND.n3337 0.034
R5384 GND.n3360 GND.n3358 0.034
R5385 GND.n3298 GND.n3296 0.034
R5386 GND.n3319 GND.n3317 0.034
R5387 GND.n3258 GND.n3256 0.034
R5388 GND.n3279 GND.n3277 0.034
R5389 GND.n4520 GND.n4518 0.034
R5390 GND.n4541 GND.n4539 0.034
R5391 GND.n4480 GND.n4478 0.034
R5392 GND.n4501 GND.n4499 0.034
R5393 GND.n4439 GND.n4437 0.034
R5394 GND.n4460 GND.n4458 0.034
R5395 GND.n4399 GND.n4397 0.034
R5396 GND.n4420 GND.n4418 0.034
R5397 GND.n4358 GND.n4356 0.034
R5398 GND.n4379 GND.n4377 0.034
R5399 GND.n4318 GND.n4316 0.034
R5400 GND.n4339 GND.n4337 0.034
R5401 GND.n4277 GND.n4275 0.034
R5402 GND.n4298 GND.n4296 0.034
R5403 GND.n4237 GND.n4235 0.034
R5404 GND.n4258 GND.n4256 0.034
R5405 GND.n4196 GND.n4194 0.034
R5406 GND.n4217 GND.n4215 0.034
R5407 GND.n4156 GND.n4154 0.034
R5408 GND.n4177 GND.n4175 0.034
R5409 GND.n4115 GND.n4113 0.034
R5410 GND.n4136 GND.n4134 0.034
R5411 GND.n4075 GND.n4073 0.034
R5412 GND.n4096 GND.n4094 0.034
R5413 GND.n4034 GND.n4032 0.034
R5414 GND.n4055 GND.n4053 0.034
R5415 GND.n3994 GND.n3992 0.034
R5416 GND.n4015 GND.n4013 0.034
R5417 GND.n3953 GND.n3951 0.034
R5418 GND.n3974 GND.n3972 0.034
R5419 GND.n3913 GND.n3911 0.034
R5420 GND.n3934 GND.n3932 0.034
R5421 GND.n5185 GND.n5183 0.034
R5422 GND.n5206 GND.n5204 0.034
R5423 GND.n5145 GND.n5143 0.034
R5424 GND.n5166 GND.n5164 0.034
R5425 GND.n5104 GND.n5102 0.034
R5426 GND.n5125 GND.n5123 0.034
R5427 GND.n5064 GND.n5062 0.034
R5428 GND.n5085 GND.n5083 0.034
R5429 GND.n5023 GND.n5021 0.034
R5430 GND.n5044 GND.n5042 0.034
R5431 GND.n4983 GND.n4981 0.034
R5432 GND.n5004 GND.n5002 0.034
R5433 GND.n4942 GND.n4940 0.034
R5434 GND.n4963 GND.n4961 0.034
R5435 GND.n4902 GND.n4900 0.034
R5436 GND.n4923 GND.n4921 0.034
R5437 GND.n4861 GND.n4859 0.034
R5438 GND.n4882 GND.n4880 0.034
R5439 GND.n4821 GND.n4819 0.034
R5440 GND.n4842 GND.n4840 0.034
R5441 GND.n4780 GND.n4778 0.034
R5442 GND.n4801 GND.n4799 0.034
R5443 GND.n4740 GND.n4738 0.034
R5444 GND.n4761 GND.n4759 0.034
R5445 GND.n4699 GND.n4697 0.034
R5446 GND.n4720 GND.n4718 0.034
R5447 GND.n4659 GND.n4657 0.034
R5448 GND.n4680 GND.n4678 0.034
R5449 GND.n4618 GND.n4616 0.034
R5450 GND.n4639 GND.n4637 0.034
R5451 GND.n4578 GND.n4576 0.034
R5452 GND.n4599 GND.n4597 0.034
R5453 GND.n100 GND.n99 0.011
R5454 GND.n273 GND.n272 0.011
R5455 GND.n610 GND.n609 0.011
R5456 GND.n1930 GND.n1929 0.011
R5457 GND.n4560 GND.n4559 0.011
R5458 GND.n9 GND.n8 0.011
R5459 GND.n100 GND.n98 0.011
R5460 GND.n273 GND.n271 0.011
R5461 GND.n610 GND.n608 0.011
R5462 GND.n1930 GND.n1928 0.011
R5463 GND.n4560 GND.n4558 0.011
R5464 GND.n9 GND.n7 0.011
R5465 GND.n7 GND.n6 0.003
R5466 GND.n98 GND.n97 0.003
R5467 GND.n271 GND.n270 0.003
R5468 GND.n608 GND.n607 0.003
R5469 GND.n1928 GND.n1927 0.003
R5470 GND.n4558 GND.n4557 0.003
R5471 GND.n75 GND.n67 0.002
R5472 GND.n86 GND.n84 0.002
R5473 GND.n35 GND.n27 0.002
R5474 GND.n46 GND.n44 0.002
R5475 GND.n247 GND.n239 0.002
R5476 GND.n258 GND.n256 0.002
R5477 GND.n207 GND.n199 0.002
R5478 GND.n218 GND.n216 0.002
R5479 GND.n166 GND.n158 0.002
R5480 GND.n177 GND.n175 0.002
R5481 GND.n126 GND.n118 0.002
R5482 GND.n137 GND.n135 0.002
R5483 GND.n582 GND.n574 0.002
R5484 GND.n593 GND.n591 0.002
R5485 GND.n542 GND.n534 0.002
R5486 GND.n553 GND.n551 0.002
R5487 GND.n501 GND.n493 0.002
R5488 GND.n512 GND.n510 0.002
R5489 GND.n461 GND.n453 0.002
R5490 GND.n472 GND.n470 0.002
R5491 GND.n420 GND.n412 0.002
R5492 GND.n431 GND.n429 0.002
R5493 GND.n380 GND.n372 0.002
R5494 GND.n391 GND.n389 0.002
R5495 GND.n339 GND.n331 0.002
R5496 GND.n350 GND.n348 0.002
R5497 GND.n299 GND.n291 0.002
R5498 GND.n310 GND.n308 0.002
R5499 GND.n1243 GND.n1235 0.002
R5500 GND.n1254 GND.n1252 0.002
R5501 GND.n1203 GND.n1195 0.002
R5502 GND.n1214 GND.n1212 0.002
R5503 GND.n1162 GND.n1154 0.002
R5504 GND.n1173 GND.n1171 0.002
R5505 GND.n1122 GND.n1114 0.002
R5506 GND.n1133 GND.n1131 0.002
R5507 GND.n1081 GND.n1073 0.002
R5508 GND.n1092 GND.n1090 0.002
R5509 GND.n1041 GND.n1033 0.002
R5510 GND.n1052 GND.n1050 0.002
R5511 GND.n1000 GND.n992 0.002
R5512 GND.n1011 GND.n1009 0.002
R5513 GND.n960 GND.n952 0.002
R5514 GND.n971 GND.n969 0.002
R5515 GND.n919 GND.n911 0.002
R5516 GND.n930 GND.n928 0.002
R5517 GND.n879 GND.n871 0.002
R5518 GND.n890 GND.n888 0.002
R5519 GND.n838 GND.n830 0.002
R5520 GND.n849 GND.n847 0.002
R5521 GND.n798 GND.n790 0.002
R5522 GND.n809 GND.n807 0.002
R5523 GND.n757 GND.n749 0.002
R5524 GND.n768 GND.n766 0.002
R5525 GND.n717 GND.n709 0.002
R5526 GND.n728 GND.n726 0.002
R5527 GND.n676 GND.n668 0.002
R5528 GND.n687 GND.n685 0.002
R5529 GND.n636 GND.n628 0.002
R5530 GND.n647 GND.n645 0.002
R5531 GND.n1898 GND.n1890 0.002
R5532 GND.n1909 GND.n1907 0.002
R5533 GND.n1858 GND.n1850 0.002
R5534 GND.n1869 GND.n1867 0.002
R5535 GND.n1817 GND.n1809 0.002
R5536 GND.n1828 GND.n1826 0.002
R5537 GND.n1777 GND.n1769 0.002
R5538 GND.n1788 GND.n1786 0.002
R5539 GND.n1736 GND.n1728 0.002
R5540 GND.n1747 GND.n1745 0.002
R5541 GND.n1696 GND.n1688 0.002
R5542 GND.n1707 GND.n1705 0.002
R5543 GND.n1655 GND.n1647 0.002
R5544 GND.n1666 GND.n1664 0.002
R5545 GND.n1615 GND.n1607 0.002
R5546 GND.n1626 GND.n1624 0.002
R5547 GND.n1574 GND.n1566 0.002
R5548 GND.n1585 GND.n1583 0.002
R5549 GND.n1534 GND.n1526 0.002
R5550 GND.n1545 GND.n1543 0.002
R5551 GND.n1493 GND.n1485 0.002
R5552 GND.n1504 GND.n1502 0.002
R5553 GND.n1453 GND.n1445 0.002
R5554 GND.n1464 GND.n1462 0.002
R5555 GND.n1412 GND.n1404 0.002
R5556 GND.n1423 GND.n1421 0.002
R5557 GND.n1372 GND.n1364 0.002
R5558 GND.n1383 GND.n1381 0.002
R5559 GND.n1331 GND.n1323 0.002
R5560 GND.n1342 GND.n1340 0.002
R5561 GND.n1291 GND.n1283 0.002
R5562 GND.n1302 GND.n1300 0.002
R5563 GND.n2563 GND.n2555 0.002
R5564 GND.n2574 GND.n2572 0.002
R5565 GND.n2523 GND.n2515 0.002
R5566 GND.n2534 GND.n2532 0.002
R5567 GND.n2482 GND.n2474 0.002
R5568 GND.n2493 GND.n2491 0.002
R5569 GND.n2442 GND.n2434 0.002
R5570 GND.n2453 GND.n2451 0.002
R5571 GND.n2401 GND.n2393 0.002
R5572 GND.n2412 GND.n2410 0.002
R5573 GND.n2361 GND.n2353 0.002
R5574 GND.n2372 GND.n2370 0.002
R5575 GND.n2320 GND.n2312 0.002
R5576 GND.n2331 GND.n2329 0.002
R5577 GND.n2280 GND.n2272 0.002
R5578 GND.n2291 GND.n2289 0.002
R5579 GND.n2239 GND.n2231 0.002
R5580 GND.n2250 GND.n2248 0.002
R5581 GND.n2199 GND.n2191 0.002
R5582 GND.n2210 GND.n2208 0.002
R5583 GND.n2158 GND.n2150 0.002
R5584 GND.n2169 GND.n2167 0.002
R5585 GND.n2118 GND.n2110 0.002
R5586 GND.n2129 GND.n2127 0.002
R5587 GND.n2077 GND.n2069 0.002
R5588 GND.n2088 GND.n2086 0.002
R5589 GND.n2037 GND.n2029 0.002
R5590 GND.n2048 GND.n2046 0.002
R5591 GND.n1996 GND.n1988 0.002
R5592 GND.n2007 GND.n2005 0.002
R5593 GND.n1956 GND.n1948 0.002
R5594 GND.n1967 GND.n1965 0.002
R5595 GND.n3218 GND.n3210 0.002
R5596 GND.n3229 GND.n3227 0.002
R5597 GND.n3178 GND.n3170 0.002
R5598 GND.n3189 GND.n3187 0.002
R5599 GND.n3137 GND.n3129 0.002
R5600 GND.n3148 GND.n3146 0.002
R5601 GND.n3097 GND.n3089 0.002
R5602 GND.n3108 GND.n3106 0.002
R5603 GND.n3056 GND.n3048 0.002
R5604 GND.n3067 GND.n3065 0.002
R5605 GND.n3016 GND.n3008 0.002
R5606 GND.n3027 GND.n3025 0.002
R5607 GND.n2975 GND.n2967 0.002
R5608 GND.n2986 GND.n2984 0.002
R5609 GND.n2935 GND.n2927 0.002
R5610 GND.n2946 GND.n2944 0.002
R5611 GND.n2894 GND.n2886 0.002
R5612 GND.n2905 GND.n2903 0.002
R5613 GND.n2854 GND.n2846 0.002
R5614 GND.n2865 GND.n2863 0.002
R5615 GND.n2813 GND.n2805 0.002
R5616 GND.n2824 GND.n2822 0.002
R5617 GND.n2773 GND.n2765 0.002
R5618 GND.n2784 GND.n2782 0.002
R5619 GND.n2732 GND.n2724 0.002
R5620 GND.n2743 GND.n2741 0.002
R5621 GND.n2692 GND.n2684 0.002
R5622 GND.n2703 GND.n2701 0.002
R5623 GND.n2651 GND.n2643 0.002
R5624 GND.n2662 GND.n2660 0.002
R5625 GND.n2611 GND.n2603 0.002
R5626 GND.n2622 GND.n2620 0.002
R5627 GND.n3873 GND.n3865 0.002
R5628 GND.n3884 GND.n3882 0.002
R5629 GND.n3833 GND.n3825 0.002
R5630 GND.n3844 GND.n3842 0.002
R5631 GND.n3792 GND.n3784 0.002
R5632 GND.n3803 GND.n3801 0.002
R5633 GND.n3752 GND.n3744 0.002
R5634 GND.n3763 GND.n3761 0.002
R5635 GND.n3711 GND.n3703 0.002
R5636 GND.n3722 GND.n3720 0.002
R5637 GND.n3671 GND.n3663 0.002
R5638 GND.n3682 GND.n3680 0.002
R5639 GND.n3630 GND.n3622 0.002
R5640 GND.n3641 GND.n3639 0.002
R5641 GND.n3590 GND.n3582 0.002
R5642 GND.n3601 GND.n3599 0.002
R5643 GND.n3549 GND.n3541 0.002
R5644 GND.n3560 GND.n3558 0.002
R5645 GND.n3509 GND.n3501 0.002
R5646 GND.n3520 GND.n3518 0.002
R5647 GND.n3468 GND.n3460 0.002
R5648 GND.n3479 GND.n3477 0.002
R5649 GND.n3428 GND.n3420 0.002
R5650 GND.n3439 GND.n3437 0.002
R5651 GND.n3387 GND.n3379 0.002
R5652 GND.n3398 GND.n3396 0.002
R5653 GND.n3347 GND.n3339 0.002
R5654 GND.n3358 GND.n3356 0.002
R5655 GND.n3306 GND.n3298 0.002
R5656 GND.n3317 GND.n3315 0.002
R5657 GND.n3266 GND.n3258 0.002
R5658 GND.n3277 GND.n3275 0.002
R5659 GND.n4528 GND.n4520 0.002
R5660 GND.n4539 GND.n4537 0.002
R5661 GND.n4488 GND.n4480 0.002
R5662 GND.n4499 GND.n4497 0.002
R5663 GND.n4447 GND.n4439 0.002
R5664 GND.n4458 GND.n4456 0.002
R5665 GND.n4407 GND.n4399 0.002
R5666 GND.n4418 GND.n4416 0.002
R5667 GND.n4366 GND.n4358 0.002
R5668 GND.n4377 GND.n4375 0.002
R5669 GND.n4326 GND.n4318 0.002
R5670 GND.n4337 GND.n4335 0.002
R5671 GND.n4285 GND.n4277 0.002
R5672 GND.n4296 GND.n4294 0.002
R5673 GND.n4245 GND.n4237 0.002
R5674 GND.n4256 GND.n4254 0.002
R5675 GND.n4204 GND.n4196 0.002
R5676 GND.n4215 GND.n4213 0.002
R5677 GND.n4164 GND.n4156 0.002
R5678 GND.n4175 GND.n4173 0.002
R5679 GND.n4123 GND.n4115 0.002
R5680 GND.n4134 GND.n4132 0.002
R5681 GND.n4083 GND.n4075 0.002
R5682 GND.n4094 GND.n4092 0.002
R5683 GND.n4042 GND.n4034 0.002
R5684 GND.n4053 GND.n4051 0.002
R5685 GND.n4002 GND.n3994 0.002
R5686 GND.n4013 GND.n4011 0.002
R5687 GND.n3961 GND.n3953 0.002
R5688 GND.n3972 GND.n3970 0.002
R5689 GND.n3921 GND.n3913 0.002
R5690 GND.n3932 GND.n3930 0.002
R5691 GND.n5193 GND.n5185 0.002
R5692 GND.n5204 GND.n5202 0.002
R5693 GND.n5153 GND.n5145 0.002
R5694 GND.n5164 GND.n5162 0.002
R5695 GND.n5112 GND.n5104 0.002
R5696 GND.n5123 GND.n5121 0.002
R5697 GND.n5072 GND.n5064 0.002
R5698 GND.n5083 GND.n5081 0.002
R5699 GND.n5031 GND.n5023 0.002
R5700 GND.n5042 GND.n5040 0.002
R5701 GND.n4991 GND.n4983 0.002
R5702 GND.n5002 GND.n5000 0.002
R5703 GND.n4950 GND.n4942 0.002
R5704 GND.n4961 GND.n4959 0.002
R5705 GND.n4910 GND.n4902 0.002
R5706 GND.n4921 GND.n4919 0.002
R5707 GND.n4869 GND.n4861 0.002
R5708 GND.n4880 GND.n4878 0.002
R5709 GND.n4829 GND.n4821 0.002
R5710 GND.n4840 GND.n4838 0.002
R5711 GND.n4788 GND.n4780 0.002
R5712 GND.n4799 GND.n4797 0.002
R5713 GND.n4748 GND.n4740 0.002
R5714 GND.n4759 GND.n4757 0.002
R5715 GND.n4707 GND.n4699 0.002
R5716 GND.n4718 GND.n4716 0.002
R5717 GND.n4667 GND.n4659 0.002
R5718 GND.n4678 GND.n4676 0.002
R5719 GND.n4626 GND.n4618 0.002
R5720 GND.n4637 GND.n4635 0.002
R5721 GND.n4586 GND.n4578 0.002
R5722 GND.n4597 GND.n4595 0.002
R5723 OUT_P.n55 OUT_P.n54 1.088
R5724 OUT_P.n57 OUT_P.n36 0.872
R5725 OUT_P.n56 OUT_P.n42 0.872
R5726 OUT_P.n55 OUT_P.n48 0.872
R5727 OUT_P.n59 OUT_P.n23 0.64
R5728 OUT_P.n58 OUT_P.n30 0.64
R5729 OUT_P.n0 OUT_P.t48 0.474
R5730 OUT_P.n9 OUT_P.t36 0.474
R5731 OUT_P.n17 OUT_P.t37 0.474
R5732 OUT_P.n24 OUT_P.t42 0.474
R5733 OUT_P.n31 OUT_P.t17 0.474
R5734 OUT_P.n37 OUT_P.t10 0.474
R5735 OUT_P.n43 OUT_P.t13 0.474
R5736 OUT_P.n60 OUT_P.n16 0.408
R5737 OUT_P.n49 OUT_P.t20 0.36
R5738 OUT_P OUT_P.n61 0.276
R5739 OUT_P.n6 OUT_P.t52 0.242
R5740 OUT_P.n5 OUT_P.t26 0.242
R5741 OUT_P.n4 OUT_P.t1 0.242
R5742 OUT_P.n3 OUT_P.t40 0.242
R5743 OUT_P.n2 OUT_P.t15 0.242
R5744 OUT_P.n1 OUT_P.t58 0.242
R5745 OUT_P.n0 OUT_P.t32 0.242
R5746 OUT_P.n14 OUT_P.t6 0.242
R5747 OUT_P.n13 OUT_P.t46 0.242
R5748 OUT_P.n12 OUT_P.t21 0.242
R5749 OUT_P.n11 OUT_P.t57 0.242
R5750 OUT_P.n10 OUT_P.t35 0.242
R5751 OUT_P.n9 OUT_P.t8 0.242
R5752 OUT_P.n22 OUT_P.t30 0.242
R5753 OUT_P.n21 OUT_P.t5 0.242
R5754 OUT_P.n20 OUT_P.t45 0.242
R5755 OUT_P.n19 OUT_P.t18 0.242
R5756 OUT_P.n18 OUT_P.t61 0.242
R5757 OUT_P.n17 OUT_P.t34 0.242
R5758 OUT_P.n28 OUT_P.t29 0.242
R5759 OUT_P.n27 OUT_P.t4 0.242
R5760 OUT_P.n26 OUT_P.t43 0.242
R5761 OUT_P.n25 OUT_P.t23 0.242
R5762 OUT_P.n24 OUT_P.t60 0.242
R5763 OUT_P.n35 OUT_P.t12 0.242
R5764 OUT_P.n34 OUT_P.t53 0.242
R5765 OUT_P.n33 OUT_P.t27 0.242
R5766 OUT_P.n32 OUT_P.t7 0.242
R5767 OUT_P.n31 OUT_P.t47 0.242
R5768 OUT_P.n41 OUT_P.t3 0.242
R5769 OUT_P.n40 OUT_P.t41 0.242
R5770 OUT_P.n39 OUT_P.t16 0.242
R5771 OUT_P.n38 OUT_P.t59 0.242
R5772 OUT_P.n37 OUT_P.t33 0.242
R5773 OUT_P.n47 OUT_P.t25 0.242
R5774 OUT_P.n46 OUT_P.t0 0.242
R5775 OUT_P.n45 OUT_P.t39 0.242
R5776 OUT_P.n44 OUT_P.t22 0.242
R5777 OUT_P.n43 OUT_P.t56 0.242
R5778 OUT_P.n8 OUT_P.n7 0.232
R5779 OUT_P.n7 OUT_P.n6 0.232
R5780 OUT_P.n6 OUT_P.n5 0.232
R5781 OUT_P.n5 OUT_P.n4 0.232
R5782 OUT_P.n4 OUT_P.n3 0.232
R5783 OUT_P.n3 OUT_P.n2 0.232
R5784 OUT_P.n2 OUT_P.n1 0.232
R5785 OUT_P.n1 OUT_P.n0 0.232
R5786 OUT_P.n16 OUT_P.n15 0.232
R5787 OUT_P.n15 OUT_P.n14 0.232
R5788 OUT_P.n14 OUT_P.n13 0.232
R5789 OUT_P.n13 OUT_P.n12 0.232
R5790 OUT_P.n12 OUT_P.n11 0.232
R5791 OUT_P.n11 OUT_P.n10 0.232
R5792 OUT_P.n10 OUT_P.n9 0.232
R5793 OUT_P.n23 OUT_P.n22 0.232
R5794 OUT_P.n22 OUT_P.n21 0.232
R5795 OUT_P.n21 OUT_P.n20 0.232
R5796 OUT_P.n20 OUT_P.n19 0.232
R5797 OUT_P.n19 OUT_P.n18 0.232
R5798 OUT_P.n18 OUT_P.n17 0.232
R5799 OUT_P.n30 OUT_P.n29 0.232
R5800 OUT_P.n29 OUT_P.n28 0.232
R5801 OUT_P.n28 OUT_P.n27 0.232
R5802 OUT_P.n27 OUT_P.n26 0.232
R5803 OUT_P.n26 OUT_P.n25 0.232
R5804 OUT_P.n25 OUT_P.n24 0.232
R5805 OUT_P.n36 OUT_P.n35 0.232
R5806 OUT_P.n35 OUT_P.n34 0.232
R5807 OUT_P.n34 OUT_P.n33 0.232
R5808 OUT_P.n33 OUT_P.n32 0.232
R5809 OUT_P.n32 OUT_P.n31 0.232
R5810 OUT_P.n42 OUT_P.n41 0.232
R5811 OUT_P.n41 OUT_P.n40 0.232
R5812 OUT_P.n40 OUT_P.n39 0.232
R5813 OUT_P.n39 OUT_P.n38 0.232
R5814 OUT_P.n38 OUT_P.n37 0.232
R5815 OUT_P.n48 OUT_P.n47 0.232
R5816 OUT_P.n47 OUT_P.n46 0.232
R5817 OUT_P.n46 OUT_P.n45 0.232
R5818 OUT_P.n45 OUT_P.n44 0.232
R5819 OUT_P.n44 OUT_P.n43 0.232
R5820 OUT_P.n54 OUT_P.n53 0.232
R5821 OUT_P.n53 OUT_P.n52 0.232
R5822 OUT_P.n52 OUT_P.n51 0.232
R5823 OUT_P.n51 OUT_P.n50 0.232
R5824 OUT_P.n50 OUT_P.n49 0.232
R5825 OUT_P.n56 OUT_P.n55 0.216
R5826 OUT_P.n57 OUT_P.n56 0.216
R5827 OUT_P.n58 OUT_P.n57 0.216
R5828 OUT_P.n59 OUT_P.n58 0.216
R5829 OUT_P.n60 OUT_P.n59 0.216
R5830 OUT_P.n61 OUT_P.n60 0.216
R5831 OUT_P.n61 OUT_P.n8 0.176
R5832 OUT_P.n8 OUT_P.t2 0.128
R5833 OUT_P.n7 OUT_P.t9 0.128
R5834 OUT_P.n16 OUT_P.t51 0.128
R5835 OUT_P.n15 OUT_P.t31 0.128
R5836 OUT_P.n23 OUT_P.t55 0.128
R5837 OUT_P.n30 OUT_P.t14 0.128
R5838 OUT_P.n29 OUT_P.t54 0.128
R5839 OUT_P.n36 OUT_P.t38 0.128
R5840 OUT_P.n42 OUT_P.t28 0.128
R5841 OUT_P.n48 OUT_P.t50 0.128
R5842 OUT_P.n54 OUT_P.t11 0.128
R5843 OUT_P.n53 OUT_P.t49 0.128
R5844 OUT_P.n52 OUT_P.t24 0.128
R5845 OUT_P.n51 OUT_P.t62 0.128
R5846 OUT_P.n50 OUT_P.t44 0.128
R5847 OUT_P.n49 OUT_P.t19 0.128
R5848 a_59376_45486.n10 a_59376_45486.t1 10.181
R5849 a_59376_45486.n10 a_59376_45486.t0 10.181
R5850 a_59376_45486.t3 a_59376_45486.n18 9.68
R5851 a_59376_45486.n1 a_59376_45486.n0 9.302
R5852 a_59376_45486.n7 a_59376_45486.n6 9.3
R5853 a_59376_45486.n5 a_59376_45486.n4 9.3
R5854 a_59376_45486.n9 a_59376_45486.n8 9
R5855 a_59376_45486.n13 a_59376_45486.n12 7.729
R5856 a_59376_45486.n13 a_59376_45486.n10 6.296
R5857 a_59376_45486.n16 a_59376_45486.n1 4.508
R5858 a_59376_45486.n15 a_59376_45486.n14 4.501
R5859 a_59376_45486.n15 a_59376_45486.n9 4.501
R5860 a_59376_45486.n16 a_59376_45486.n3 4.494
R5861 a_59376_45486.n18 a_59376_45486.t2 1.259
R5862 a_59376_45486.n12 a_59376_45486.n11 0.536
R5863 a_59376_45486.n18 a_59376_45486.n17 0.415
R5864 a_59376_45486.n14 a_59376_45486.n13 0.151
R5865 a_59376_45486.n7 a_59376_45486.n5 0.028
R5866 a_59376_45486.n3 a_59376_45486.n2 0.025
R5867 a_59376_45486.n17 a_59376_45486.n16 0.021
R5868 a_59376_45486.n9 a_59376_45486.n7 0.012
R5869 a_59376_45486.n16 a_59376_45486.n15 0.006
R5870 bit5.n247 bit5.t65 552.693
R5871 bit5.n2 bit5.t5 300.446
R5872 bit5.n0 bit5.t43 300.446
R5873 bit5.n9 bit5.t12 300.446
R5874 bit5.n7 bit5.t40 300.446
R5875 bit5.n16 bit5.t37 300.446
R5876 bit5.n14 bit5.t61 300.446
R5877 bit5.n23 bit5.t33 300.446
R5878 bit5.n21 bit5.t59 300.446
R5879 bit5.n30 bit5.t28 300.446
R5880 bit5.n28 bit5.t55 300.446
R5881 bit5.n37 bit5.t24 300.446
R5882 bit5.n35 bit5.t60 300.446
R5883 bit5.n44 bit5.t31 300.446
R5884 bit5.n42 bit5.t58 300.446
R5885 bit5.n53 bit5.t46 300.446
R5886 bit5.n51 bit5.t3 300.446
R5887 bit5.n65 bit5.t52 300.446
R5888 bit5.n63 bit5.t18 300.446
R5889 bit5.n72 bit5.t53 300.446
R5890 bit5.n70 bit5.t16 300.446
R5891 bit5.n79 bit5.t15 300.446
R5892 bit5.n77 bit5.t42 300.446
R5893 bit5.n86 bit5.t11 300.446
R5894 bit5.n84 bit5.t39 300.446
R5895 bit5.n93 bit5.t8 300.446
R5896 bit5.n91 bit5.t35 300.446
R5897 bit5.n100 bit5.t4 300.446
R5898 bit5.n98 bit5.t41 300.446
R5899 bit5.n107 bit5.t10 300.446
R5900 bit5.n105 bit5.t36 300.446
R5901 bit5.n114 bit5.t21 300.446
R5902 bit5.n112 bit5.t50 300.446
R5903 bit5.n129 bit5.t45 300.446
R5904 bit5.n127 bit5.t13 300.446
R5905 bit5.n136 bit5.t49 300.446
R5906 bit5.n134 bit5.t9 300.446
R5907 bit5.n143 bit5.t6 300.446
R5908 bit5.n141 bit5.t34 300.446
R5909 bit5.n150 bit5.t2 300.446
R5910 bit5.n148 bit5.t29 300.446
R5911 bit5.n157 bit5.t64 300.446
R5912 bit5.n155 bit5.t25 300.446
R5913 bit5.n164 bit5.t63 300.446
R5914 bit5.n162 bit5.t32 300.446
R5915 bit5.n171 bit5.t1 300.446
R5916 bit5.n169 bit5.t26 300.446
R5917 bit5.n178 bit5.t17 300.446
R5918 bit5.n176 bit5.t44 300.446
R5919 bit5.n193 bit5.t30 300.446
R5920 bit5.n191 bit5.t20 300.446
R5921 bit5.n200 bit5.t38 300.446
R5922 bit5.n198 bit5.t51 300.446
R5923 bit5.n207 bit5.t54 300.446
R5924 bit5.n205 bit5.t0 300.446
R5925 bit5.n214 bit5.t19 300.446
R5926 bit5.n212 bit5.t27 300.446
R5927 bit5.n221 bit5.t48 300.446
R5928 bit5.n219 bit5.t57 300.446
R5929 bit5.n228 bit5.t7 300.446
R5930 bit5.n226 bit5.t62 300.446
R5931 bit5.n235 bit5.t14 300.446
R5932 bit5.n233 bit5.t22 300.446
R5933 bit5.n242 bit5.t47 300.446
R5934 bit5.n240 bit5.t56 300.446
R5935 bit5.n247 bit5.t23 279.56
R5936 bit5.n248 bit5.n247 120.317
R5937 bit5.n52 bit5.n51 27.537
R5938 bit5.n5 bit5.n2 27.536
R5939 bit5.n12 bit5.n9 27.536
R5940 bit5.n19 bit5.n16 27.536
R5941 bit5.n26 bit5.n23 27.536
R5942 bit5.n33 bit5.n30 27.536
R5943 bit5.n40 bit5.n37 27.536
R5944 bit5.n47 bit5.n44 27.536
R5945 bit5.n68 bit5.n65 27.536
R5946 bit5.n75 bit5.n72 27.536
R5947 bit5.n82 bit5.n79 27.536
R5948 bit5.n89 bit5.n86 27.536
R5949 bit5.n96 bit5.n93 27.536
R5950 bit5.n103 bit5.n100 27.536
R5951 bit5.n110 bit5.n107 27.536
R5952 bit5.n117 bit5.n114 27.536
R5953 bit5.n132 bit5.n129 27.536
R5954 bit5.n139 bit5.n136 27.536
R5955 bit5.n146 bit5.n143 27.536
R5956 bit5.n153 bit5.n150 27.536
R5957 bit5.n160 bit5.n157 27.536
R5958 bit5.n167 bit5.n164 27.536
R5959 bit5.n174 bit5.n171 27.536
R5960 bit5.n181 bit5.n178 27.536
R5961 bit5.n196 bit5.n193 27.536
R5962 bit5.n203 bit5.n200 27.536
R5963 bit5.n210 bit5.n207 27.536
R5964 bit5.n217 bit5.n214 27.536
R5965 bit5.n224 bit5.n221 27.536
R5966 bit5.n231 bit5.n228 27.536
R5967 bit5.n238 bit5.n235 27.536
R5968 bit5.n245 bit5.n242 27.536
R5969 bit5.n1 bit5.n0 24.127
R5970 bit5.n8 bit5.n7 24.127
R5971 bit5.n15 bit5.n14 24.127
R5972 bit5.n22 bit5.n21 24.127
R5973 bit5.n29 bit5.n28 24.127
R5974 bit5.n36 bit5.n35 24.127
R5975 bit5.n43 bit5.n42 24.127
R5976 bit5.n54 bit5.n53 24.127
R5977 bit5.n64 bit5.n63 24.127
R5978 bit5.n71 bit5.n70 24.127
R5979 bit5.n78 bit5.n77 24.127
R5980 bit5.n85 bit5.n84 24.127
R5981 bit5.n92 bit5.n91 24.127
R5982 bit5.n99 bit5.n98 24.127
R5983 bit5.n106 bit5.n105 24.127
R5984 bit5.n113 bit5.n112 24.127
R5985 bit5.n128 bit5.n127 24.127
R5986 bit5.n135 bit5.n134 24.127
R5987 bit5.n142 bit5.n141 24.127
R5988 bit5.n149 bit5.n148 24.127
R5989 bit5.n156 bit5.n155 24.127
R5990 bit5.n163 bit5.n162 24.127
R5991 bit5.n170 bit5.n169 24.127
R5992 bit5.n177 bit5.n176 24.127
R5993 bit5.n192 bit5.n191 24.127
R5994 bit5.n199 bit5.n198 24.127
R5995 bit5.n206 bit5.n205 24.127
R5996 bit5.n213 bit5.n212 24.127
R5997 bit5.n220 bit5.n219 24.127
R5998 bit5.n227 bit5.n226 24.127
R5999 bit5.n234 bit5.n233 24.127
R6000 bit5.n241 bit5.n240 24.127
R6001 bit5.n4 bit5.n3 8.764
R6002 bit5.n11 bit5.n10 8.764
R6003 bit5.n18 bit5.n17 8.764
R6004 bit5.n25 bit5.n24 8.764
R6005 bit5.n32 bit5.n31 8.764
R6006 bit5.n39 bit5.n38 8.764
R6007 bit5.n46 bit5.n45 8.764
R6008 bit5.n50 bit5.n49 8.764
R6009 bit5.n67 bit5.n66 8.764
R6010 bit5.n74 bit5.n73 8.764
R6011 bit5.n81 bit5.n80 8.764
R6012 bit5.n88 bit5.n87 8.764
R6013 bit5.n95 bit5.n94 8.764
R6014 bit5.n102 bit5.n101 8.764
R6015 bit5.n109 bit5.n108 8.764
R6016 bit5.n116 bit5.n115 8.764
R6017 bit5.n131 bit5.n130 8.764
R6018 bit5.n138 bit5.n137 8.764
R6019 bit5.n145 bit5.n144 8.764
R6020 bit5.n152 bit5.n151 8.764
R6021 bit5.n159 bit5.n158 8.764
R6022 bit5.n166 bit5.n165 8.764
R6023 bit5.n173 bit5.n172 8.764
R6024 bit5.n180 bit5.n179 8.764
R6025 bit5.n195 bit5.n194 8.764
R6026 bit5.n202 bit5.n201 8.764
R6027 bit5.n209 bit5.n208 8.764
R6028 bit5.n216 bit5.n215 8.764
R6029 bit5.n223 bit5.n222 8.764
R6030 bit5.n230 bit5.n229 8.764
R6031 bit5.n237 bit5.n236 8.764
R6032 bit5.n244 bit5.n243 8.764
R6033 bit5.n6 bit5.n1 4.662
R6034 bit5.n13 bit5.n8 4.662
R6035 bit5.n20 bit5.n15 4.662
R6036 bit5.n27 bit5.n22 4.662
R6037 bit5.n34 bit5.n29 4.662
R6038 bit5.n41 bit5.n36 4.662
R6039 bit5.n48 bit5.n43 4.662
R6040 bit5.n69 bit5.n64 4.662
R6041 bit5.n76 bit5.n71 4.662
R6042 bit5.n83 bit5.n78 4.662
R6043 bit5.n90 bit5.n85 4.662
R6044 bit5.n97 bit5.n92 4.662
R6045 bit5.n104 bit5.n99 4.662
R6046 bit5.n111 bit5.n106 4.662
R6047 bit5.n118 bit5.n113 4.662
R6048 bit5.n133 bit5.n128 4.662
R6049 bit5.n140 bit5.n135 4.662
R6050 bit5.n147 bit5.n142 4.662
R6051 bit5.n154 bit5.n149 4.662
R6052 bit5.n161 bit5.n156 4.662
R6053 bit5.n168 bit5.n163 4.662
R6054 bit5.n175 bit5.n170 4.662
R6055 bit5.n182 bit5.n177 4.662
R6056 bit5.n197 bit5.n192 4.662
R6057 bit5.n204 bit5.n199 4.662
R6058 bit5.n211 bit5.n206 4.662
R6059 bit5.n218 bit5.n213 4.662
R6060 bit5.n225 bit5.n220 4.662
R6061 bit5.n232 bit5.n227 4.662
R6062 bit5.n239 bit5.n234 4.662
R6063 bit5.n246 bit5.n241 4.662
R6064 bit5.n55 bit5.n54 4.661
R6065 bit5.n5 bit5.n4 3.401
R6066 bit5.n12 bit5.n11 3.401
R6067 bit5.n19 bit5.n18 3.401
R6068 bit5.n26 bit5.n25 3.401
R6069 bit5.n33 bit5.n32 3.401
R6070 bit5.n40 bit5.n39 3.401
R6071 bit5.n47 bit5.n46 3.401
R6072 bit5.n68 bit5.n67 3.401
R6073 bit5.n75 bit5.n74 3.401
R6074 bit5.n82 bit5.n81 3.401
R6075 bit5.n89 bit5.n88 3.401
R6076 bit5.n96 bit5.n95 3.401
R6077 bit5.n103 bit5.n102 3.401
R6078 bit5.n110 bit5.n109 3.401
R6079 bit5.n117 bit5.n116 3.401
R6080 bit5.n132 bit5.n131 3.401
R6081 bit5.n139 bit5.n138 3.401
R6082 bit5.n146 bit5.n145 3.401
R6083 bit5.n153 bit5.n152 3.401
R6084 bit5.n160 bit5.n159 3.401
R6085 bit5.n167 bit5.n166 3.401
R6086 bit5.n174 bit5.n173 3.401
R6087 bit5.n181 bit5.n180 3.401
R6088 bit5.n196 bit5.n195 3.401
R6089 bit5.n203 bit5.n202 3.401
R6090 bit5.n210 bit5.n209 3.401
R6091 bit5.n217 bit5.n216 3.401
R6092 bit5.n224 bit5.n223 3.401
R6093 bit5.n231 bit5.n230 3.401
R6094 bit5.n238 bit5.n237 3.401
R6095 bit5.n245 bit5.n244 3.401
R6096 bit5.n52 bit5.n50 3.401
R6097 bit5.n126 bit5.n62 1.218
R6098 bit5.n56 bit5.n55 0.873
R6099 bit5.n119 bit5.n118 0.873
R6100 bit5.n183 bit5.n182 0.873
R6101 bit5.n126 bit5.n125 0.726
R6102 bit5.n190 bit5.n189 0.726
R6103 bit5.n256 bit5.n255 0.726
R6104 bit5.n55 bit5.n52 0.626
R6105 bit5.n6 bit5.n5 0.626
R6106 bit5.n13 bit5.n12 0.626
R6107 bit5.n20 bit5.n19 0.626
R6108 bit5.n27 bit5.n26 0.626
R6109 bit5.n34 bit5.n33 0.626
R6110 bit5.n41 bit5.n40 0.626
R6111 bit5.n48 bit5.n47 0.626
R6112 bit5.n69 bit5.n68 0.626
R6113 bit5.n76 bit5.n75 0.626
R6114 bit5.n83 bit5.n82 0.626
R6115 bit5.n90 bit5.n89 0.626
R6116 bit5.n97 bit5.n96 0.626
R6117 bit5.n104 bit5.n103 0.626
R6118 bit5.n111 bit5.n110 0.626
R6119 bit5.n118 bit5.n117 0.626
R6120 bit5.n133 bit5.n132 0.626
R6121 bit5.n140 bit5.n139 0.626
R6122 bit5.n147 bit5.n146 0.626
R6123 bit5.n154 bit5.n153 0.626
R6124 bit5.n161 bit5.n160 0.626
R6125 bit5.n168 bit5.n167 0.626
R6126 bit5.n175 bit5.n174 0.626
R6127 bit5.n182 bit5.n181 0.626
R6128 bit5.n197 bit5.n196 0.626
R6129 bit5.n204 bit5.n203 0.626
R6130 bit5.n211 bit5.n210 0.626
R6131 bit5.n218 bit5.n217 0.626
R6132 bit5.n225 bit5.n224 0.626
R6133 bit5.n232 bit5.n231 0.626
R6134 bit5.n239 bit5.n238 0.626
R6135 bit5.n246 bit5.n245 0.626
R6136 bit5.n62 bit5.n61 0.575
R6137 bit5.n61 bit5.n60 0.575
R6138 bit5.n60 bit5.n59 0.575
R6139 bit5.n59 bit5.n58 0.575
R6140 bit5.n58 bit5.n57 0.575
R6141 bit5.n57 bit5.n56 0.575
R6142 bit5.n125 bit5.n124 0.575
R6143 bit5.n124 bit5.n123 0.575
R6144 bit5.n123 bit5.n122 0.575
R6145 bit5.n122 bit5.n121 0.575
R6146 bit5.n121 bit5.n120 0.575
R6147 bit5.n120 bit5.n119 0.575
R6148 bit5.n189 bit5.n188 0.575
R6149 bit5.n188 bit5.n187 0.575
R6150 bit5.n187 bit5.n186 0.575
R6151 bit5.n186 bit5.n185 0.575
R6152 bit5.n185 bit5.n184 0.575
R6153 bit5.n184 bit5.n183 0.575
R6154 bit5.n255 bit5.n254 0.575
R6155 bit5.n254 bit5.n253 0.575
R6156 bit5.n253 bit5.n252 0.575
R6157 bit5.n252 bit5.n251 0.575
R6158 bit5.n251 bit5.n250 0.575
R6159 bit5.n250 bit5.n249 0.575
R6160 bit5.n249 bit5.n248 0.575
R6161 bit5.n190 bit5.n126 0.492
R6162 bit5.n256 bit5.n190 0.492
R6163 bit5.n62 bit5.n6 0.298
R6164 bit5.n61 bit5.n13 0.298
R6165 bit5.n60 bit5.n20 0.298
R6166 bit5.n59 bit5.n27 0.298
R6167 bit5.n58 bit5.n34 0.298
R6168 bit5.n57 bit5.n41 0.298
R6169 bit5.n56 bit5.n48 0.298
R6170 bit5.n125 bit5.n69 0.298
R6171 bit5.n124 bit5.n76 0.298
R6172 bit5.n123 bit5.n83 0.298
R6173 bit5.n122 bit5.n90 0.298
R6174 bit5.n121 bit5.n97 0.298
R6175 bit5.n120 bit5.n104 0.298
R6176 bit5.n119 bit5.n111 0.298
R6177 bit5.n189 bit5.n133 0.298
R6178 bit5.n188 bit5.n140 0.298
R6179 bit5.n187 bit5.n147 0.298
R6180 bit5.n186 bit5.n154 0.298
R6181 bit5.n185 bit5.n161 0.298
R6182 bit5.n184 bit5.n168 0.298
R6183 bit5.n183 bit5.n175 0.298
R6184 bit5.n255 bit5.n197 0.298
R6185 bit5.n254 bit5.n204 0.298
R6186 bit5.n253 bit5.n211 0.298
R6187 bit5.n252 bit5.n218 0.298
R6188 bit5.n251 bit5.n225 0.298
R6189 bit5.n250 bit5.n232 0.298
R6190 bit5.n249 bit5.n239 0.298
R6191 bit5.n248 bit5.n246 0.298
R6192 bit5 bit5.n256 0.125
R6193 a_50466_6042.n26 a_50466_6042.t0 10.181
R6194 a_50466_6042.n18 a_50466_6042.t1 10.181
R6195 a_50466_6042.t3 a_50466_6042.n39 9.68
R6196 a_50466_6042.n3 a_50466_6042.n2 9.302
R6197 a_50466_6042.n13 a_50466_6042.n12 9.302
R6198 a_50466_6042.n32 a_50466_6042.n31 9.3
R6199 a_50466_6042.n34 a_50466_6042.n33 9.3
R6200 a_50466_6042.n7 a_50466_6042.n6 9.3
R6201 a_50466_6042.n5 a_50466_6042.n4 9.3
R6202 a_50466_6042.n36 a_50466_6042.n35 9
R6203 a_50466_6042.n9 a_50466_6042.n8 9
R6204 a_50466_6042.n27 a_50466_6042.n25 7.729
R6205 a_50466_6042.n19 a_50466_6042.n17 7.729
R6206 a_50466_6042.n27 a_50466_6042.n26 6.296
R6207 a_50466_6042.n19 a_50466_6042.n18 6.296
R6208 a_50466_6042.n30 a_50466_6042.n3 4.508
R6209 a_50466_6042.n14 a_50466_6042.n13 4.508
R6210 a_50466_6042.n37 a_50466_6042.n36 4.496
R6211 a_50466_6042.n21 a_50466_6042.n20 4.496
R6212 a_50466_6042.n29 a_50466_6042.n28 4.495
R6213 a_50466_6042.n10 a_50466_6042.n9 4.495
R6214 a_50466_6042.n14 a_50466_6042.n11 4.494
R6215 a_50466_6042.n30 a_50466_6042.n1 4.494
R6216 a_50466_6042.n39 a_50466_6042.t2 1.087
R6217 a_50466_6042.n25 a_50466_6042.n24 0.536
R6218 a_50466_6042.n17 a_50466_6042.n16 0.536
R6219 a_50466_6042.n39 a_50466_6042.n38 0.255
R6220 a_50466_6042.n28 a_50466_6042.n27 0.151
R6221 a_50466_6042.n20 a_50466_6042.n19 0.151
R6222 a_50466_6042.n23 a_50466_6042.n22 0.125
R6223 a_50466_6042.n34 a_50466_6042.n32 0.028
R6224 a_50466_6042.n7 a_50466_6042.n5 0.028
R6225 a_50466_6042.n1 a_50466_6042.n0 0.025
R6226 a_50466_6042.n20 a_50466_6042.n15 0.024
R6227 a_50466_6042.n36 a_50466_6042.n34 0.012
R6228 a_50466_6042.n9 a_50466_6042.n7 0.012
R6229 a_50466_6042.n29 a_50466_6042.n23 0.011
R6230 a_50466_6042.n30 a_50466_6042.n29 0.011
R6231 a_50466_6042.n14 a_50466_6042.n10 0.011
R6232 a_50466_6042.n38 a_50466_6042.n37 0.01
R6233 a_50466_6042.n22 a_50466_6042.n21 0.01
R6234 a_50466_6042.n21 a_50466_6042.n14 0.01
R6235 a_50466_6042.n37 a_50466_6042.n30 0.01
R6236 a_50176_5966.n10 a_50176_5966.t1 10.181
R6237 a_50176_5966.n10 a_50176_5966.t2 10.181
R6238 a_50176_5966.t0 a_50176_5966.n18 9.68
R6239 a_50176_5966.n1 a_50176_5966.n0 9.302
R6240 a_50176_5966.n7 a_50176_5966.n6 9.3
R6241 a_50176_5966.n5 a_50176_5966.n4 9.3
R6242 a_50176_5966.n9 a_50176_5966.n8 9
R6243 a_50176_5966.n13 a_50176_5966.n12 7.729
R6244 a_50176_5966.n13 a_50176_5966.n10 6.296
R6245 a_50176_5966.n16 a_50176_5966.n1 4.508
R6246 a_50176_5966.n15 a_50176_5966.n14 4.501
R6247 a_50176_5966.n15 a_50176_5966.n9 4.501
R6248 a_50176_5966.n16 a_50176_5966.n3 4.494
R6249 a_50176_5966.n18 a_50176_5966.t3 1.259
R6250 a_50176_5966.n12 a_50176_5966.n11 0.536
R6251 a_50176_5966.n18 a_50176_5966.n17 0.415
R6252 a_50176_5966.n14 a_50176_5966.n13 0.151
R6253 a_50176_5966.n7 a_50176_5966.n5 0.028
R6254 a_50176_5966.n3 a_50176_5966.n2 0.025
R6255 a_50176_5966.n17 a_50176_5966.n16 0.021
R6256 a_50176_5966.n9 a_50176_5966.n7 0.012
R6257 a_50176_5966.n16 a_50176_5966.n15 0.006
R6258 a_4176_94886.n10 a_4176_94886.t1 10.181
R6259 a_4176_94886.n10 a_4176_94886.t2 10.181
R6260 a_4176_94886.t0 a_4176_94886.n18 9.68
R6261 a_4176_94886.n1 a_4176_94886.n0 9.302
R6262 a_4176_94886.n7 a_4176_94886.n6 9.3
R6263 a_4176_94886.n5 a_4176_94886.n4 9.3
R6264 a_4176_94886.n9 a_4176_94886.n8 9
R6265 a_4176_94886.n13 a_4176_94886.n12 7.729
R6266 a_4176_94886.n13 a_4176_94886.n10 6.296
R6267 a_4176_94886.n16 a_4176_94886.n1 4.508
R6268 a_4176_94886.n15 a_4176_94886.n14 4.501
R6269 a_4176_94886.n15 a_4176_94886.n9 4.501
R6270 a_4176_94886.n16 a_4176_94886.n3 4.494
R6271 a_4176_94886.n18 a_4176_94886.t3 1.259
R6272 a_4176_94886.n12 a_4176_94886.n11 0.536
R6273 a_4176_94886.n18 a_4176_94886.n17 0.415
R6274 a_4176_94886.n14 a_4176_94886.n13 0.151
R6275 a_4176_94886.n7 a_4176_94886.n5 0.028
R6276 a_4176_94886.n3 a_4176_94886.n2 0.025
R6277 a_4176_94886.n17 a_4176_94886.n16 0.021
R6278 a_4176_94886.n9 a_4176_94886.n7 0.012
R6279 a_4176_94886.n16 a_4176_94886.n15 0.006
R6280 a_n436_94366.t1 a_n436_94366.n1 139.026
R6281 a_n436_94366.n1 a_n436_94366.t2 85.389
R6282 a_n436_94366.n1 a_n436_94366.n0 54.371
R6283 a_n436_94366.n0 a_n436_94366.t3 9.633
R6284 a_n436_94366.n0 a_n436_94366.t0 9.587
R6285 a_4176_55366.n10 a_4176_55366.t0 10.181
R6286 a_4176_55366.n10 a_4176_55366.t1 10.181
R6287 a_4176_55366.t3 a_4176_55366.n18 9.68
R6288 a_4176_55366.n1 a_4176_55366.n0 9.302
R6289 a_4176_55366.n7 a_4176_55366.n6 9.3
R6290 a_4176_55366.n5 a_4176_55366.n4 9.3
R6291 a_4176_55366.n9 a_4176_55366.n8 9
R6292 a_4176_55366.n13 a_4176_55366.n12 7.729
R6293 a_4176_55366.n13 a_4176_55366.n10 6.296
R6294 a_4176_55366.n16 a_4176_55366.n1 4.508
R6295 a_4176_55366.n15 a_4176_55366.n14 4.501
R6296 a_4176_55366.n15 a_4176_55366.n9 4.501
R6297 a_4176_55366.n16 a_4176_55366.n3 4.494
R6298 a_4176_55366.n18 a_4176_55366.t2 1.259
R6299 a_4176_55366.n12 a_4176_55366.n11 0.536
R6300 a_4176_55366.n18 a_4176_55366.n17 0.415
R6301 a_4176_55366.n14 a_4176_55366.n13 0.151
R6302 a_4176_55366.n7 a_4176_55366.n5 0.028
R6303 a_4176_55366.n3 a_4176_55366.n2 0.025
R6304 a_4176_55366.n17 a_4176_55366.n16 0.021
R6305 a_4176_55366.n9 a_4176_55366.n7 0.012
R6306 a_4176_55366.n16 a_4176_55366.n15 0.006
R6307 a_13376_15846.n10 a_13376_15846.t1 10.181
R6308 a_13376_15846.n10 a_13376_15846.t0 10.181
R6309 a_13376_15846.t3 a_13376_15846.n18 9.68
R6310 a_13376_15846.n1 a_13376_15846.n0 9.302
R6311 a_13376_15846.n7 a_13376_15846.n6 9.3
R6312 a_13376_15846.n5 a_13376_15846.n4 9.3
R6313 a_13376_15846.n9 a_13376_15846.n8 9
R6314 a_13376_15846.n13 a_13376_15846.n12 7.729
R6315 a_13376_15846.n13 a_13376_15846.n10 6.296
R6316 a_13376_15846.n16 a_13376_15846.n1 4.508
R6317 a_13376_15846.n15 a_13376_15846.n14 4.501
R6318 a_13376_15846.n15 a_13376_15846.n9 4.501
R6319 a_13376_15846.n16 a_13376_15846.n3 4.494
R6320 a_13376_15846.n18 a_13376_15846.t2 1.259
R6321 a_13376_15846.n12 a_13376_15846.n11 0.536
R6322 a_13376_15846.n18 a_13376_15846.n17 0.415
R6323 a_13376_15846.n14 a_13376_15846.n13 0.151
R6324 a_13376_15846.n7 a_13376_15846.n5 0.028
R6325 a_13376_15846.n3 a_13376_15846.n2 0.025
R6326 a_13376_15846.n17 a_13376_15846.n16 0.021
R6327 a_13376_15846.n9 a_13376_15846.n7 0.012
R6328 a_13376_15846.n16 a_13376_15846.n15 0.006
R6329 a_13666_15922.n26 a_13666_15922.t2 10.181
R6330 a_13666_15922.n18 a_13666_15922.t1 10.181
R6331 a_13666_15922.t0 a_13666_15922.n39 9.68
R6332 a_13666_15922.n3 a_13666_15922.n2 9.302
R6333 a_13666_15922.n13 a_13666_15922.n12 9.302
R6334 a_13666_15922.n32 a_13666_15922.n31 9.3
R6335 a_13666_15922.n34 a_13666_15922.n33 9.3
R6336 a_13666_15922.n7 a_13666_15922.n6 9.3
R6337 a_13666_15922.n5 a_13666_15922.n4 9.3
R6338 a_13666_15922.n36 a_13666_15922.n35 9
R6339 a_13666_15922.n9 a_13666_15922.n8 9
R6340 a_13666_15922.n27 a_13666_15922.n25 7.729
R6341 a_13666_15922.n19 a_13666_15922.n17 7.729
R6342 a_13666_15922.n27 a_13666_15922.n26 6.296
R6343 a_13666_15922.n19 a_13666_15922.n18 6.296
R6344 a_13666_15922.n30 a_13666_15922.n3 4.508
R6345 a_13666_15922.n14 a_13666_15922.n13 4.508
R6346 a_13666_15922.n37 a_13666_15922.n36 4.496
R6347 a_13666_15922.n21 a_13666_15922.n20 4.496
R6348 a_13666_15922.n29 a_13666_15922.n28 4.495
R6349 a_13666_15922.n10 a_13666_15922.n9 4.495
R6350 a_13666_15922.n14 a_13666_15922.n11 4.494
R6351 a_13666_15922.n30 a_13666_15922.n1 4.494
R6352 a_13666_15922.n39 a_13666_15922.t3 1.087
R6353 a_13666_15922.n25 a_13666_15922.n24 0.536
R6354 a_13666_15922.n17 a_13666_15922.n16 0.536
R6355 a_13666_15922.n39 a_13666_15922.n38 0.255
R6356 a_13666_15922.n28 a_13666_15922.n27 0.151
R6357 a_13666_15922.n20 a_13666_15922.n19 0.151
R6358 a_13666_15922.n23 a_13666_15922.n22 0.125
R6359 a_13666_15922.n34 a_13666_15922.n32 0.028
R6360 a_13666_15922.n7 a_13666_15922.n5 0.028
R6361 a_13666_15922.n1 a_13666_15922.n0 0.025
R6362 a_13666_15922.n20 a_13666_15922.n15 0.024
R6363 a_13666_15922.n36 a_13666_15922.n34 0.012
R6364 a_13666_15922.n9 a_13666_15922.n7 0.012
R6365 a_13666_15922.n29 a_13666_15922.n23 0.011
R6366 a_13666_15922.n30 a_13666_15922.n29 0.011
R6367 a_13666_15922.n14 a_13666_15922.n10 0.011
R6368 a_13666_15922.n38 a_13666_15922.n37 0.01
R6369 a_13666_15922.n22 a_13666_15922.n21 0.01
R6370 a_13666_15922.n21 a_13666_15922.n14 0.01
R6371 a_13666_15922.n37 a_13666_15922.n30 0.01
R6372 a_4176_15846.n10 a_4176_15846.t2 10.181
R6373 a_4176_15846.n10 a_4176_15846.t1 10.181
R6374 a_4176_15846.t0 a_4176_15846.n18 9.68
R6375 a_4176_15846.n1 a_4176_15846.n0 9.302
R6376 a_4176_15846.n7 a_4176_15846.n6 9.3
R6377 a_4176_15846.n5 a_4176_15846.n4 9.3
R6378 a_4176_15846.n9 a_4176_15846.n8 9
R6379 a_4176_15846.n13 a_4176_15846.n12 7.729
R6380 a_4176_15846.n13 a_4176_15846.n10 6.296
R6381 a_4176_15846.n16 a_4176_15846.n1 4.508
R6382 a_4176_15846.n15 a_4176_15846.n14 4.501
R6383 a_4176_15846.n15 a_4176_15846.n9 4.501
R6384 a_4176_15846.n16 a_4176_15846.n3 4.494
R6385 a_4176_15846.n18 a_4176_15846.t3 1.259
R6386 a_4176_15846.n12 a_4176_15846.n11 0.536
R6387 a_4176_15846.n18 a_4176_15846.n17 0.415
R6388 a_4176_15846.n14 a_4176_15846.n13 0.151
R6389 a_4176_15846.n7 a_4176_15846.n5 0.028
R6390 a_4176_15846.n3 a_4176_15846.n2 0.025
R6391 a_4176_15846.n17 a_4176_15846.n16 0.021
R6392 a_4176_15846.n9 a_4176_15846.n7 0.012
R6393 a_4176_15846.n16 a_4176_15846.n15 0.006
R6394 a_n436_5446.t25 a_n436_5446.n63 139.026
R6395 a_n436_5446.n63 a_n436_5446.t24 85.389
R6396 a_n436_5446.n63 a_n436_5446.n62 54.371
R6397 a_n436_5446.n0 a_n436_5446.t44 9.633
R6398 a_n436_5446.n15 a_n436_5446.t54 9.633
R6399 a_n436_5446.n31 a_n436_5446.t8 9.633
R6400 a_n436_5446.n0 a_n436_5446.t35 9.587
R6401 a_n436_5446.n1 a_n436_5446.t65 9.587
R6402 a_n436_5446.n2 a_n436_5446.t59 9.587
R6403 a_n436_5446.n3 a_n436_5446.t27 9.587
R6404 a_n436_5446.n4 a_n436_5446.t51 9.587
R6405 a_n436_5446.n5 a_n436_5446.t42 9.587
R6406 a_n436_5446.n6 a_n436_5446.t53 9.587
R6407 a_n436_5446.n7 a_n436_5446.t21 9.587
R6408 a_n436_5446.n8 a_n436_5446.t7 9.587
R6409 a_n436_5446.n9 a_n436_5446.t57 9.587
R6410 a_n436_5446.n10 a_n436_5446.t28 9.587
R6411 a_n436_5446.n11 a_n436_5446.t15 9.587
R6412 a_n436_5446.n12 a_n436_5446.t5 9.587
R6413 a_n436_5446.n13 a_n436_5446.t16 9.587
R6414 a_n436_5446.n14 a_n436_5446.t62 9.587
R6415 a_n436_5446.n15 a_n436_5446.t32 9.587
R6416 a_n436_5446.n16 a_n436_5446.t50 9.587
R6417 a_n436_5446.n17 a_n436_5446.t55 9.587
R6418 a_n436_5446.n18 a_n436_5446.t63 9.587
R6419 a_n436_5446.n19 a_n436_5446.t13 9.587
R6420 a_n436_5446.n20 a_n436_5446.t43 9.587
R6421 a_n436_5446.n21 a_n436_5446.t46 9.587
R6422 a_n436_5446.n22 a_n436_5446.t11 9.587
R6423 a_n436_5446.n23 a_n436_5446.t30 9.587
R6424 a_n436_5446.n24 a_n436_5446.t64 9.587
R6425 a_n436_5446.n25 a_n436_5446.t52 9.587
R6426 a_n436_5446.n26 a_n436_5446.t38 9.587
R6427 a_n436_5446.n27 a_n436_5446.t29 9.587
R6428 a_n436_5446.n28 a_n436_5446.t22 9.587
R6429 a_n436_5446.n29 a_n436_5446.t1 9.587
R6430 a_n436_5446.n31 a_n436_5446.t4 9.587
R6431 a_n436_5446.n32 a_n436_5446.t41 9.587
R6432 a_n436_5446.n33 a_n436_5446.t9 9.587
R6433 a_n436_5446.n34 a_n436_5446.t3 9.587
R6434 a_n436_5446.n35 a_n436_5446.t31 9.587
R6435 a_n436_5446.n36 a_n436_5446.t49 9.587
R6436 a_n436_5446.n37 a_n436_5446.t17 9.587
R6437 a_n436_5446.n38 a_n436_5446.t61 9.587
R6438 a_n436_5446.n39 a_n436_5446.t12 9.587
R6439 a_n436_5446.n40 a_n436_5446.t47 9.587
R6440 a_n436_5446.n41 a_n436_5446.t45 9.587
R6441 a_n436_5446.n42 a_n436_5446.t34 9.587
R6442 a_n436_5446.n43 a_n436_5446.t19 9.587
R6443 a_n436_5446.n44 a_n436_5446.t36 9.587
R6444 a_n436_5446.n45 a_n436_5446.t39 9.587
R6445 a_n436_5446.n62 a_n436_5446.t14 9.587
R6446 a_n436_5446.n61 a_n436_5446.t10 9.587
R6447 a_n436_5446.n60 a_n436_5446.t56 9.587
R6448 a_n436_5446.n59 a_n436_5446.t48 9.587
R6449 a_n436_5446.n58 a_n436_5446.t40 9.587
R6450 a_n436_5446.n57 a_n436_5446.t33 9.587
R6451 a_n436_5446.n56 a_n436_5446.t6 9.587
R6452 a_n436_5446.n55 a_n436_5446.t26 9.587
R6453 a_n436_5446.n54 a_n436_5446.t60 9.587
R6454 a_n436_5446.n53 a_n436_5446.t23 9.587
R6455 a_n436_5446.n52 a_n436_5446.t2 9.587
R6456 a_n436_5446.n51 a_n436_5446.t58 9.587
R6457 a_n436_5446.n50 a_n436_5446.t37 9.587
R6458 a_n436_5446.n49 a_n436_5446.t20 9.587
R6459 a_n436_5446.n48 a_n436_5446.t18 9.587
R6460 a_n436_5446.n47 a_n436_5446.t0 9.587
R6461 a_n436_5446.n30 a_n436_5446.n14 0.945
R6462 a_n436_5446.n47 a_n436_5446.n46 0.945
R6463 a_n436_5446.n13 a_n436_5446.n12 0.528
R6464 a_n436_5446.n11 a_n436_5446.n10 0.528
R6465 a_n436_5446.n9 a_n436_5446.n8 0.528
R6466 a_n436_5446.n7 a_n436_5446.n6 0.528
R6467 a_n436_5446.n5 a_n436_5446.n4 0.528
R6468 a_n436_5446.n3 a_n436_5446.n2 0.528
R6469 a_n436_5446.n1 a_n436_5446.n0 0.528
R6470 a_n436_5446.n28 a_n436_5446.n27 0.528
R6471 a_n436_5446.n26 a_n436_5446.n25 0.528
R6472 a_n436_5446.n24 a_n436_5446.n23 0.528
R6473 a_n436_5446.n22 a_n436_5446.n21 0.528
R6474 a_n436_5446.n20 a_n436_5446.n19 0.528
R6475 a_n436_5446.n18 a_n436_5446.n17 0.528
R6476 a_n436_5446.n16 a_n436_5446.n15 0.528
R6477 a_n436_5446.n44 a_n436_5446.n43 0.528
R6478 a_n436_5446.n42 a_n436_5446.n41 0.528
R6479 a_n436_5446.n40 a_n436_5446.n39 0.528
R6480 a_n436_5446.n38 a_n436_5446.n37 0.528
R6481 a_n436_5446.n36 a_n436_5446.n35 0.528
R6482 a_n436_5446.n34 a_n436_5446.n33 0.528
R6483 a_n436_5446.n32 a_n436_5446.n31 0.528
R6484 a_n436_5446.n49 a_n436_5446.n48 0.528
R6485 a_n436_5446.n51 a_n436_5446.n50 0.528
R6486 a_n436_5446.n53 a_n436_5446.n52 0.528
R6487 a_n436_5446.n55 a_n436_5446.n54 0.528
R6488 a_n436_5446.n57 a_n436_5446.n56 0.528
R6489 a_n436_5446.n59 a_n436_5446.n58 0.528
R6490 a_n436_5446.n61 a_n436_5446.n60 0.528
R6491 a_n436_5446.n46 a_n436_5446.n30 0.492
R6492 a_n436_5446.n30 a_n436_5446.n29 0.453
R6493 a_n436_5446.n46 a_n436_5446.n45 0.453
R6494 a_n436_5446.n14 a_n436_5446.n13 0.046
R6495 a_n436_5446.n12 a_n436_5446.n11 0.046
R6496 a_n436_5446.n10 a_n436_5446.n9 0.046
R6497 a_n436_5446.n8 a_n436_5446.n7 0.046
R6498 a_n436_5446.n6 a_n436_5446.n5 0.046
R6499 a_n436_5446.n4 a_n436_5446.n3 0.046
R6500 a_n436_5446.n2 a_n436_5446.n1 0.046
R6501 a_n436_5446.n29 a_n436_5446.n28 0.046
R6502 a_n436_5446.n27 a_n436_5446.n26 0.046
R6503 a_n436_5446.n25 a_n436_5446.n24 0.046
R6504 a_n436_5446.n23 a_n436_5446.n22 0.046
R6505 a_n436_5446.n21 a_n436_5446.n20 0.046
R6506 a_n436_5446.n19 a_n436_5446.n18 0.046
R6507 a_n436_5446.n17 a_n436_5446.n16 0.046
R6508 a_n436_5446.n45 a_n436_5446.n44 0.046
R6509 a_n436_5446.n43 a_n436_5446.n42 0.046
R6510 a_n436_5446.n41 a_n436_5446.n40 0.046
R6511 a_n436_5446.n39 a_n436_5446.n38 0.046
R6512 a_n436_5446.n37 a_n436_5446.n36 0.046
R6513 a_n436_5446.n35 a_n436_5446.n34 0.046
R6514 a_n436_5446.n33 a_n436_5446.n32 0.046
R6515 a_n436_5446.n48 a_n436_5446.n47 0.046
R6516 a_n436_5446.n50 a_n436_5446.n49 0.046
R6517 a_n436_5446.n52 a_n436_5446.n51 0.046
R6518 a_n436_5446.n54 a_n436_5446.n53 0.046
R6519 a_n436_5446.n56 a_n436_5446.n55 0.046
R6520 a_n436_5446.n58 a_n436_5446.n57 0.046
R6521 a_n436_5446.n60 a_n436_5446.n59 0.046
R6522 a_n436_5446.n62 a_n436_5446.n61 0.046
R6523 a_31776_25726.n10 a_31776_25726.t1 10.181
R6524 a_31776_25726.n10 a_31776_25726.t0 10.181
R6525 a_31776_25726.t3 a_31776_25726.n18 9.68
R6526 a_31776_25726.n1 a_31776_25726.n0 9.302
R6527 a_31776_25726.n7 a_31776_25726.n6 9.3
R6528 a_31776_25726.n5 a_31776_25726.n4 9.3
R6529 a_31776_25726.n9 a_31776_25726.n8 9
R6530 a_31776_25726.n13 a_31776_25726.n12 7.729
R6531 a_31776_25726.n13 a_31776_25726.n10 6.296
R6532 a_31776_25726.n16 a_31776_25726.n1 4.508
R6533 a_31776_25726.n15 a_31776_25726.n14 4.501
R6534 a_31776_25726.n15 a_31776_25726.n9 4.501
R6535 a_31776_25726.n16 a_31776_25726.n3 4.494
R6536 a_31776_25726.n18 a_31776_25726.t2 1.259
R6537 a_31776_25726.n12 a_31776_25726.n11 0.536
R6538 a_31776_25726.n18 a_31776_25726.n17 0.415
R6539 a_31776_25726.n14 a_31776_25726.n13 0.151
R6540 a_31776_25726.n7 a_31776_25726.n5 0.028
R6541 a_31776_25726.n3 a_31776_25726.n2 0.025
R6542 a_31776_25726.n17 a_31776_25726.n16 0.021
R6543 a_31776_25726.n9 a_31776_25726.n7 0.012
R6544 a_31776_25726.n16 a_31776_25726.n15 0.006
R6545 a_68866_45562.n26 a_68866_45562.t1 10.181
R6546 a_68866_45562.n18 a_68866_45562.t0 10.181
R6547 a_68866_45562.t3 a_68866_45562.n39 9.68
R6548 a_68866_45562.n3 a_68866_45562.n2 9.302
R6549 a_68866_45562.n13 a_68866_45562.n12 9.302
R6550 a_68866_45562.n32 a_68866_45562.n31 9.3
R6551 a_68866_45562.n34 a_68866_45562.n33 9.3
R6552 a_68866_45562.n7 a_68866_45562.n6 9.3
R6553 a_68866_45562.n5 a_68866_45562.n4 9.3
R6554 a_68866_45562.n36 a_68866_45562.n35 9
R6555 a_68866_45562.n9 a_68866_45562.n8 9
R6556 a_68866_45562.n27 a_68866_45562.n25 7.729
R6557 a_68866_45562.n19 a_68866_45562.n17 7.729
R6558 a_68866_45562.n27 a_68866_45562.n26 6.296
R6559 a_68866_45562.n19 a_68866_45562.n18 6.296
R6560 a_68866_45562.n30 a_68866_45562.n3 4.508
R6561 a_68866_45562.n14 a_68866_45562.n13 4.508
R6562 a_68866_45562.n37 a_68866_45562.n36 4.496
R6563 a_68866_45562.n21 a_68866_45562.n20 4.496
R6564 a_68866_45562.n29 a_68866_45562.n28 4.495
R6565 a_68866_45562.n10 a_68866_45562.n9 4.495
R6566 a_68866_45562.n14 a_68866_45562.n11 4.494
R6567 a_68866_45562.n30 a_68866_45562.n1 4.494
R6568 a_68866_45562.n39 a_68866_45562.t2 1.087
R6569 a_68866_45562.n25 a_68866_45562.n24 0.536
R6570 a_68866_45562.n17 a_68866_45562.n16 0.536
R6571 a_68866_45562.n39 a_68866_45562.n38 0.255
R6572 a_68866_45562.n28 a_68866_45562.n27 0.151
R6573 a_68866_45562.n20 a_68866_45562.n19 0.151
R6574 a_68866_45562.n23 a_68866_45562.n22 0.125
R6575 a_68866_45562.n34 a_68866_45562.n32 0.028
R6576 a_68866_45562.n7 a_68866_45562.n5 0.028
R6577 a_68866_45562.n1 a_68866_45562.n0 0.025
R6578 a_68866_45562.n20 a_68866_45562.n15 0.024
R6579 a_68866_45562.n36 a_68866_45562.n34 0.012
R6580 a_68866_45562.n9 a_68866_45562.n7 0.012
R6581 a_68866_45562.n29 a_68866_45562.n23 0.011
R6582 a_68866_45562.n30 a_68866_45562.n29 0.011
R6583 a_68866_45562.n14 a_68866_45562.n10 0.011
R6584 a_68866_45562.n38 a_68866_45562.n37 0.01
R6585 a_68866_45562.n22 a_68866_45562.n21 0.01
R6586 a_68866_45562.n21 a_68866_45562.n14 0.01
R6587 a_68866_45562.n37 a_68866_45562.n30 0.01
R6588 a_n436_44966.t9 a_n436_44966.n31 139.026
R6589 a_n436_44966.n31 a_n436_44966.t8 85.389
R6590 a_n436_44966.n31 a_n436_44966.n30 54.371
R6591 a_n436_44966.n0 a_n436_44966.t21 9.633
R6592 a_n436_44966.n0 a_n436_44966.t32 9.587
R6593 a_n436_44966.n1 a_n436_44966.t11 9.587
R6594 a_n436_44966.n2 a_n436_44966.t7 9.587
R6595 a_n436_44966.n3 a_n436_44966.t15 9.587
R6596 a_n436_44966.n4 a_n436_44966.t4 9.587
R6597 a_n436_44966.n5 a_n436_44966.t18 9.587
R6598 a_n436_44966.n6 a_n436_44966.t5 9.587
R6599 a_n436_44966.n7 a_n436_44966.t19 9.587
R6600 a_n436_44966.n8 a_n436_44966.t23 9.587
R6601 a_n436_44966.n9 a_n436_44966.t17 9.587
R6602 a_n436_44966.n10 a_n436_44966.t25 9.587
R6603 a_n436_44966.n11 a_n436_44966.t29 9.587
R6604 a_n436_44966.n12 a_n436_44966.t6 9.587
R6605 a_n436_44966.n13 a_n436_44966.t31 9.587
R6606 a_n436_44966.n14 a_n436_44966.t1 9.587
R6607 a_n436_44966.n30 a_n436_44966.t13 9.587
R6608 a_n436_44966.n29 a_n436_44966.t20 9.587
R6609 a_n436_44966.n28 a_n436_44966.t14 9.587
R6610 a_n436_44966.n27 a_n436_44966.t28 9.587
R6611 a_n436_44966.n26 a_n436_44966.t26 9.587
R6612 a_n436_44966.n25 a_n436_44966.t0 9.587
R6613 a_n436_44966.n24 a_n436_44966.t3 9.587
R6614 a_n436_44966.n23 a_n436_44966.t2 9.587
R6615 a_n436_44966.n22 a_n436_44966.t27 9.587
R6616 a_n436_44966.n21 a_n436_44966.t12 9.587
R6617 a_n436_44966.n20 a_n436_44966.t30 9.587
R6618 a_n436_44966.n19 a_n436_44966.t16 9.587
R6619 a_n436_44966.n18 a_n436_44966.t22 9.587
R6620 a_n436_44966.n17 a_n436_44966.t10 9.587
R6621 a_n436_44966.n16 a_n436_44966.t24 9.587
R6622 a_n436_44966.n15 a_n436_44966.t33 9.587
R6623 a_n436_44966.n15 a_n436_44966.n14 1.398
R6624 a_n436_44966.n13 a_n436_44966.n12 0.528
R6625 a_n436_44966.n11 a_n436_44966.n10 0.528
R6626 a_n436_44966.n9 a_n436_44966.n8 0.528
R6627 a_n436_44966.n7 a_n436_44966.n6 0.528
R6628 a_n436_44966.n5 a_n436_44966.n4 0.528
R6629 a_n436_44966.n3 a_n436_44966.n2 0.528
R6630 a_n436_44966.n1 a_n436_44966.n0 0.528
R6631 a_n436_44966.n17 a_n436_44966.n16 0.528
R6632 a_n436_44966.n19 a_n436_44966.n18 0.528
R6633 a_n436_44966.n21 a_n436_44966.n20 0.528
R6634 a_n436_44966.n23 a_n436_44966.n22 0.528
R6635 a_n436_44966.n25 a_n436_44966.n24 0.528
R6636 a_n436_44966.n27 a_n436_44966.n26 0.528
R6637 a_n436_44966.n29 a_n436_44966.n28 0.528
R6638 a_n436_44966.n14 a_n436_44966.n13 0.046
R6639 a_n436_44966.n12 a_n436_44966.n11 0.046
R6640 a_n436_44966.n10 a_n436_44966.n9 0.046
R6641 a_n436_44966.n8 a_n436_44966.n7 0.046
R6642 a_n436_44966.n6 a_n436_44966.n5 0.046
R6643 a_n436_44966.n4 a_n436_44966.n3 0.046
R6644 a_n436_44966.n2 a_n436_44966.n1 0.046
R6645 a_n436_44966.n16 a_n436_44966.n15 0.046
R6646 a_n436_44966.n18 a_n436_44966.n17 0.046
R6647 a_n436_44966.n20 a_n436_44966.n19 0.046
R6648 a_n436_44966.n22 a_n436_44966.n21 0.046
R6649 a_n436_44966.n24 a_n436_44966.n23 0.046
R6650 a_n436_44966.n26 a_n436_44966.n25 0.046
R6651 a_n436_44966.n28 a_n436_44966.n27 0.046
R6652 a_n436_44966.n30 a_n436_44966.n29 0.046
R6653 a_50466_45562.n26 a_50466_45562.t0 10.181
R6654 a_50466_45562.n18 a_50466_45562.t1 10.181
R6655 a_50466_45562.t2 a_50466_45562.n39 9.68
R6656 a_50466_45562.n3 a_50466_45562.n2 9.302
R6657 a_50466_45562.n13 a_50466_45562.n12 9.302
R6658 a_50466_45562.n32 a_50466_45562.n31 9.3
R6659 a_50466_45562.n34 a_50466_45562.n33 9.3
R6660 a_50466_45562.n7 a_50466_45562.n6 9.3
R6661 a_50466_45562.n5 a_50466_45562.n4 9.3
R6662 a_50466_45562.n36 a_50466_45562.n35 9
R6663 a_50466_45562.n9 a_50466_45562.n8 9
R6664 a_50466_45562.n27 a_50466_45562.n25 7.729
R6665 a_50466_45562.n19 a_50466_45562.n17 7.729
R6666 a_50466_45562.n27 a_50466_45562.n26 6.296
R6667 a_50466_45562.n19 a_50466_45562.n18 6.296
R6668 a_50466_45562.n30 a_50466_45562.n3 4.508
R6669 a_50466_45562.n14 a_50466_45562.n13 4.508
R6670 a_50466_45562.n37 a_50466_45562.n36 4.496
R6671 a_50466_45562.n21 a_50466_45562.n20 4.496
R6672 a_50466_45562.n29 a_50466_45562.n28 4.495
R6673 a_50466_45562.n10 a_50466_45562.n9 4.495
R6674 a_50466_45562.n14 a_50466_45562.n11 4.494
R6675 a_50466_45562.n30 a_50466_45562.n1 4.494
R6676 a_50466_45562.n39 a_50466_45562.t3 1.087
R6677 a_50466_45562.n25 a_50466_45562.n24 0.536
R6678 a_50466_45562.n17 a_50466_45562.n16 0.536
R6679 a_50466_45562.n39 a_50466_45562.n38 0.255
R6680 a_50466_45562.n28 a_50466_45562.n27 0.151
R6681 a_50466_45562.n20 a_50466_45562.n19 0.151
R6682 a_50466_45562.n23 a_50466_45562.n22 0.125
R6683 a_50466_45562.n34 a_50466_45562.n32 0.028
R6684 a_50466_45562.n7 a_50466_45562.n5 0.028
R6685 a_50466_45562.n1 a_50466_45562.n0 0.025
R6686 a_50466_45562.n20 a_50466_45562.n15 0.024
R6687 a_50466_45562.n36 a_50466_45562.n34 0.012
R6688 a_50466_45562.n9 a_50466_45562.n7 0.012
R6689 a_50466_45562.n29 a_50466_45562.n23 0.011
R6690 a_50466_45562.n30 a_50466_45562.n29 0.011
R6691 a_50466_45562.n14 a_50466_45562.n10 0.011
R6692 a_50466_45562.n38 a_50466_45562.n37 0.01
R6693 a_50466_45562.n22 a_50466_45562.n21 0.01
R6694 a_50466_45562.n21 a_50466_45562.n14 0.01
R6695 a_50466_45562.n37 a_50466_45562.n30 0.01
R6696 a_50176_45486.n10 a_50176_45486.t0 10.181
R6697 a_50176_45486.n10 a_50176_45486.t1 10.181
R6698 a_50176_45486.t3 a_50176_45486.n18 9.68
R6699 a_50176_45486.n1 a_50176_45486.n0 9.302
R6700 a_50176_45486.n7 a_50176_45486.n6 9.3
R6701 a_50176_45486.n5 a_50176_45486.n4 9.3
R6702 a_50176_45486.n9 a_50176_45486.n8 9
R6703 a_50176_45486.n13 a_50176_45486.n12 7.729
R6704 a_50176_45486.n13 a_50176_45486.n10 6.296
R6705 a_50176_45486.n16 a_50176_45486.n1 4.508
R6706 a_50176_45486.n15 a_50176_45486.n14 4.501
R6707 a_50176_45486.n15 a_50176_45486.n9 4.501
R6708 a_50176_45486.n16 a_50176_45486.n3 4.494
R6709 a_50176_45486.n18 a_50176_45486.t2 1.259
R6710 a_50176_45486.n12 a_50176_45486.n11 0.536
R6711 a_50176_45486.n18 a_50176_45486.n17 0.415
R6712 a_50176_45486.n14 a_50176_45486.n13 0.151
R6713 a_50176_45486.n7 a_50176_45486.n5 0.028
R6714 a_50176_45486.n3 a_50176_45486.n2 0.025
R6715 a_50176_45486.n17 a_50176_45486.n16 0.021
R6716 a_50176_45486.n9 a_50176_45486.n7 0.012
R6717 a_50176_45486.n16 a_50176_45486.n15 0.006
R6718 a_50176_55366.n10 a_50176_55366.t0 10.181
R6719 a_50176_55366.n10 a_50176_55366.t1 10.181
R6720 a_50176_55366.t2 a_50176_55366.n18 9.68
R6721 a_50176_55366.n1 a_50176_55366.n0 9.302
R6722 a_50176_55366.n7 a_50176_55366.n6 9.3
R6723 a_50176_55366.n5 a_50176_55366.n4 9.3
R6724 a_50176_55366.n9 a_50176_55366.n8 9
R6725 a_50176_55366.n13 a_50176_55366.n12 7.729
R6726 a_50176_55366.n13 a_50176_55366.n10 6.296
R6727 a_50176_55366.n16 a_50176_55366.n1 4.508
R6728 a_50176_55366.n15 a_50176_55366.n14 4.501
R6729 a_50176_55366.n15 a_50176_55366.n9 4.501
R6730 a_50176_55366.n16 a_50176_55366.n3 4.494
R6731 a_50176_55366.n18 a_50176_55366.t3 1.259
R6732 a_50176_55366.n12 a_50176_55366.n11 0.536
R6733 a_50176_55366.n18 a_50176_55366.n17 0.415
R6734 a_50176_55366.n14 a_50176_55366.n13 0.151
R6735 a_50176_55366.n7 a_50176_55366.n5 0.028
R6736 a_50176_55366.n3 a_50176_55366.n2 0.025
R6737 a_50176_55366.n17 a_50176_55366.n16 0.021
R6738 a_50176_55366.n9 a_50176_55366.n7 0.012
R6739 a_50176_55366.n16 a_50176_55366.n15 0.006
R6740 OUT_N.n61 OUT_N.n5 1.013
R6741 OUT_N.n58 OUT_N.n23 1.013
R6742 OUT_N.n59 OUT_N.n17 1.013
R6743 OUT_N.n60 OUT_N.n11 1.013
R6744 OUT_N.n56 OUT_N.n37 0.781
R6745 OUT_N.n57 OUT_N.n30 0.781
R6746 OUT_N.n55 OUT_N.n45 0.549
R6747 OUT_N.n55 OUT_N.n54 0.532
R6748 OUT_N.n0 OUT_N.t9 0.359
R6749 OUT_N.n46 OUT_N.t41 0.359
R6750 OUT_N.n38 OUT_N.t23 0.359
R6751 OUT_N.n31 OUT_N.t27 0.359
R6752 OUT_N.n24 OUT_N.t33 0.359
R6753 OUT_N.n18 OUT_N.t24 0.359
R6754 OUT_N.n12 OUT_N.t30 0.359
R6755 OUT_N.n6 OUT_N.t36 0.359
R6756 OUT_N OUT_N.n61 0.257
R6757 OUT_N.n1 OUT_N.n0 0.23
R6758 OUT_N.n2 OUT_N.n1 0.23
R6759 OUT_N.n3 OUT_N.n2 0.23
R6760 OUT_N.n4 OUT_N.n3 0.23
R6761 OUT_N.n5 OUT_N.n4 0.23
R6762 OUT_N.n47 OUT_N.n46 0.23
R6763 OUT_N.n48 OUT_N.n47 0.23
R6764 OUT_N.n49 OUT_N.n48 0.23
R6765 OUT_N.n50 OUT_N.n49 0.23
R6766 OUT_N.n51 OUT_N.n50 0.23
R6767 OUT_N.n52 OUT_N.n51 0.23
R6768 OUT_N.n53 OUT_N.n52 0.23
R6769 OUT_N.n54 OUT_N.n53 0.23
R6770 OUT_N.n39 OUT_N.n38 0.23
R6771 OUT_N.n40 OUT_N.n39 0.23
R6772 OUT_N.n41 OUT_N.n40 0.23
R6773 OUT_N.n42 OUT_N.n41 0.23
R6774 OUT_N.n43 OUT_N.n42 0.23
R6775 OUT_N.n44 OUT_N.n43 0.23
R6776 OUT_N.n45 OUT_N.n44 0.23
R6777 OUT_N.n32 OUT_N.n31 0.23
R6778 OUT_N.n33 OUT_N.n32 0.23
R6779 OUT_N.n34 OUT_N.n33 0.23
R6780 OUT_N.n35 OUT_N.n34 0.23
R6781 OUT_N.n36 OUT_N.n35 0.23
R6782 OUT_N.n37 OUT_N.n36 0.23
R6783 OUT_N.n25 OUT_N.n24 0.23
R6784 OUT_N.n26 OUT_N.n25 0.23
R6785 OUT_N.n27 OUT_N.n26 0.23
R6786 OUT_N.n28 OUT_N.n27 0.23
R6787 OUT_N.n29 OUT_N.n28 0.23
R6788 OUT_N.n30 OUT_N.n29 0.23
R6789 OUT_N.n19 OUT_N.n18 0.23
R6790 OUT_N.n20 OUT_N.n19 0.23
R6791 OUT_N.n21 OUT_N.n20 0.23
R6792 OUT_N.n22 OUT_N.n21 0.23
R6793 OUT_N.n23 OUT_N.n22 0.23
R6794 OUT_N.n13 OUT_N.n12 0.23
R6795 OUT_N.n14 OUT_N.n13 0.23
R6796 OUT_N.n15 OUT_N.n14 0.23
R6797 OUT_N.n16 OUT_N.n15 0.23
R6798 OUT_N.n17 OUT_N.n16 0.23
R6799 OUT_N.n7 OUT_N.n6 0.23
R6800 OUT_N.n8 OUT_N.n7 0.23
R6801 OUT_N.n9 OUT_N.n8 0.23
R6802 OUT_N.n10 OUT_N.n9 0.23
R6803 OUT_N.n11 OUT_N.n10 0.23
R6804 OUT_N.n60 OUT_N.n59 0.215
R6805 OUT_N.n59 OUT_N.n58 0.215
R6806 OUT_N.n58 OUT_N.n57 0.215
R6807 OUT_N.n57 OUT_N.n56 0.215
R6808 OUT_N.n56 OUT_N.n55 0.215
R6809 OUT_N.n61 OUT_N.n60 0.214
R6810 OUT_N.n5 OUT_N.t13 0.129
R6811 OUT_N.n4 OUT_N.t51 0.129
R6812 OUT_N.n3 OUT_N.t25 0.129
R6813 OUT_N.n2 OUT_N.t0 0.129
R6814 OUT_N.n1 OUT_N.t48 0.129
R6815 OUT_N.n0 OUT_N.t19 0.129
R6816 OUT_N.n54 OUT_N.t4 0.129
R6817 OUT_N.n53 OUT_N.t12 0.129
R6818 OUT_N.n52 OUT_N.t53 0.129
R6819 OUT_N.n51 OUT_N.t28 0.129
R6820 OUT_N.n50 OUT_N.t3 0.129
R6821 OUT_N.n49 OUT_N.t44 0.129
R6822 OUT_N.n48 OUT_N.t17 0.129
R6823 OUT_N.n47 OUT_N.t60 0.129
R6824 OUT_N.n46 OUT_N.t38 0.129
R6825 OUT_N.n45 OUT_N.t52 0.129
R6826 OUT_N.n44 OUT_N.t34 0.129
R6827 OUT_N.n43 OUT_N.t7 0.129
R6828 OUT_N.n42 OUT_N.t49 0.129
R6829 OUT_N.n41 OUT_N.t21 0.129
R6830 OUT_N.n40 OUT_N.t59 0.129
R6831 OUT_N.n39 OUT_N.t40 0.129
R6832 OUT_N.n38 OUT_N.t11 0.129
R6833 OUT_N.n37 OUT_N.t57 0.129
R6834 OUT_N.n36 OUT_N.t31 0.129
R6835 OUT_N.n35 OUT_N.t6 0.129
R6836 OUT_N.n34 OUT_N.t47 0.129
R6837 OUT_N.n33 OUT_N.t20 0.129
R6838 OUT_N.n32 OUT_N.t62 0.129
R6839 OUT_N.n31 OUT_N.t39 0.129
R6840 OUT_N.n30 OUT_N.t15 0.129
R6841 OUT_N.n29 OUT_N.t54 0.129
R6842 OUT_N.n28 OUT_N.t29 0.129
R6843 OUT_N.n27 OUT_N.t5 0.129
R6844 OUT_N.n26 OUT_N.t45 0.129
R6845 OUT_N.n25 OUT_N.t22 0.129
R6846 OUT_N.n24 OUT_N.t61 0.129
R6847 OUT_N.n23 OUT_N.t46 0.129
R6848 OUT_N.n22 OUT_N.t18 0.129
R6849 OUT_N.n21 OUT_N.t56 0.129
R6850 OUT_N.n20 OUT_N.t32 0.129
R6851 OUT_N.n19 OUT_N.t10 0.129
R6852 OUT_N.n18 OUT_N.t50 0.129
R6853 OUT_N.n17 OUT_N.t2 0.129
R6854 OUT_N.n16 OUT_N.t43 0.129
R6855 OUT_N.n15 OUT_N.t16 0.129
R6856 OUT_N.n14 OUT_N.t55 0.129
R6857 OUT_N.n13 OUT_N.t37 0.129
R6858 OUT_N.n12 OUT_N.t8 0.129
R6859 OUT_N.n11 OUT_N.t26 0.129
R6860 OUT_N.n10 OUT_N.t1 0.129
R6861 OUT_N.n9 OUT_N.t42 0.129
R6862 OUT_N.n8 OUT_N.t14 0.129
R6863 OUT_N.n7 OUT_N.t58 0.129
R6864 OUT_N.n6 OUT_N.t35 0.129
R6865 a_68866_35682.n26 a_68866_35682.t0 10.181
R6866 a_68866_35682.n18 a_68866_35682.t1 10.181
R6867 a_68866_35682.t3 a_68866_35682.n39 9.68
R6868 a_68866_35682.n3 a_68866_35682.n2 9.302
R6869 a_68866_35682.n13 a_68866_35682.n12 9.302
R6870 a_68866_35682.n32 a_68866_35682.n31 9.3
R6871 a_68866_35682.n34 a_68866_35682.n33 9.3
R6872 a_68866_35682.n7 a_68866_35682.n6 9.3
R6873 a_68866_35682.n5 a_68866_35682.n4 9.3
R6874 a_68866_35682.n36 a_68866_35682.n35 9
R6875 a_68866_35682.n9 a_68866_35682.n8 9
R6876 a_68866_35682.n27 a_68866_35682.n25 7.729
R6877 a_68866_35682.n19 a_68866_35682.n17 7.729
R6878 a_68866_35682.n27 a_68866_35682.n26 6.296
R6879 a_68866_35682.n19 a_68866_35682.n18 6.296
R6880 a_68866_35682.n30 a_68866_35682.n3 4.508
R6881 a_68866_35682.n14 a_68866_35682.n13 4.508
R6882 a_68866_35682.n37 a_68866_35682.n36 4.496
R6883 a_68866_35682.n21 a_68866_35682.n20 4.496
R6884 a_68866_35682.n29 a_68866_35682.n28 4.495
R6885 a_68866_35682.n10 a_68866_35682.n9 4.495
R6886 a_68866_35682.n14 a_68866_35682.n11 4.494
R6887 a_68866_35682.n30 a_68866_35682.n1 4.494
R6888 a_68866_35682.n39 a_68866_35682.t2 1.087
R6889 a_68866_35682.n25 a_68866_35682.n24 0.536
R6890 a_68866_35682.n17 a_68866_35682.n16 0.536
R6891 a_68866_35682.n39 a_68866_35682.n38 0.255
R6892 a_68866_35682.n28 a_68866_35682.n27 0.151
R6893 a_68866_35682.n20 a_68866_35682.n19 0.151
R6894 a_68866_35682.n23 a_68866_35682.n22 0.125
R6895 a_68866_35682.n34 a_68866_35682.n32 0.028
R6896 a_68866_35682.n7 a_68866_35682.n5 0.028
R6897 a_68866_35682.n1 a_68866_35682.n0 0.025
R6898 a_68866_35682.n20 a_68866_35682.n15 0.024
R6899 a_68866_35682.n36 a_68866_35682.n34 0.012
R6900 a_68866_35682.n9 a_68866_35682.n7 0.012
R6901 a_68866_35682.n29 a_68866_35682.n23 0.011
R6902 a_68866_35682.n30 a_68866_35682.n29 0.011
R6903 a_68866_35682.n14 a_68866_35682.n10 0.011
R6904 a_68866_35682.n38 a_68866_35682.n37 0.01
R6905 a_68866_35682.n22 a_68866_35682.n21 0.01
R6906 a_68866_35682.n21 a_68866_35682.n14 0.01
R6907 a_68866_35682.n37 a_68866_35682.n30 0.01
R6908 a_31776_45486.n10 a_31776_45486.t2 10.181
R6909 a_31776_45486.n10 a_31776_45486.t1 10.181
R6910 a_31776_45486.t0 a_31776_45486.n18 9.68
R6911 a_31776_45486.n1 a_31776_45486.n0 9.302
R6912 a_31776_45486.n7 a_31776_45486.n6 9.3
R6913 a_31776_45486.n5 a_31776_45486.n4 9.3
R6914 a_31776_45486.n9 a_31776_45486.n8 9
R6915 a_31776_45486.n13 a_31776_45486.n12 7.729
R6916 a_31776_45486.n13 a_31776_45486.n10 6.296
R6917 a_31776_45486.n16 a_31776_45486.n1 4.508
R6918 a_31776_45486.n15 a_31776_45486.n14 4.501
R6919 a_31776_45486.n15 a_31776_45486.n9 4.501
R6920 a_31776_45486.n16 a_31776_45486.n3 4.494
R6921 a_31776_45486.n18 a_31776_45486.t3 1.259
R6922 a_31776_45486.n12 a_31776_45486.n11 0.536
R6923 a_31776_45486.n18 a_31776_45486.n17 0.415
R6924 a_31776_45486.n14 a_31776_45486.n13 0.151
R6925 a_31776_45486.n7 a_31776_45486.n5 0.028
R6926 a_31776_45486.n3 a_31776_45486.n2 0.025
R6927 a_31776_45486.n17 a_31776_45486.n16 0.021
R6928 a_31776_45486.n9 a_31776_45486.n7 0.012
R6929 a_31776_45486.n16 a_31776_45486.n15 0.006
R6930 a_59666_55442.n26 a_59666_55442.t2 10.181
R6931 a_59666_55442.n18 a_59666_55442.t1 10.181
R6932 a_59666_55442.t0 a_59666_55442.n39 9.68
R6933 a_59666_55442.n3 a_59666_55442.n2 9.302
R6934 a_59666_55442.n13 a_59666_55442.n12 9.302
R6935 a_59666_55442.n32 a_59666_55442.n31 9.3
R6936 a_59666_55442.n34 a_59666_55442.n33 9.3
R6937 a_59666_55442.n7 a_59666_55442.n6 9.3
R6938 a_59666_55442.n5 a_59666_55442.n4 9.3
R6939 a_59666_55442.n36 a_59666_55442.n35 9
R6940 a_59666_55442.n9 a_59666_55442.n8 9
R6941 a_59666_55442.n27 a_59666_55442.n25 7.729
R6942 a_59666_55442.n19 a_59666_55442.n17 7.729
R6943 a_59666_55442.n27 a_59666_55442.n26 6.296
R6944 a_59666_55442.n19 a_59666_55442.n18 6.296
R6945 a_59666_55442.n30 a_59666_55442.n3 4.508
R6946 a_59666_55442.n14 a_59666_55442.n13 4.508
R6947 a_59666_55442.n37 a_59666_55442.n36 4.496
R6948 a_59666_55442.n21 a_59666_55442.n20 4.496
R6949 a_59666_55442.n29 a_59666_55442.n28 4.495
R6950 a_59666_55442.n10 a_59666_55442.n9 4.495
R6951 a_59666_55442.n14 a_59666_55442.n11 4.494
R6952 a_59666_55442.n30 a_59666_55442.n1 4.494
R6953 a_59666_55442.n39 a_59666_55442.t3 1.087
R6954 a_59666_55442.n25 a_59666_55442.n24 0.536
R6955 a_59666_55442.n17 a_59666_55442.n16 0.536
R6956 a_59666_55442.n39 a_59666_55442.n38 0.255
R6957 a_59666_55442.n28 a_59666_55442.n27 0.151
R6958 a_59666_55442.n20 a_59666_55442.n19 0.151
R6959 a_59666_55442.n23 a_59666_55442.n22 0.125
R6960 a_59666_55442.n34 a_59666_55442.n32 0.028
R6961 a_59666_55442.n7 a_59666_55442.n5 0.028
R6962 a_59666_55442.n1 a_59666_55442.n0 0.025
R6963 a_59666_55442.n20 a_59666_55442.n15 0.024
R6964 a_59666_55442.n36 a_59666_55442.n34 0.012
R6965 a_59666_55442.n9 a_59666_55442.n7 0.012
R6966 a_59666_55442.n29 a_59666_55442.n23 0.011
R6967 a_59666_55442.n30 a_59666_55442.n29 0.011
R6968 a_59666_55442.n14 a_59666_55442.n10 0.011
R6969 a_59666_55442.n38 a_59666_55442.n37 0.01
R6970 a_59666_55442.n22 a_59666_55442.n21 0.01
R6971 a_59666_55442.n21 a_59666_55442.n14 0.01
R6972 a_59666_55442.n37 a_59666_55442.n30 0.01
R6973 a_13376_35606.n10 a_13376_35606.t1 10.181
R6974 a_13376_35606.n10 a_13376_35606.t0 10.181
R6975 a_13376_35606.t3 a_13376_35606.n18 9.68
R6976 a_13376_35606.n1 a_13376_35606.n0 9.302
R6977 a_13376_35606.n7 a_13376_35606.n6 9.3
R6978 a_13376_35606.n5 a_13376_35606.n4 9.3
R6979 a_13376_35606.n9 a_13376_35606.n8 9
R6980 a_13376_35606.n13 a_13376_35606.n12 7.729
R6981 a_13376_35606.n13 a_13376_35606.n10 6.296
R6982 a_13376_35606.n16 a_13376_35606.n1 4.508
R6983 a_13376_35606.n15 a_13376_35606.n14 4.501
R6984 a_13376_35606.n15 a_13376_35606.n9 4.501
R6985 a_13376_35606.n16 a_13376_35606.n3 4.494
R6986 a_13376_35606.n18 a_13376_35606.t2 1.259
R6987 a_13376_35606.n12 a_13376_35606.n11 0.536
R6988 a_13376_35606.n18 a_13376_35606.n17 0.415
R6989 a_13376_35606.n14 a_13376_35606.n13 0.151
R6990 a_13376_35606.n7 a_13376_35606.n5 0.028
R6991 a_13376_35606.n3 a_13376_35606.n2 0.025
R6992 a_13376_35606.n17 a_13376_35606.n16 0.021
R6993 a_13376_35606.n9 a_13376_35606.n7 0.012
R6994 a_13376_35606.n16 a_13376_35606.n15 0.006
R6995 a_40976_15846.n10 a_40976_15846.t1 10.181
R6996 a_40976_15846.n10 a_40976_15846.t0 10.181
R6997 a_40976_15846.t3 a_40976_15846.n18 9.68
R6998 a_40976_15846.n1 a_40976_15846.n0 9.302
R6999 a_40976_15846.n7 a_40976_15846.n6 9.3
R7000 a_40976_15846.n5 a_40976_15846.n4 9.3
R7001 a_40976_15846.n9 a_40976_15846.n8 9
R7002 a_40976_15846.n13 a_40976_15846.n12 7.729
R7003 a_40976_15846.n13 a_40976_15846.n10 6.296
R7004 a_40976_15846.n16 a_40976_15846.n1 4.508
R7005 a_40976_15846.n15 a_40976_15846.n14 4.501
R7006 a_40976_15846.n15 a_40976_15846.n9 4.501
R7007 a_40976_15846.n16 a_40976_15846.n3 4.494
R7008 a_40976_15846.n18 a_40976_15846.t2 1.259
R7009 a_40976_15846.n12 a_40976_15846.n11 0.536
R7010 a_40976_15846.n18 a_40976_15846.n17 0.415
R7011 a_40976_15846.n14 a_40976_15846.n13 0.151
R7012 a_40976_15846.n7 a_40976_15846.n5 0.028
R7013 a_40976_15846.n3 a_40976_15846.n2 0.025
R7014 a_40976_15846.n17 a_40976_15846.n16 0.021
R7015 a_40976_15846.n9 a_40976_15846.n7 0.012
R7016 a_40976_15846.n16 a_40976_15846.n15 0.006
R7017 a_41266_15922.n26 a_41266_15922.t2 10.181
R7018 a_41266_15922.n18 a_41266_15922.t1 10.181
R7019 a_41266_15922.t0 a_41266_15922.n39 9.68
R7020 a_41266_15922.n3 a_41266_15922.n2 9.302
R7021 a_41266_15922.n13 a_41266_15922.n12 9.302
R7022 a_41266_15922.n32 a_41266_15922.n31 9.3
R7023 a_41266_15922.n34 a_41266_15922.n33 9.3
R7024 a_41266_15922.n7 a_41266_15922.n6 9.3
R7025 a_41266_15922.n5 a_41266_15922.n4 9.3
R7026 a_41266_15922.n36 a_41266_15922.n35 9
R7027 a_41266_15922.n9 a_41266_15922.n8 9
R7028 a_41266_15922.n27 a_41266_15922.n25 7.729
R7029 a_41266_15922.n19 a_41266_15922.n17 7.729
R7030 a_41266_15922.n27 a_41266_15922.n26 6.296
R7031 a_41266_15922.n19 a_41266_15922.n18 6.296
R7032 a_41266_15922.n30 a_41266_15922.n3 4.508
R7033 a_41266_15922.n14 a_41266_15922.n13 4.508
R7034 a_41266_15922.n37 a_41266_15922.n36 4.496
R7035 a_41266_15922.n21 a_41266_15922.n20 4.496
R7036 a_41266_15922.n29 a_41266_15922.n28 4.495
R7037 a_41266_15922.n10 a_41266_15922.n9 4.495
R7038 a_41266_15922.n14 a_41266_15922.n11 4.494
R7039 a_41266_15922.n30 a_41266_15922.n1 4.494
R7040 a_41266_15922.n39 a_41266_15922.t3 1.087
R7041 a_41266_15922.n25 a_41266_15922.n24 0.536
R7042 a_41266_15922.n17 a_41266_15922.n16 0.536
R7043 a_41266_15922.n39 a_41266_15922.n38 0.255
R7044 a_41266_15922.n28 a_41266_15922.n27 0.151
R7045 a_41266_15922.n20 a_41266_15922.n19 0.151
R7046 a_41266_15922.n23 a_41266_15922.n22 0.125
R7047 a_41266_15922.n34 a_41266_15922.n32 0.028
R7048 a_41266_15922.n7 a_41266_15922.n5 0.028
R7049 a_41266_15922.n1 a_41266_15922.n0 0.025
R7050 a_41266_15922.n20 a_41266_15922.n15 0.024
R7051 a_41266_15922.n36 a_41266_15922.n34 0.012
R7052 a_41266_15922.n9 a_41266_15922.n7 0.012
R7053 a_41266_15922.n29 a_41266_15922.n23 0.011
R7054 a_41266_15922.n30 a_41266_15922.n29 0.011
R7055 a_41266_15922.n14 a_41266_15922.n10 0.011
R7056 a_41266_15922.n38 a_41266_15922.n37 0.01
R7057 a_41266_15922.n22 a_41266_15922.n21 0.01
R7058 a_41266_15922.n21 a_41266_15922.n14 0.01
R7059 a_41266_15922.n37 a_41266_15922.n30 0.01
R7060 a_32066_55442.n26 a_32066_55442.t2 10.181
R7061 a_32066_55442.n18 a_32066_55442.t1 10.181
R7062 a_32066_55442.t0 a_32066_55442.n39 9.68
R7063 a_32066_55442.n3 a_32066_55442.n2 9.302
R7064 a_32066_55442.n13 a_32066_55442.n12 9.302
R7065 a_32066_55442.n32 a_32066_55442.n31 9.3
R7066 a_32066_55442.n34 a_32066_55442.n33 9.3
R7067 a_32066_55442.n7 a_32066_55442.n6 9.3
R7068 a_32066_55442.n5 a_32066_55442.n4 9.3
R7069 a_32066_55442.n36 a_32066_55442.n35 9
R7070 a_32066_55442.n9 a_32066_55442.n8 9
R7071 a_32066_55442.n27 a_32066_55442.n25 7.729
R7072 a_32066_55442.n19 a_32066_55442.n17 7.729
R7073 a_32066_55442.n27 a_32066_55442.n26 6.296
R7074 a_32066_55442.n19 a_32066_55442.n18 6.296
R7075 a_32066_55442.n30 a_32066_55442.n3 4.508
R7076 a_32066_55442.n14 a_32066_55442.n13 4.508
R7077 a_32066_55442.n37 a_32066_55442.n36 4.496
R7078 a_32066_55442.n21 a_32066_55442.n20 4.496
R7079 a_32066_55442.n29 a_32066_55442.n28 4.495
R7080 a_32066_55442.n10 a_32066_55442.n9 4.495
R7081 a_32066_55442.n14 a_32066_55442.n11 4.494
R7082 a_32066_55442.n30 a_32066_55442.n1 4.494
R7083 a_32066_55442.n39 a_32066_55442.t3 1.087
R7084 a_32066_55442.n25 a_32066_55442.n24 0.536
R7085 a_32066_55442.n17 a_32066_55442.n16 0.536
R7086 a_32066_55442.n39 a_32066_55442.n38 0.255
R7087 a_32066_55442.n28 a_32066_55442.n27 0.151
R7088 a_32066_55442.n20 a_32066_55442.n19 0.151
R7089 a_32066_55442.n23 a_32066_55442.n22 0.125
R7090 a_32066_55442.n34 a_32066_55442.n32 0.028
R7091 a_32066_55442.n7 a_32066_55442.n5 0.028
R7092 a_32066_55442.n1 a_32066_55442.n0 0.025
R7093 a_32066_55442.n20 a_32066_55442.n15 0.024
R7094 a_32066_55442.n36 a_32066_55442.n34 0.012
R7095 a_32066_55442.n9 a_32066_55442.n7 0.012
R7096 a_32066_55442.n29 a_32066_55442.n23 0.011
R7097 a_32066_55442.n30 a_32066_55442.n29 0.011
R7098 a_32066_55442.n14 a_32066_55442.n10 0.011
R7099 a_32066_55442.n38 a_32066_55442.n37 0.01
R7100 a_32066_55442.n22 a_32066_55442.n21 0.01
R7101 a_32066_55442.n21 a_32066_55442.n14 0.01
R7102 a_32066_55442.n37 a_32066_55442.n30 0.01
R7103 a_31776_55366.n10 a_31776_55366.t0 10.181
R7104 a_31776_55366.n10 a_31776_55366.t1 10.181
R7105 a_31776_55366.t2 a_31776_55366.n18 9.68
R7106 a_31776_55366.n1 a_31776_55366.n0 9.302
R7107 a_31776_55366.n7 a_31776_55366.n6 9.3
R7108 a_31776_55366.n5 a_31776_55366.n4 9.3
R7109 a_31776_55366.n9 a_31776_55366.n8 9
R7110 a_31776_55366.n13 a_31776_55366.n12 7.729
R7111 a_31776_55366.n13 a_31776_55366.n10 6.296
R7112 a_31776_55366.n16 a_31776_55366.n1 4.508
R7113 a_31776_55366.n15 a_31776_55366.n14 4.501
R7114 a_31776_55366.n15 a_31776_55366.n9 4.501
R7115 a_31776_55366.n16 a_31776_55366.n3 4.494
R7116 a_31776_55366.n18 a_31776_55366.t3 1.259
R7117 a_31776_55366.n12 a_31776_55366.n11 0.536
R7118 a_31776_55366.n18 a_31776_55366.n17 0.415
R7119 a_31776_55366.n14 a_31776_55366.n13 0.151
R7120 a_31776_55366.n7 a_31776_55366.n5 0.028
R7121 a_31776_55366.n3 a_31776_55366.n2 0.025
R7122 a_31776_55366.n17 a_31776_55366.n16 0.021
R7123 a_31776_55366.n9 a_31776_55366.n7 0.012
R7124 a_31776_55366.n16 a_31776_55366.n15 0.006
R7125 a_4466_65322.n26 a_4466_65322.t0 10.181
R7126 a_4466_65322.n18 a_4466_65322.t3 10.181
R7127 a_4466_65322.t1 a_4466_65322.n39 9.68
R7128 a_4466_65322.n3 a_4466_65322.n2 9.302
R7129 a_4466_65322.n13 a_4466_65322.n12 9.302
R7130 a_4466_65322.n32 a_4466_65322.n31 9.3
R7131 a_4466_65322.n34 a_4466_65322.n33 9.3
R7132 a_4466_65322.n7 a_4466_65322.n6 9.3
R7133 a_4466_65322.n5 a_4466_65322.n4 9.3
R7134 a_4466_65322.n36 a_4466_65322.n35 9
R7135 a_4466_65322.n9 a_4466_65322.n8 9
R7136 a_4466_65322.n27 a_4466_65322.n25 7.729
R7137 a_4466_65322.n19 a_4466_65322.n17 7.729
R7138 a_4466_65322.n27 a_4466_65322.n26 6.296
R7139 a_4466_65322.n19 a_4466_65322.n18 6.296
R7140 a_4466_65322.n30 a_4466_65322.n3 4.508
R7141 a_4466_65322.n14 a_4466_65322.n13 4.508
R7142 a_4466_65322.n37 a_4466_65322.n36 4.496
R7143 a_4466_65322.n21 a_4466_65322.n20 4.496
R7144 a_4466_65322.n29 a_4466_65322.n28 4.495
R7145 a_4466_65322.n10 a_4466_65322.n9 4.495
R7146 a_4466_65322.n14 a_4466_65322.n11 4.494
R7147 a_4466_65322.n30 a_4466_65322.n1 4.494
R7148 a_4466_65322.n39 a_4466_65322.t2 1.087
R7149 a_4466_65322.n25 a_4466_65322.n24 0.536
R7150 a_4466_65322.n17 a_4466_65322.n16 0.536
R7151 a_4466_65322.n39 a_4466_65322.n38 0.255
R7152 a_4466_65322.n28 a_4466_65322.n27 0.151
R7153 a_4466_65322.n20 a_4466_65322.n19 0.151
R7154 a_4466_65322.n23 a_4466_65322.n22 0.125
R7155 a_4466_65322.n34 a_4466_65322.n32 0.028
R7156 a_4466_65322.n7 a_4466_65322.n5 0.028
R7157 a_4466_65322.n1 a_4466_65322.n0 0.025
R7158 a_4466_65322.n20 a_4466_65322.n15 0.024
R7159 a_4466_65322.n36 a_4466_65322.n34 0.012
R7160 a_4466_65322.n9 a_4466_65322.n7 0.012
R7161 a_4466_65322.n29 a_4466_65322.n23 0.011
R7162 a_4466_65322.n30 a_4466_65322.n29 0.011
R7163 a_4466_65322.n14 a_4466_65322.n10 0.011
R7164 a_4466_65322.n38 a_4466_65322.n37 0.01
R7165 a_4466_65322.n22 a_4466_65322.n21 0.01
R7166 a_4466_65322.n21 a_4466_65322.n14 0.01
R7167 a_4466_65322.n37 a_4466_65322.n30 0.01
R7168 a_n436_64726.t2 a_n436_64726.n15 139.026
R7169 a_n436_64726.n15 a_n436_64726.t9 85.389
R7170 a_n436_64726.n15 a_n436_64726.n14 54.371
R7171 a_n436_64726.n0 a_n436_64726.t7 9.633
R7172 a_n436_64726.n14 a_n436_64726.t3 9.587
R7173 a_n436_64726.n13 a_n436_64726.t5 9.587
R7174 a_n436_64726.n12 a_n436_64726.t8 9.587
R7175 a_n436_64726.n11 a_n436_64726.t4 9.587
R7176 a_n436_64726.n10 a_n436_64726.t10 9.587
R7177 a_n436_64726.n9 a_n436_64726.t13 9.587
R7178 a_n436_64726.n8 a_n436_64726.t12 9.587
R7179 a_n436_64726.n7 a_n436_64726.t14 9.587
R7180 a_n436_64726.n6 a_n436_64726.t6 9.587
R7181 a_n436_64726.n5 a_n436_64726.t1 9.587
R7182 a_n436_64726.n4 a_n436_64726.t11 9.587
R7183 a_n436_64726.n3 a_n436_64726.t15 9.587
R7184 a_n436_64726.n2 a_n436_64726.t16 9.587
R7185 a_n436_64726.n1 a_n436_64726.t0 9.587
R7186 a_n436_64726.n0 a_n436_64726.t17 9.587
R7187 a_n436_64726.n1 a_n436_64726.n0 0.528
R7188 a_n436_64726.n3 a_n436_64726.n2 0.528
R7189 a_n436_64726.n5 a_n436_64726.n4 0.528
R7190 a_n436_64726.n7 a_n436_64726.n6 0.528
R7191 a_n436_64726.n9 a_n436_64726.n8 0.528
R7192 a_n436_64726.n11 a_n436_64726.n10 0.528
R7193 a_n436_64726.n13 a_n436_64726.n12 0.528
R7194 a_n436_64726.n2 a_n436_64726.n1 0.046
R7195 a_n436_64726.n4 a_n436_64726.n3 0.046
R7196 a_n436_64726.n6 a_n436_64726.n5 0.046
R7197 a_n436_64726.n8 a_n436_64726.n7 0.046
R7198 a_n436_64726.n10 a_n436_64726.n9 0.046
R7199 a_n436_64726.n12 a_n436_64726.n11 0.046
R7200 a_n436_64726.n14 a_n436_64726.n13 0.046
R7201 a_22576_55366.n10 a_22576_55366.t0 10.181
R7202 a_22576_55366.n10 a_22576_55366.t1 10.181
R7203 a_22576_55366.t2 a_22576_55366.n18 9.68
R7204 a_22576_55366.n1 a_22576_55366.n0 9.302
R7205 a_22576_55366.n7 a_22576_55366.n6 9.3
R7206 a_22576_55366.n5 a_22576_55366.n4 9.3
R7207 a_22576_55366.n9 a_22576_55366.n8 9
R7208 a_22576_55366.n13 a_22576_55366.n12 7.729
R7209 a_22576_55366.n13 a_22576_55366.n10 6.296
R7210 a_22576_55366.n16 a_22576_55366.n1 4.508
R7211 a_22576_55366.n15 a_22576_55366.n14 4.501
R7212 a_22576_55366.n15 a_22576_55366.n9 4.501
R7213 a_22576_55366.n16 a_22576_55366.n3 4.494
R7214 a_22576_55366.n18 a_22576_55366.t3 1.259
R7215 a_22576_55366.n12 a_22576_55366.n11 0.536
R7216 a_22576_55366.n18 a_22576_55366.n17 0.415
R7217 a_22576_55366.n14 a_22576_55366.n13 0.151
R7218 a_22576_55366.n7 a_22576_55366.n5 0.028
R7219 a_22576_55366.n3 a_22576_55366.n2 0.025
R7220 a_22576_55366.n17 a_22576_55366.n16 0.021
R7221 a_22576_55366.n9 a_22576_55366.n7 0.012
R7222 a_22576_55366.n16 a_22576_55366.n15 0.006
R7223 a_50466_65322.n26 a_50466_65322.t0 10.181
R7224 a_50466_65322.n18 a_50466_65322.t2 10.181
R7225 a_50466_65322.t3 a_50466_65322.n39 9.68
R7226 a_50466_65322.n3 a_50466_65322.n2 9.302
R7227 a_50466_65322.n13 a_50466_65322.n12 9.302
R7228 a_50466_65322.n32 a_50466_65322.n31 9.3
R7229 a_50466_65322.n34 a_50466_65322.n33 9.3
R7230 a_50466_65322.n7 a_50466_65322.n6 9.3
R7231 a_50466_65322.n5 a_50466_65322.n4 9.3
R7232 a_50466_65322.n36 a_50466_65322.n35 9
R7233 a_50466_65322.n9 a_50466_65322.n8 9
R7234 a_50466_65322.n27 a_50466_65322.n25 7.729
R7235 a_50466_65322.n19 a_50466_65322.n17 7.729
R7236 a_50466_65322.n27 a_50466_65322.n26 6.296
R7237 a_50466_65322.n19 a_50466_65322.n18 6.296
R7238 a_50466_65322.n30 a_50466_65322.n3 4.508
R7239 a_50466_65322.n14 a_50466_65322.n13 4.508
R7240 a_50466_65322.n37 a_50466_65322.n36 4.496
R7241 a_50466_65322.n21 a_50466_65322.n20 4.496
R7242 a_50466_65322.n29 a_50466_65322.n28 4.495
R7243 a_50466_65322.n10 a_50466_65322.n9 4.495
R7244 a_50466_65322.n14 a_50466_65322.n11 4.494
R7245 a_50466_65322.n30 a_50466_65322.n1 4.494
R7246 a_50466_65322.n39 a_50466_65322.t1 1.087
R7247 a_50466_65322.n25 a_50466_65322.n24 0.536
R7248 a_50466_65322.n17 a_50466_65322.n16 0.536
R7249 a_50466_65322.n39 a_50466_65322.n38 0.255
R7250 a_50466_65322.n28 a_50466_65322.n27 0.151
R7251 a_50466_65322.n20 a_50466_65322.n19 0.151
R7252 a_50466_65322.n23 a_50466_65322.n22 0.125
R7253 a_50466_65322.n34 a_50466_65322.n32 0.028
R7254 a_50466_65322.n7 a_50466_65322.n5 0.028
R7255 a_50466_65322.n1 a_50466_65322.n0 0.025
R7256 a_50466_65322.n20 a_50466_65322.n15 0.024
R7257 a_50466_65322.n36 a_50466_65322.n34 0.012
R7258 a_50466_65322.n9 a_50466_65322.n7 0.012
R7259 a_50466_65322.n29 a_50466_65322.n23 0.011
R7260 a_50466_65322.n30 a_50466_65322.n29 0.011
R7261 a_50466_65322.n14 a_50466_65322.n10 0.011
R7262 a_50466_65322.n38 a_50466_65322.n37 0.01
R7263 a_50466_65322.n22 a_50466_65322.n21 0.01
R7264 a_50466_65322.n21 a_50466_65322.n14 0.01
R7265 a_50466_65322.n37 a_50466_65322.n30 0.01
R7266 a_4466_55442.n26 a_4466_55442.t0 10.181
R7267 a_4466_55442.n18 a_4466_55442.t1 10.181
R7268 a_4466_55442.t3 a_4466_55442.n39 9.68
R7269 a_4466_55442.n3 a_4466_55442.n2 9.302
R7270 a_4466_55442.n13 a_4466_55442.n12 9.302
R7271 a_4466_55442.n32 a_4466_55442.n31 9.3
R7272 a_4466_55442.n34 a_4466_55442.n33 9.3
R7273 a_4466_55442.n7 a_4466_55442.n6 9.3
R7274 a_4466_55442.n5 a_4466_55442.n4 9.3
R7275 a_4466_55442.n36 a_4466_55442.n35 9
R7276 a_4466_55442.n9 a_4466_55442.n8 9
R7277 a_4466_55442.n27 a_4466_55442.n25 7.729
R7278 a_4466_55442.n19 a_4466_55442.n17 7.729
R7279 a_4466_55442.n27 a_4466_55442.n26 6.296
R7280 a_4466_55442.n19 a_4466_55442.n18 6.296
R7281 a_4466_55442.n30 a_4466_55442.n3 4.508
R7282 a_4466_55442.n14 a_4466_55442.n13 4.508
R7283 a_4466_55442.n37 a_4466_55442.n36 4.496
R7284 a_4466_55442.n21 a_4466_55442.n20 4.496
R7285 a_4466_55442.n29 a_4466_55442.n28 4.495
R7286 a_4466_55442.n10 a_4466_55442.n9 4.495
R7287 a_4466_55442.n14 a_4466_55442.n11 4.494
R7288 a_4466_55442.n30 a_4466_55442.n1 4.494
R7289 a_4466_55442.n39 a_4466_55442.t2 1.087
R7290 a_4466_55442.n25 a_4466_55442.n24 0.536
R7291 a_4466_55442.n17 a_4466_55442.n16 0.536
R7292 a_4466_55442.n39 a_4466_55442.n38 0.255
R7293 a_4466_55442.n28 a_4466_55442.n27 0.151
R7294 a_4466_55442.n20 a_4466_55442.n19 0.151
R7295 a_4466_55442.n23 a_4466_55442.n22 0.125
R7296 a_4466_55442.n34 a_4466_55442.n32 0.028
R7297 a_4466_55442.n7 a_4466_55442.n5 0.028
R7298 a_4466_55442.n1 a_4466_55442.n0 0.025
R7299 a_4466_55442.n20 a_4466_55442.n15 0.024
R7300 a_4466_55442.n36 a_4466_55442.n34 0.012
R7301 a_4466_55442.n9 a_4466_55442.n7 0.012
R7302 a_4466_55442.n29 a_4466_55442.n23 0.011
R7303 a_4466_55442.n30 a_4466_55442.n29 0.011
R7304 a_4466_55442.n14 a_4466_55442.n10 0.011
R7305 a_4466_55442.n38 a_4466_55442.n37 0.01
R7306 a_4466_55442.n22 a_4466_55442.n21 0.01
R7307 a_4466_55442.n21 a_4466_55442.n14 0.01
R7308 a_4466_55442.n37 a_4466_55442.n30 0.01
R7309 a_4466_35682.n26 a_4466_35682.t0 10.181
R7310 a_4466_35682.n18 a_4466_35682.t1 10.181
R7311 a_4466_35682.t2 a_4466_35682.n39 9.68
R7312 a_4466_35682.n3 a_4466_35682.n2 9.302
R7313 a_4466_35682.n13 a_4466_35682.n12 9.302
R7314 a_4466_35682.n32 a_4466_35682.n31 9.3
R7315 a_4466_35682.n34 a_4466_35682.n33 9.3
R7316 a_4466_35682.n7 a_4466_35682.n6 9.3
R7317 a_4466_35682.n5 a_4466_35682.n4 9.3
R7318 a_4466_35682.n36 a_4466_35682.n35 9
R7319 a_4466_35682.n9 a_4466_35682.n8 9
R7320 a_4466_35682.n27 a_4466_35682.n25 7.729
R7321 a_4466_35682.n19 a_4466_35682.n17 7.729
R7322 a_4466_35682.n27 a_4466_35682.n26 6.296
R7323 a_4466_35682.n19 a_4466_35682.n18 6.296
R7324 a_4466_35682.n30 a_4466_35682.n3 4.508
R7325 a_4466_35682.n14 a_4466_35682.n13 4.508
R7326 a_4466_35682.n37 a_4466_35682.n36 4.496
R7327 a_4466_35682.n21 a_4466_35682.n20 4.496
R7328 a_4466_35682.n29 a_4466_35682.n28 4.495
R7329 a_4466_35682.n10 a_4466_35682.n9 4.495
R7330 a_4466_35682.n14 a_4466_35682.n11 4.494
R7331 a_4466_35682.n30 a_4466_35682.n1 4.494
R7332 a_4466_35682.n39 a_4466_35682.t3 1.087
R7333 a_4466_35682.n25 a_4466_35682.n24 0.536
R7334 a_4466_35682.n17 a_4466_35682.n16 0.536
R7335 a_4466_35682.n39 a_4466_35682.n38 0.255
R7336 a_4466_35682.n28 a_4466_35682.n27 0.151
R7337 a_4466_35682.n20 a_4466_35682.n19 0.151
R7338 a_4466_35682.n23 a_4466_35682.n22 0.125
R7339 a_4466_35682.n34 a_4466_35682.n32 0.028
R7340 a_4466_35682.n7 a_4466_35682.n5 0.028
R7341 a_4466_35682.n1 a_4466_35682.n0 0.025
R7342 a_4466_35682.n20 a_4466_35682.n15 0.024
R7343 a_4466_35682.n36 a_4466_35682.n34 0.012
R7344 a_4466_35682.n9 a_4466_35682.n7 0.012
R7345 a_4466_35682.n29 a_4466_35682.n23 0.011
R7346 a_4466_35682.n30 a_4466_35682.n29 0.011
R7347 a_4466_35682.n14 a_4466_35682.n10 0.011
R7348 a_4466_35682.n38 a_4466_35682.n37 0.01
R7349 a_4466_35682.n22 a_4466_35682.n21 0.01
R7350 a_4466_35682.n21 a_4466_35682.n14 0.01
R7351 a_4466_35682.n37 a_4466_35682.n30 0.01
R7352 a_4176_35606.n10 a_4176_35606.t0 10.181
R7353 a_4176_35606.n10 a_4176_35606.t1 10.181
R7354 a_4176_35606.t3 a_4176_35606.n18 9.68
R7355 a_4176_35606.n1 a_4176_35606.n0 9.302
R7356 a_4176_35606.n7 a_4176_35606.n6 9.3
R7357 a_4176_35606.n5 a_4176_35606.n4 9.3
R7358 a_4176_35606.n9 a_4176_35606.n8 9
R7359 a_4176_35606.n13 a_4176_35606.n12 7.729
R7360 a_4176_35606.n13 a_4176_35606.n10 6.296
R7361 a_4176_35606.n16 a_4176_35606.n1 4.508
R7362 a_4176_35606.n15 a_4176_35606.n14 4.501
R7363 a_4176_35606.n15 a_4176_35606.n9 4.501
R7364 a_4176_35606.n16 a_4176_35606.n3 4.494
R7365 a_4176_35606.n18 a_4176_35606.t2 1.259
R7366 a_4176_35606.n12 a_4176_35606.n11 0.536
R7367 a_4176_35606.n18 a_4176_35606.n17 0.415
R7368 a_4176_35606.n14 a_4176_35606.n13 0.151
R7369 a_4176_35606.n7 a_4176_35606.n5 0.028
R7370 a_4176_35606.n3 a_4176_35606.n2 0.025
R7371 a_4176_35606.n17 a_4176_35606.n16 0.021
R7372 a_4176_35606.n9 a_4176_35606.n7 0.012
R7373 a_4176_35606.n16 a_4176_35606.n15 0.006
R7374 a_22576_25726.n10 a_22576_25726.t1 10.181
R7375 a_22576_25726.n10 a_22576_25726.t0 10.181
R7376 a_22576_25726.t3 a_22576_25726.n18 9.68
R7377 a_22576_25726.n1 a_22576_25726.n0 9.302
R7378 a_22576_25726.n7 a_22576_25726.n6 9.3
R7379 a_22576_25726.n5 a_22576_25726.n4 9.3
R7380 a_22576_25726.n9 a_22576_25726.n8 9
R7381 a_22576_25726.n13 a_22576_25726.n12 7.729
R7382 a_22576_25726.n13 a_22576_25726.n10 6.296
R7383 a_22576_25726.n16 a_22576_25726.n1 4.508
R7384 a_22576_25726.n15 a_22576_25726.n14 4.501
R7385 a_22576_25726.n15 a_22576_25726.n9 4.501
R7386 a_22576_25726.n16 a_22576_25726.n3 4.494
R7387 a_22576_25726.n18 a_22576_25726.t2 1.259
R7388 a_22576_25726.n12 a_22576_25726.n11 0.536
R7389 a_22576_25726.n18 a_22576_25726.n17 0.415
R7390 a_22576_25726.n14 a_22576_25726.n13 0.151
R7391 a_22576_25726.n7 a_22576_25726.n5 0.028
R7392 a_22576_25726.n3 a_22576_25726.n2 0.025
R7393 a_22576_25726.n17 a_22576_25726.n16 0.021
R7394 a_22576_25726.n9 a_22576_25726.n7 0.012
R7395 a_22576_25726.n16 a_22576_25726.n15 0.006
R7396 a_22866_25802.n26 a_22866_25802.t2 10.181
R7397 a_22866_25802.n18 a_22866_25802.t1 10.181
R7398 a_22866_25802.t0 a_22866_25802.n39 9.68
R7399 a_22866_25802.n3 a_22866_25802.n2 9.302
R7400 a_22866_25802.n13 a_22866_25802.n12 9.302
R7401 a_22866_25802.n32 a_22866_25802.n31 9.3
R7402 a_22866_25802.n34 a_22866_25802.n33 9.3
R7403 a_22866_25802.n7 a_22866_25802.n6 9.3
R7404 a_22866_25802.n5 a_22866_25802.n4 9.3
R7405 a_22866_25802.n36 a_22866_25802.n35 9
R7406 a_22866_25802.n9 a_22866_25802.n8 9
R7407 a_22866_25802.n27 a_22866_25802.n25 7.729
R7408 a_22866_25802.n19 a_22866_25802.n17 7.729
R7409 a_22866_25802.n27 a_22866_25802.n26 6.296
R7410 a_22866_25802.n19 a_22866_25802.n18 6.296
R7411 a_22866_25802.n30 a_22866_25802.n3 4.508
R7412 a_22866_25802.n14 a_22866_25802.n13 4.508
R7413 a_22866_25802.n37 a_22866_25802.n36 4.496
R7414 a_22866_25802.n21 a_22866_25802.n20 4.496
R7415 a_22866_25802.n29 a_22866_25802.n28 4.495
R7416 a_22866_25802.n10 a_22866_25802.n9 4.495
R7417 a_22866_25802.n14 a_22866_25802.n11 4.494
R7418 a_22866_25802.n30 a_22866_25802.n1 4.494
R7419 a_22866_25802.n39 a_22866_25802.t3 1.087
R7420 a_22866_25802.n25 a_22866_25802.n24 0.536
R7421 a_22866_25802.n17 a_22866_25802.n16 0.536
R7422 a_22866_25802.n39 a_22866_25802.n38 0.255
R7423 a_22866_25802.n28 a_22866_25802.n27 0.151
R7424 a_22866_25802.n20 a_22866_25802.n19 0.151
R7425 a_22866_25802.n23 a_22866_25802.n22 0.125
R7426 a_22866_25802.n34 a_22866_25802.n32 0.028
R7427 a_22866_25802.n7 a_22866_25802.n5 0.028
R7428 a_22866_25802.n1 a_22866_25802.n0 0.025
R7429 a_22866_25802.n20 a_22866_25802.n15 0.024
R7430 a_22866_25802.n36 a_22866_25802.n34 0.012
R7431 a_22866_25802.n9 a_22866_25802.n7 0.012
R7432 a_22866_25802.n29 a_22866_25802.n23 0.011
R7433 a_22866_25802.n30 a_22866_25802.n29 0.011
R7434 a_22866_25802.n14 a_22866_25802.n10 0.011
R7435 a_22866_25802.n38 a_22866_25802.n37 0.01
R7436 a_22866_25802.n22 a_22866_25802.n21 0.01
R7437 a_22866_25802.n21 a_22866_25802.n14 0.01
R7438 a_22866_25802.n37 a_22866_25802.n30 0.01
R7439 bit2.n28 bit2.t9 552.693
R7440 bit2.n2 bit2.t7 300.446
R7441 bit2.n0 bit2.t2 300.446
R7442 bit2.n9 bit2.t6 300.446
R7443 bit2.n7 bit2.t4 300.446
R7444 bit2.n16 bit2.t8 300.446
R7445 bit2.n14 bit2.t3 300.446
R7446 bit2.n25 bit2.t0 300.446
R7447 bit2.n23 bit2.t5 300.446
R7448 bit2.n28 bit2.t1 279.56
R7449 bit2.n29 bit2.n28 120.317
R7450 bit2.n24 bit2.n23 27.537
R7451 bit2.n5 bit2.n2 27.536
R7452 bit2.n12 bit2.n9 27.536
R7453 bit2.n19 bit2.n16 27.536
R7454 bit2.n1 bit2.n0 24.127
R7455 bit2.n8 bit2.n7 24.127
R7456 bit2.n15 bit2.n14 24.127
R7457 bit2.n26 bit2.n25 24.127
R7458 bit2.n4 bit2.n3 8.764
R7459 bit2.n11 bit2.n10 8.764
R7460 bit2.n18 bit2.n17 8.764
R7461 bit2.n22 bit2.n21 8.764
R7462 bit2.n6 bit2.n1 4.662
R7463 bit2.n13 bit2.n8 4.662
R7464 bit2.n20 bit2.n15 4.662
R7465 bit2.n27 bit2.n26 4.661
R7466 bit2.n5 bit2.n4 3.401
R7467 bit2.n12 bit2.n11 3.401
R7468 bit2.n19 bit2.n18 3.401
R7469 bit2.n24 bit2.n22 3.401
R7470 bit2 bit2.n32 3.151
R7471 bit2.n27 bit2.n24 0.626
R7472 bit2.n6 bit2.n5 0.626
R7473 bit2.n13 bit2.n12 0.626
R7474 bit2.n20 bit2.n19 0.626
R7475 bit2.n32 bit2.n31 0.575
R7476 bit2.n31 bit2.n30 0.575
R7477 bit2.n30 bit2.n29 0.575
R7478 bit2.n32 bit2.n6 0.298
R7479 bit2.n31 bit2.n13 0.298
R7480 bit2.n30 bit2.n20 0.298
R7481 bit2.n29 bit2.n27 0.298
R7482 a_4176_75126.n10 a_4176_75126.t1 10.181
R7483 a_4176_75126.n10 a_4176_75126.t0 10.181
R7484 a_4176_75126.t3 a_4176_75126.n18 9.68
R7485 a_4176_75126.n1 a_4176_75126.n0 9.302
R7486 a_4176_75126.n7 a_4176_75126.n6 9.3
R7487 a_4176_75126.n5 a_4176_75126.n4 9.3
R7488 a_4176_75126.n9 a_4176_75126.n8 9
R7489 a_4176_75126.n13 a_4176_75126.n12 7.729
R7490 a_4176_75126.n13 a_4176_75126.n10 6.296
R7491 a_4176_75126.n16 a_4176_75126.n1 4.508
R7492 a_4176_75126.n15 a_4176_75126.n14 4.501
R7493 a_4176_75126.n15 a_4176_75126.n9 4.501
R7494 a_4176_75126.n16 a_4176_75126.n3 4.494
R7495 a_4176_75126.n18 a_4176_75126.t2 1.259
R7496 a_4176_75126.n12 a_4176_75126.n11 0.536
R7497 a_4176_75126.n18 a_4176_75126.n17 0.415
R7498 a_4176_75126.n14 a_4176_75126.n13 0.151
R7499 a_4176_75126.n7 a_4176_75126.n5 0.028
R7500 a_4176_75126.n3 a_4176_75126.n2 0.025
R7501 a_4176_75126.n17 a_4176_75126.n16 0.021
R7502 a_4176_75126.n9 a_4176_75126.n7 0.012
R7503 a_4176_75126.n16 a_4176_75126.n15 0.006
R7504 a_4466_75202.n26 a_4466_75202.t1 10.181
R7505 a_4466_75202.n18 a_4466_75202.t0 10.181
R7506 a_4466_75202.t3 a_4466_75202.n39 9.68
R7507 a_4466_75202.n3 a_4466_75202.n2 9.302
R7508 a_4466_75202.n13 a_4466_75202.n12 9.302
R7509 a_4466_75202.n32 a_4466_75202.n31 9.3
R7510 a_4466_75202.n34 a_4466_75202.n33 9.3
R7511 a_4466_75202.n7 a_4466_75202.n6 9.3
R7512 a_4466_75202.n5 a_4466_75202.n4 9.3
R7513 a_4466_75202.n36 a_4466_75202.n35 9
R7514 a_4466_75202.n9 a_4466_75202.n8 9
R7515 a_4466_75202.n27 a_4466_75202.n25 7.729
R7516 a_4466_75202.n19 a_4466_75202.n17 7.729
R7517 a_4466_75202.n27 a_4466_75202.n26 6.296
R7518 a_4466_75202.n19 a_4466_75202.n18 6.296
R7519 a_4466_75202.n30 a_4466_75202.n3 4.508
R7520 a_4466_75202.n14 a_4466_75202.n13 4.508
R7521 a_4466_75202.n37 a_4466_75202.n36 4.496
R7522 a_4466_75202.n21 a_4466_75202.n20 4.496
R7523 a_4466_75202.n29 a_4466_75202.n28 4.495
R7524 a_4466_75202.n10 a_4466_75202.n9 4.495
R7525 a_4466_75202.n14 a_4466_75202.n11 4.494
R7526 a_4466_75202.n30 a_4466_75202.n1 4.494
R7527 a_4466_75202.n39 a_4466_75202.t2 1.087
R7528 a_4466_75202.n25 a_4466_75202.n24 0.536
R7529 a_4466_75202.n17 a_4466_75202.n16 0.536
R7530 a_4466_75202.n39 a_4466_75202.n38 0.255
R7531 a_4466_75202.n28 a_4466_75202.n27 0.151
R7532 a_4466_75202.n20 a_4466_75202.n19 0.151
R7533 a_4466_75202.n23 a_4466_75202.n22 0.125
R7534 a_4466_75202.n34 a_4466_75202.n32 0.028
R7535 a_4466_75202.n7 a_4466_75202.n5 0.028
R7536 a_4466_75202.n1 a_4466_75202.n0 0.025
R7537 a_4466_75202.n20 a_4466_75202.n15 0.024
R7538 a_4466_75202.n36 a_4466_75202.n34 0.012
R7539 a_4466_75202.n9 a_4466_75202.n7 0.012
R7540 a_4466_75202.n29 a_4466_75202.n23 0.011
R7541 a_4466_75202.n30 a_4466_75202.n29 0.011
R7542 a_4466_75202.n14 a_4466_75202.n10 0.011
R7543 a_4466_75202.n38 a_4466_75202.n37 0.01
R7544 a_4466_75202.n22 a_4466_75202.n21 0.01
R7545 a_4466_75202.n21 a_4466_75202.n14 0.01
R7546 a_4466_75202.n37 a_4466_75202.n30 0.01
R7547 a_4466_94962.n26 a_4466_94962.t0 10.181
R7548 a_4466_94962.n18 a_4466_94962.t1 10.181
R7549 a_4466_94962.t3 a_4466_94962.n39 9.68
R7550 a_4466_94962.n3 a_4466_94962.n2 9.302
R7551 a_4466_94962.n13 a_4466_94962.n12 9.302
R7552 a_4466_94962.n32 a_4466_94962.n31 9.3
R7553 a_4466_94962.n34 a_4466_94962.n33 9.3
R7554 a_4466_94962.n7 a_4466_94962.n6 9.3
R7555 a_4466_94962.n5 a_4466_94962.n4 9.3
R7556 a_4466_94962.n36 a_4466_94962.n35 9
R7557 a_4466_94962.n9 a_4466_94962.n8 9
R7558 a_4466_94962.n27 a_4466_94962.n25 7.729
R7559 a_4466_94962.n19 a_4466_94962.n17 7.729
R7560 a_4466_94962.n27 a_4466_94962.n26 6.296
R7561 a_4466_94962.n19 a_4466_94962.n18 6.296
R7562 a_4466_94962.n30 a_4466_94962.n3 4.508
R7563 a_4466_94962.n14 a_4466_94962.n13 4.508
R7564 a_4466_94962.n37 a_4466_94962.n36 4.496
R7565 a_4466_94962.n21 a_4466_94962.n20 4.496
R7566 a_4466_94962.n29 a_4466_94962.n28 4.495
R7567 a_4466_94962.n10 a_4466_94962.n9 4.495
R7568 a_4466_94962.n14 a_4466_94962.n11 4.494
R7569 a_4466_94962.n30 a_4466_94962.n1 4.494
R7570 a_4466_94962.n39 a_4466_94962.t2 1.087
R7571 a_4466_94962.n25 a_4466_94962.n24 0.536
R7572 a_4466_94962.n17 a_4466_94962.n16 0.536
R7573 a_4466_94962.n39 a_4466_94962.n38 0.255
R7574 a_4466_94962.n28 a_4466_94962.n27 0.151
R7575 a_4466_94962.n20 a_4466_94962.n19 0.151
R7576 a_4466_94962.n23 a_4466_94962.n22 0.125
R7577 a_4466_94962.n34 a_4466_94962.n32 0.028
R7578 a_4466_94962.n7 a_4466_94962.n5 0.028
R7579 a_4466_94962.n1 a_4466_94962.n0 0.025
R7580 a_4466_94962.n20 a_4466_94962.n15 0.024
R7581 a_4466_94962.n36 a_4466_94962.n34 0.012
R7582 a_4466_94962.n9 a_4466_94962.n7 0.012
R7583 a_4466_94962.n29 a_4466_94962.n23 0.011
R7584 a_4466_94962.n30 a_4466_94962.n29 0.011
R7585 a_4466_94962.n14 a_4466_94962.n10 0.011
R7586 a_4466_94962.n38 a_4466_94962.n37 0.01
R7587 a_4466_94962.n22 a_4466_94962.n21 0.01
R7588 a_4466_94962.n21 a_4466_94962.n14 0.01
R7589 a_4466_94962.n37 a_4466_94962.n30 0.01
R7590 a_13376_65246.n10 a_13376_65246.t0 10.181
R7591 a_13376_65246.n10 a_13376_65246.t3 10.181
R7592 a_13376_65246.t1 a_13376_65246.n18 9.68
R7593 a_13376_65246.n1 a_13376_65246.n0 9.302
R7594 a_13376_65246.n7 a_13376_65246.n6 9.3
R7595 a_13376_65246.n5 a_13376_65246.n4 9.3
R7596 a_13376_65246.n9 a_13376_65246.n8 9
R7597 a_13376_65246.n13 a_13376_65246.n12 7.729
R7598 a_13376_65246.n13 a_13376_65246.n10 6.296
R7599 a_13376_65246.n16 a_13376_65246.n1 4.508
R7600 a_13376_65246.n15 a_13376_65246.n14 4.501
R7601 a_13376_65246.n15 a_13376_65246.n9 4.501
R7602 a_13376_65246.n16 a_13376_65246.n3 4.494
R7603 a_13376_65246.n18 a_13376_65246.t2 1.259
R7604 a_13376_65246.n12 a_13376_65246.n11 0.536
R7605 a_13376_65246.n18 a_13376_65246.n17 0.415
R7606 a_13376_65246.n14 a_13376_65246.n13 0.151
R7607 a_13376_65246.n7 a_13376_65246.n5 0.028
R7608 a_13376_65246.n3 a_13376_65246.n2 0.025
R7609 a_13376_65246.n17 a_13376_65246.n16 0.021
R7610 a_13376_65246.n9 a_13376_65246.n7 0.012
R7611 a_13376_65246.n16 a_13376_65246.n15 0.006
R7612 a_32066_45562.n26 a_32066_45562.t2 10.181
R7613 a_32066_45562.n18 a_32066_45562.t1 10.181
R7614 a_32066_45562.t0 a_32066_45562.n39 9.68
R7615 a_32066_45562.n3 a_32066_45562.n2 9.302
R7616 a_32066_45562.n13 a_32066_45562.n12 9.302
R7617 a_32066_45562.n32 a_32066_45562.n31 9.3
R7618 a_32066_45562.n34 a_32066_45562.n33 9.3
R7619 a_32066_45562.n7 a_32066_45562.n6 9.3
R7620 a_32066_45562.n5 a_32066_45562.n4 9.3
R7621 a_32066_45562.n36 a_32066_45562.n35 9
R7622 a_32066_45562.n9 a_32066_45562.n8 9
R7623 a_32066_45562.n27 a_32066_45562.n25 7.729
R7624 a_32066_45562.n19 a_32066_45562.n17 7.729
R7625 a_32066_45562.n27 a_32066_45562.n26 6.296
R7626 a_32066_45562.n19 a_32066_45562.n18 6.296
R7627 a_32066_45562.n30 a_32066_45562.n3 4.508
R7628 a_32066_45562.n14 a_32066_45562.n13 4.508
R7629 a_32066_45562.n37 a_32066_45562.n36 4.496
R7630 a_32066_45562.n21 a_32066_45562.n20 4.496
R7631 a_32066_45562.n29 a_32066_45562.n28 4.495
R7632 a_32066_45562.n10 a_32066_45562.n9 4.495
R7633 a_32066_45562.n14 a_32066_45562.n11 4.494
R7634 a_32066_45562.n30 a_32066_45562.n1 4.494
R7635 a_32066_45562.n39 a_32066_45562.t3 1.087
R7636 a_32066_45562.n25 a_32066_45562.n24 0.536
R7637 a_32066_45562.n17 a_32066_45562.n16 0.536
R7638 a_32066_45562.n39 a_32066_45562.n38 0.255
R7639 a_32066_45562.n28 a_32066_45562.n27 0.151
R7640 a_32066_45562.n20 a_32066_45562.n19 0.151
R7641 a_32066_45562.n23 a_32066_45562.n22 0.125
R7642 a_32066_45562.n34 a_32066_45562.n32 0.028
R7643 a_32066_45562.n7 a_32066_45562.n5 0.028
R7644 a_32066_45562.n1 a_32066_45562.n0 0.025
R7645 a_32066_45562.n20 a_32066_45562.n15 0.024
R7646 a_32066_45562.n36 a_32066_45562.n34 0.012
R7647 a_32066_45562.n9 a_32066_45562.n7 0.012
R7648 a_32066_45562.n29 a_32066_45562.n23 0.011
R7649 a_32066_45562.n30 a_32066_45562.n29 0.011
R7650 a_32066_45562.n14 a_32066_45562.n10 0.011
R7651 a_32066_45562.n38 a_32066_45562.n37 0.01
R7652 a_32066_45562.n22 a_32066_45562.n21 0.01
R7653 a_32066_45562.n21 a_32066_45562.n14 0.01
R7654 a_32066_45562.n37 a_32066_45562.n30 0.01
R7655 a_13666_55442.n26 a_13666_55442.t2 10.181
R7656 a_13666_55442.n18 a_13666_55442.t1 10.181
R7657 a_13666_55442.t0 a_13666_55442.n39 9.68
R7658 a_13666_55442.n3 a_13666_55442.n2 9.302
R7659 a_13666_55442.n13 a_13666_55442.n12 9.302
R7660 a_13666_55442.n32 a_13666_55442.n31 9.3
R7661 a_13666_55442.n34 a_13666_55442.n33 9.3
R7662 a_13666_55442.n7 a_13666_55442.n6 9.3
R7663 a_13666_55442.n5 a_13666_55442.n4 9.3
R7664 a_13666_55442.n36 a_13666_55442.n35 9
R7665 a_13666_55442.n9 a_13666_55442.n8 9
R7666 a_13666_55442.n27 a_13666_55442.n25 7.729
R7667 a_13666_55442.n19 a_13666_55442.n17 7.729
R7668 a_13666_55442.n27 a_13666_55442.n26 6.296
R7669 a_13666_55442.n19 a_13666_55442.n18 6.296
R7670 a_13666_55442.n30 a_13666_55442.n3 4.508
R7671 a_13666_55442.n14 a_13666_55442.n13 4.508
R7672 a_13666_55442.n37 a_13666_55442.n36 4.496
R7673 a_13666_55442.n21 a_13666_55442.n20 4.496
R7674 a_13666_55442.n29 a_13666_55442.n28 4.495
R7675 a_13666_55442.n10 a_13666_55442.n9 4.495
R7676 a_13666_55442.n14 a_13666_55442.n11 4.494
R7677 a_13666_55442.n30 a_13666_55442.n1 4.494
R7678 a_13666_55442.n39 a_13666_55442.t3 1.087
R7679 a_13666_55442.n25 a_13666_55442.n24 0.536
R7680 a_13666_55442.n17 a_13666_55442.n16 0.536
R7681 a_13666_55442.n39 a_13666_55442.n38 0.255
R7682 a_13666_55442.n28 a_13666_55442.n27 0.151
R7683 a_13666_55442.n20 a_13666_55442.n19 0.151
R7684 a_13666_55442.n23 a_13666_55442.n22 0.125
R7685 a_13666_55442.n34 a_13666_55442.n32 0.028
R7686 a_13666_55442.n7 a_13666_55442.n5 0.028
R7687 a_13666_55442.n1 a_13666_55442.n0 0.025
R7688 a_13666_55442.n20 a_13666_55442.n15 0.024
R7689 a_13666_55442.n36 a_13666_55442.n34 0.012
R7690 a_13666_55442.n9 a_13666_55442.n7 0.012
R7691 a_13666_55442.n29 a_13666_55442.n23 0.011
R7692 a_13666_55442.n30 a_13666_55442.n29 0.011
R7693 a_13666_55442.n14 a_13666_55442.n10 0.011
R7694 a_13666_55442.n38 a_13666_55442.n37 0.01
R7695 a_13666_55442.n22 a_13666_55442.n21 0.01
R7696 a_13666_55442.n21 a_13666_55442.n14 0.01
R7697 a_13666_55442.n37 a_13666_55442.n30 0.01
R7698 a_13376_55366.n10 a_13376_55366.t0 10.181
R7699 a_13376_55366.n10 a_13376_55366.t1 10.181
R7700 a_13376_55366.t2 a_13376_55366.n18 9.68
R7701 a_13376_55366.n1 a_13376_55366.n0 9.302
R7702 a_13376_55366.n7 a_13376_55366.n6 9.3
R7703 a_13376_55366.n5 a_13376_55366.n4 9.3
R7704 a_13376_55366.n9 a_13376_55366.n8 9
R7705 a_13376_55366.n13 a_13376_55366.n12 7.729
R7706 a_13376_55366.n13 a_13376_55366.n10 6.296
R7707 a_13376_55366.n16 a_13376_55366.n1 4.508
R7708 a_13376_55366.n15 a_13376_55366.n14 4.501
R7709 a_13376_55366.n15 a_13376_55366.n9 4.501
R7710 a_13376_55366.n16 a_13376_55366.n3 4.494
R7711 a_13376_55366.n18 a_13376_55366.t3 1.259
R7712 a_13376_55366.n12 a_13376_55366.n11 0.536
R7713 a_13376_55366.n18 a_13376_55366.n17 0.415
R7714 a_13376_55366.n14 a_13376_55366.n13 0.151
R7715 a_13376_55366.n7 a_13376_55366.n5 0.028
R7716 a_13376_55366.n3 a_13376_55366.n2 0.025
R7717 a_13376_55366.n17 a_13376_55366.n16 0.021
R7718 a_13376_55366.n9 a_13376_55366.n7 0.012
R7719 a_13376_55366.n16 a_13376_55366.n15 0.006
R7720 a_4466_6042.n26 a_4466_6042.t2 10.181
R7721 a_4466_6042.n18 a_4466_6042.t1 10.181
R7722 a_4466_6042.t0 a_4466_6042.n39 9.68
R7723 a_4466_6042.n3 a_4466_6042.n2 9.302
R7724 a_4466_6042.n13 a_4466_6042.n12 9.302
R7725 a_4466_6042.n32 a_4466_6042.n31 9.3
R7726 a_4466_6042.n34 a_4466_6042.n33 9.3
R7727 a_4466_6042.n7 a_4466_6042.n6 9.3
R7728 a_4466_6042.n5 a_4466_6042.n4 9.3
R7729 a_4466_6042.n36 a_4466_6042.n35 9
R7730 a_4466_6042.n9 a_4466_6042.n8 9
R7731 a_4466_6042.n27 a_4466_6042.n25 7.729
R7732 a_4466_6042.n19 a_4466_6042.n17 7.729
R7733 a_4466_6042.n27 a_4466_6042.n26 6.296
R7734 a_4466_6042.n19 a_4466_6042.n18 6.296
R7735 a_4466_6042.n30 a_4466_6042.n3 4.508
R7736 a_4466_6042.n14 a_4466_6042.n13 4.508
R7737 a_4466_6042.n37 a_4466_6042.n36 4.496
R7738 a_4466_6042.n21 a_4466_6042.n20 4.496
R7739 a_4466_6042.n29 a_4466_6042.n28 4.495
R7740 a_4466_6042.n10 a_4466_6042.n9 4.495
R7741 a_4466_6042.n14 a_4466_6042.n11 4.494
R7742 a_4466_6042.n30 a_4466_6042.n1 4.494
R7743 a_4466_6042.n39 a_4466_6042.t3 1.087
R7744 a_4466_6042.n25 a_4466_6042.n24 0.536
R7745 a_4466_6042.n17 a_4466_6042.n16 0.536
R7746 a_4466_6042.n39 a_4466_6042.n38 0.255
R7747 a_4466_6042.n28 a_4466_6042.n27 0.151
R7748 a_4466_6042.n20 a_4466_6042.n19 0.151
R7749 a_4466_6042.n23 a_4466_6042.n22 0.125
R7750 a_4466_6042.n34 a_4466_6042.n32 0.028
R7751 a_4466_6042.n7 a_4466_6042.n5 0.028
R7752 a_4466_6042.n1 a_4466_6042.n0 0.025
R7753 a_4466_6042.n20 a_4466_6042.n15 0.024
R7754 a_4466_6042.n36 a_4466_6042.n34 0.012
R7755 a_4466_6042.n9 a_4466_6042.n7 0.012
R7756 a_4466_6042.n29 a_4466_6042.n23 0.011
R7757 a_4466_6042.n30 a_4466_6042.n29 0.011
R7758 a_4466_6042.n14 a_4466_6042.n10 0.011
R7759 a_4466_6042.n38 a_4466_6042.n37 0.01
R7760 a_4466_6042.n22 a_4466_6042.n21 0.01
R7761 a_4466_6042.n21 a_4466_6042.n14 0.01
R7762 a_4466_6042.n37 a_4466_6042.n30 0.01
R7763 a_40976_25726.n10 a_40976_25726.t2 10.181
R7764 a_40976_25726.n10 a_40976_25726.t1 10.181
R7765 a_40976_25726.t0 a_40976_25726.n18 9.68
R7766 a_40976_25726.n1 a_40976_25726.n0 9.302
R7767 a_40976_25726.n7 a_40976_25726.n6 9.3
R7768 a_40976_25726.n5 a_40976_25726.n4 9.3
R7769 a_40976_25726.n9 a_40976_25726.n8 9
R7770 a_40976_25726.n13 a_40976_25726.n12 7.729
R7771 a_40976_25726.n13 a_40976_25726.n10 6.296
R7772 a_40976_25726.n16 a_40976_25726.n1 4.508
R7773 a_40976_25726.n15 a_40976_25726.n14 4.501
R7774 a_40976_25726.n15 a_40976_25726.n9 4.501
R7775 a_40976_25726.n16 a_40976_25726.n3 4.494
R7776 a_40976_25726.n18 a_40976_25726.t3 1.259
R7777 a_40976_25726.n12 a_40976_25726.n11 0.536
R7778 a_40976_25726.n18 a_40976_25726.n17 0.415
R7779 a_40976_25726.n14 a_40976_25726.n13 0.151
R7780 a_40976_25726.n7 a_40976_25726.n5 0.028
R7781 a_40976_25726.n3 a_40976_25726.n2 0.025
R7782 a_40976_25726.n17 a_40976_25726.n16 0.021
R7783 a_40976_25726.n9 a_40976_25726.n7 0.012
R7784 a_40976_25726.n16 a_40976_25726.n15 0.006
R7785 a_68576_35606.n10 a_68576_35606.t2 10.181
R7786 a_68576_35606.n10 a_68576_35606.t1 10.181
R7787 a_68576_35606.t0 a_68576_35606.n18 9.68
R7788 a_68576_35606.n1 a_68576_35606.n0 9.302
R7789 a_68576_35606.n7 a_68576_35606.n6 9.3
R7790 a_68576_35606.n5 a_68576_35606.n4 9.3
R7791 a_68576_35606.n9 a_68576_35606.n8 9
R7792 a_68576_35606.n13 a_68576_35606.n12 7.729
R7793 a_68576_35606.n13 a_68576_35606.n10 6.296
R7794 a_68576_35606.n16 a_68576_35606.n1 4.508
R7795 a_68576_35606.n15 a_68576_35606.n14 4.501
R7796 a_68576_35606.n15 a_68576_35606.n9 4.501
R7797 a_68576_35606.n16 a_68576_35606.n3 4.494
R7798 a_68576_35606.n18 a_68576_35606.t3 1.259
R7799 a_68576_35606.n12 a_68576_35606.n11 0.536
R7800 a_68576_35606.n18 a_68576_35606.n17 0.415
R7801 a_68576_35606.n14 a_68576_35606.n13 0.151
R7802 a_68576_35606.n7 a_68576_35606.n5 0.028
R7803 a_68576_35606.n3 a_68576_35606.n2 0.025
R7804 a_68576_35606.n17 a_68576_35606.n16 0.021
R7805 a_68576_35606.n9 a_68576_35606.n7 0.012
R7806 a_68576_35606.n16 a_68576_35606.n15 0.006
R7807 a_32066_6042.n26 a_32066_6042.t1 10.181
R7808 a_32066_6042.n18 a_32066_6042.t0 10.181
R7809 a_32066_6042.t2 a_32066_6042.n39 9.68
R7810 a_32066_6042.n3 a_32066_6042.n2 9.302
R7811 a_32066_6042.n13 a_32066_6042.n12 9.302
R7812 a_32066_6042.n32 a_32066_6042.n31 9.3
R7813 a_32066_6042.n34 a_32066_6042.n33 9.3
R7814 a_32066_6042.n7 a_32066_6042.n6 9.3
R7815 a_32066_6042.n5 a_32066_6042.n4 9.3
R7816 a_32066_6042.n36 a_32066_6042.n35 9
R7817 a_32066_6042.n9 a_32066_6042.n8 9
R7818 a_32066_6042.n27 a_32066_6042.n25 7.729
R7819 a_32066_6042.n19 a_32066_6042.n17 7.729
R7820 a_32066_6042.n27 a_32066_6042.n26 6.296
R7821 a_32066_6042.n19 a_32066_6042.n18 6.296
R7822 a_32066_6042.n30 a_32066_6042.n3 4.508
R7823 a_32066_6042.n14 a_32066_6042.n13 4.508
R7824 a_32066_6042.n37 a_32066_6042.n36 4.496
R7825 a_32066_6042.n21 a_32066_6042.n20 4.496
R7826 a_32066_6042.n29 a_32066_6042.n28 4.495
R7827 a_32066_6042.n10 a_32066_6042.n9 4.495
R7828 a_32066_6042.n14 a_32066_6042.n11 4.494
R7829 a_32066_6042.n30 a_32066_6042.n1 4.494
R7830 a_32066_6042.n39 a_32066_6042.t3 1.087
R7831 a_32066_6042.n25 a_32066_6042.n24 0.536
R7832 a_32066_6042.n17 a_32066_6042.n16 0.536
R7833 a_32066_6042.n39 a_32066_6042.n38 0.255
R7834 a_32066_6042.n28 a_32066_6042.n27 0.151
R7835 a_32066_6042.n20 a_32066_6042.n19 0.151
R7836 a_32066_6042.n23 a_32066_6042.n22 0.125
R7837 a_32066_6042.n34 a_32066_6042.n32 0.028
R7838 a_32066_6042.n7 a_32066_6042.n5 0.028
R7839 a_32066_6042.n1 a_32066_6042.n0 0.025
R7840 a_32066_6042.n20 a_32066_6042.n15 0.024
R7841 a_32066_6042.n36 a_32066_6042.n34 0.012
R7842 a_32066_6042.n9 a_32066_6042.n7 0.012
R7843 a_32066_6042.n29 a_32066_6042.n23 0.011
R7844 a_32066_6042.n30 a_32066_6042.n29 0.011
R7845 a_32066_6042.n14 a_32066_6042.n10 0.011
R7846 a_32066_6042.n38 a_32066_6042.n37 0.01
R7847 a_32066_6042.n22 a_32066_6042.n21 0.01
R7848 a_32066_6042.n21 a_32066_6042.n14 0.01
R7849 a_32066_6042.n37 a_32066_6042.n30 0.01
R7850 a_22866_55442.n26 a_22866_55442.t1 10.181
R7851 a_22866_55442.n18 a_22866_55442.t2 10.181
R7852 a_22866_55442.t0 a_22866_55442.n39 9.68
R7853 a_22866_55442.n3 a_22866_55442.n2 9.302
R7854 a_22866_55442.n13 a_22866_55442.n12 9.302
R7855 a_22866_55442.n32 a_22866_55442.n31 9.3
R7856 a_22866_55442.n34 a_22866_55442.n33 9.3
R7857 a_22866_55442.n7 a_22866_55442.n6 9.3
R7858 a_22866_55442.n5 a_22866_55442.n4 9.3
R7859 a_22866_55442.n36 a_22866_55442.n35 9
R7860 a_22866_55442.n9 a_22866_55442.n8 9
R7861 a_22866_55442.n27 a_22866_55442.n25 7.729
R7862 a_22866_55442.n19 a_22866_55442.n17 7.729
R7863 a_22866_55442.n27 a_22866_55442.n26 6.296
R7864 a_22866_55442.n19 a_22866_55442.n18 6.296
R7865 a_22866_55442.n30 a_22866_55442.n3 4.508
R7866 a_22866_55442.n14 a_22866_55442.n13 4.508
R7867 a_22866_55442.n37 a_22866_55442.n36 4.496
R7868 a_22866_55442.n21 a_22866_55442.n20 4.496
R7869 a_22866_55442.n29 a_22866_55442.n28 4.495
R7870 a_22866_55442.n10 a_22866_55442.n9 4.495
R7871 a_22866_55442.n14 a_22866_55442.n11 4.494
R7872 a_22866_55442.n30 a_22866_55442.n1 4.494
R7873 a_22866_55442.n39 a_22866_55442.t3 1.087
R7874 a_22866_55442.n25 a_22866_55442.n24 0.536
R7875 a_22866_55442.n17 a_22866_55442.n16 0.536
R7876 a_22866_55442.n39 a_22866_55442.n38 0.255
R7877 a_22866_55442.n28 a_22866_55442.n27 0.151
R7878 a_22866_55442.n20 a_22866_55442.n19 0.151
R7879 a_22866_55442.n23 a_22866_55442.n22 0.125
R7880 a_22866_55442.n34 a_22866_55442.n32 0.028
R7881 a_22866_55442.n7 a_22866_55442.n5 0.028
R7882 a_22866_55442.n1 a_22866_55442.n0 0.025
R7883 a_22866_55442.n20 a_22866_55442.n15 0.024
R7884 a_22866_55442.n36 a_22866_55442.n34 0.012
R7885 a_22866_55442.n9 a_22866_55442.n7 0.012
R7886 a_22866_55442.n29 a_22866_55442.n23 0.011
R7887 a_22866_55442.n30 a_22866_55442.n29 0.011
R7888 a_22866_55442.n14 a_22866_55442.n10 0.011
R7889 a_22866_55442.n38 a_22866_55442.n37 0.01
R7890 a_22866_55442.n22 a_22866_55442.n21 0.01
R7891 a_22866_55442.n21 a_22866_55442.n14 0.01
R7892 a_22866_55442.n37 a_22866_55442.n30 0.01
R7893 a_22576_35606.n10 a_22576_35606.t0 10.181
R7894 a_22576_35606.n10 a_22576_35606.t1 10.181
R7895 a_22576_35606.t2 a_22576_35606.n18 9.68
R7896 a_22576_35606.n1 a_22576_35606.n0 9.302
R7897 a_22576_35606.n7 a_22576_35606.n6 9.3
R7898 a_22576_35606.n5 a_22576_35606.n4 9.3
R7899 a_22576_35606.n9 a_22576_35606.n8 9
R7900 a_22576_35606.n13 a_22576_35606.n12 7.729
R7901 a_22576_35606.n13 a_22576_35606.n10 6.296
R7902 a_22576_35606.n16 a_22576_35606.n1 4.508
R7903 a_22576_35606.n15 a_22576_35606.n14 4.501
R7904 a_22576_35606.n15 a_22576_35606.n9 4.501
R7905 a_22576_35606.n16 a_22576_35606.n3 4.494
R7906 a_22576_35606.n18 a_22576_35606.t3 1.259
R7907 a_22576_35606.n12 a_22576_35606.n11 0.536
R7908 a_22576_35606.n18 a_22576_35606.n17 0.415
R7909 a_22576_35606.n14 a_22576_35606.n13 0.151
R7910 a_22576_35606.n7 a_22576_35606.n5 0.028
R7911 a_22576_35606.n3 a_22576_35606.n2 0.025
R7912 a_22576_35606.n17 a_22576_35606.n16 0.021
R7913 a_22576_35606.n9 a_22576_35606.n7 0.012
R7914 a_22576_35606.n16 a_22576_35606.n15 0.006
R7915 a_41266_55442.n26 a_41266_55442.t1 10.181
R7916 a_41266_55442.n18 a_41266_55442.t0 10.181
R7917 a_41266_55442.t3 a_41266_55442.n39 9.68
R7918 a_41266_55442.n3 a_41266_55442.n2 9.302
R7919 a_41266_55442.n13 a_41266_55442.n12 9.302
R7920 a_41266_55442.n32 a_41266_55442.n31 9.3
R7921 a_41266_55442.n34 a_41266_55442.n33 9.3
R7922 a_41266_55442.n7 a_41266_55442.n6 9.3
R7923 a_41266_55442.n5 a_41266_55442.n4 9.3
R7924 a_41266_55442.n36 a_41266_55442.n35 9
R7925 a_41266_55442.n9 a_41266_55442.n8 9
R7926 a_41266_55442.n27 a_41266_55442.n25 7.729
R7927 a_41266_55442.n19 a_41266_55442.n17 7.729
R7928 a_41266_55442.n27 a_41266_55442.n26 6.296
R7929 a_41266_55442.n19 a_41266_55442.n18 6.296
R7930 a_41266_55442.n30 a_41266_55442.n3 4.508
R7931 a_41266_55442.n14 a_41266_55442.n13 4.508
R7932 a_41266_55442.n37 a_41266_55442.n36 4.496
R7933 a_41266_55442.n21 a_41266_55442.n20 4.496
R7934 a_41266_55442.n29 a_41266_55442.n28 4.495
R7935 a_41266_55442.n10 a_41266_55442.n9 4.495
R7936 a_41266_55442.n14 a_41266_55442.n11 4.494
R7937 a_41266_55442.n30 a_41266_55442.n1 4.494
R7938 a_41266_55442.n39 a_41266_55442.t2 1.087
R7939 a_41266_55442.n25 a_41266_55442.n24 0.536
R7940 a_41266_55442.n17 a_41266_55442.n16 0.536
R7941 a_41266_55442.n39 a_41266_55442.n38 0.255
R7942 a_41266_55442.n28 a_41266_55442.n27 0.151
R7943 a_41266_55442.n20 a_41266_55442.n19 0.151
R7944 a_41266_55442.n23 a_41266_55442.n22 0.125
R7945 a_41266_55442.n34 a_41266_55442.n32 0.028
R7946 a_41266_55442.n7 a_41266_55442.n5 0.028
R7947 a_41266_55442.n1 a_41266_55442.n0 0.025
R7948 a_41266_55442.n20 a_41266_55442.n15 0.024
R7949 a_41266_55442.n36 a_41266_55442.n34 0.012
R7950 a_41266_55442.n9 a_41266_55442.n7 0.012
R7951 a_41266_55442.n29 a_41266_55442.n23 0.011
R7952 a_41266_55442.n30 a_41266_55442.n29 0.011
R7953 a_41266_55442.n14 a_41266_55442.n10 0.011
R7954 a_41266_55442.n38 a_41266_55442.n37 0.01
R7955 a_41266_55442.n22 a_41266_55442.n21 0.01
R7956 a_41266_55442.n21 a_41266_55442.n14 0.01
R7957 a_41266_55442.n37 a_41266_55442.n30 0.01
R7958 a_40976_55366.n10 a_40976_55366.t0 10.181
R7959 a_40976_55366.n10 a_40976_55366.t1 10.181
R7960 a_40976_55366.t2 a_40976_55366.n18 9.68
R7961 a_40976_55366.n1 a_40976_55366.n0 9.302
R7962 a_40976_55366.n7 a_40976_55366.n6 9.3
R7963 a_40976_55366.n5 a_40976_55366.n4 9.3
R7964 a_40976_55366.n9 a_40976_55366.n8 9
R7965 a_40976_55366.n13 a_40976_55366.n12 7.729
R7966 a_40976_55366.n13 a_40976_55366.n10 6.296
R7967 a_40976_55366.n16 a_40976_55366.n1 4.508
R7968 a_40976_55366.n15 a_40976_55366.n14 4.501
R7969 a_40976_55366.n15 a_40976_55366.n9 4.501
R7970 a_40976_55366.n16 a_40976_55366.n3 4.494
R7971 a_40976_55366.n18 a_40976_55366.t3 1.259
R7972 a_40976_55366.n12 a_40976_55366.n11 0.536
R7973 a_40976_55366.n18 a_40976_55366.n17 0.415
R7974 a_40976_55366.n14 a_40976_55366.n13 0.151
R7975 a_40976_55366.n7 a_40976_55366.n5 0.028
R7976 a_40976_55366.n3 a_40976_55366.n2 0.025
R7977 a_40976_55366.n17 a_40976_55366.n16 0.021
R7978 a_40976_55366.n9 a_40976_55366.n7 0.012
R7979 a_40976_55366.n16 a_40976_55366.n15 0.006
R7980 a_50176_15846.n10 a_50176_15846.t1 10.181
R7981 a_50176_15846.n10 a_50176_15846.t0 10.181
R7982 a_50176_15846.t3 a_50176_15846.n18 9.68
R7983 a_50176_15846.n1 a_50176_15846.n0 9.302
R7984 a_50176_15846.n7 a_50176_15846.n6 9.3
R7985 a_50176_15846.n5 a_50176_15846.n4 9.3
R7986 a_50176_15846.n9 a_50176_15846.n8 9
R7987 a_50176_15846.n13 a_50176_15846.n12 7.729
R7988 a_50176_15846.n13 a_50176_15846.n10 6.296
R7989 a_50176_15846.n16 a_50176_15846.n1 4.508
R7990 a_50176_15846.n15 a_50176_15846.n14 4.501
R7991 a_50176_15846.n15 a_50176_15846.n9 4.501
R7992 a_50176_15846.n16 a_50176_15846.n3 4.494
R7993 a_50176_15846.n18 a_50176_15846.t2 1.259
R7994 a_50176_15846.n12 a_50176_15846.n11 0.536
R7995 a_50176_15846.n18 a_50176_15846.n17 0.415
R7996 a_50176_15846.n14 a_50176_15846.n13 0.151
R7997 a_50176_15846.n7 a_50176_15846.n5 0.028
R7998 a_50176_15846.n3 a_50176_15846.n2 0.025
R7999 a_50176_15846.n17 a_50176_15846.n16 0.021
R8000 a_50176_15846.n9 a_50176_15846.n7 0.012
R8001 a_50176_15846.n16 a_50176_15846.n15 0.006
R8002 a_50466_15922.n26 a_50466_15922.t1 10.181
R8003 a_50466_15922.n18 a_50466_15922.t0 10.181
R8004 a_50466_15922.t3 a_50466_15922.n39 9.68
R8005 a_50466_15922.n3 a_50466_15922.n2 9.302
R8006 a_50466_15922.n13 a_50466_15922.n12 9.302
R8007 a_50466_15922.n32 a_50466_15922.n31 9.3
R8008 a_50466_15922.n34 a_50466_15922.n33 9.3
R8009 a_50466_15922.n7 a_50466_15922.n6 9.3
R8010 a_50466_15922.n5 a_50466_15922.n4 9.3
R8011 a_50466_15922.n36 a_50466_15922.n35 9
R8012 a_50466_15922.n9 a_50466_15922.n8 9
R8013 a_50466_15922.n27 a_50466_15922.n25 7.729
R8014 a_50466_15922.n19 a_50466_15922.n17 7.729
R8015 a_50466_15922.n27 a_50466_15922.n26 6.296
R8016 a_50466_15922.n19 a_50466_15922.n18 6.296
R8017 a_50466_15922.n30 a_50466_15922.n3 4.508
R8018 a_50466_15922.n14 a_50466_15922.n13 4.508
R8019 a_50466_15922.n37 a_50466_15922.n36 4.496
R8020 a_50466_15922.n21 a_50466_15922.n20 4.496
R8021 a_50466_15922.n29 a_50466_15922.n28 4.495
R8022 a_50466_15922.n10 a_50466_15922.n9 4.495
R8023 a_50466_15922.n14 a_50466_15922.n11 4.494
R8024 a_50466_15922.n30 a_50466_15922.n1 4.494
R8025 a_50466_15922.n39 a_50466_15922.t2 1.087
R8026 a_50466_15922.n25 a_50466_15922.n24 0.536
R8027 a_50466_15922.n17 a_50466_15922.n16 0.536
R8028 a_50466_15922.n39 a_50466_15922.n38 0.255
R8029 a_50466_15922.n28 a_50466_15922.n27 0.151
R8030 a_50466_15922.n20 a_50466_15922.n19 0.151
R8031 a_50466_15922.n23 a_50466_15922.n22 0.125
R8032 a_50466_15922.n34 a_50466_15922.n32 0.028
R8033 a_50466_15922.n7 a_50466_15922.n5 0.028
R8034 a_50466_15922.n1 a_50466_15922.n0 0.025
R8035 a_50466_15922.n20 a_50466_15922.n15 0.024
R8036 a_50466_15922.n36 a_50466_15922.n34 0.012
R8037 a_50466_15922.n9 a_50466_15922.n7 0.012
R8038 a_50466_15922.n29 a_50466_15922.n23 0.011
R8039 a_50466_15922.n30 a_50466_15922.n29 0.011
R8040 a_50466_15922.n14 a_50466_15922.n10 0.011
R8041 a_50466_15922.n38 a_50466_15922.n37 0.01
R8042 a_50466_15922.n22 a_50466_15922.n21 0.01
R8043 a_50466_15922.n21 a_50466_15922.n14 0.01
R8044 a_50466_15922.n37 a_50466_15922.n30 0.01
R8045 a_13376_45486.n10 a_13376_45486.t1 10.181
R8046 a_13376_45486.n10 a_13376_45486.t0 10.181
R8047 a_13376_45486.t2 a_13376_45486.n18 9.68
R8048 a_13376_45486.n1 a_13376_45486.n0 9.302
R8049 a_13376_45486.n7 a_13376_45486.n6 9.3
R8050 a_13376_45486.n5 a_13376_45486.n4 9.3
R8051 a_13376_45486.n9 a_13376_45486.n8 9
R8052 a_13376_45486.n13 a_13376_45486.n12 7.729
R8053 a_13376_45486.n13 a_13376_45486.n10 6.296
R8054 a_13376_45486.n16 a_13376_45486.n1 4.508
R8055 a_13376_45486.n15 a_13376_45486.n14 4.501
R8056 a_13376_45486.n15 a_13376_45486.n9 4.501
R8057 a_13376_45486.n16 a_13376_45486.n3 4.494
R8058 a_13376_45486.n18 a_13376_45486.t3 1.259
R8059 a_13376_45486.n12 a_13376_45486.n11 0.536
R8060 a_13376_45486.n18 a_13376_45486.n17 0.415
R8061 a_13376_45486.n14 a_13376_45486.n13 0.151
R8062 a_13376_45486.n7 a_13376_45486.n5 0.028
R8063 a_13376_45486.n3 a_13376_45486.n2 0.025
R8064 a_13376_45486.n17 a_13376_45486.n16 0.021
R8065 a_13376_45486.n9 a_13376_45486.n7 0.012
R8066 a_13376_45486.n16 a_13376_45486.n15 0.006
R8067 a_22576_5966.n10 a_22576_5966.t1 10.181
R8068 a_22576_5966.n10 a_22576_5966.t0 10.181
R8069 a_22576_5966.t3 a_22576_5966.n18 9.68
R8070 a_22576_5966.n1 a_22576_5966.n0 9.302
R8071 a_22576_5966.n7 a_22576_5966.n6 9.3
R8072 a_22576_5966.n5 a_22576_5966.n4 9.3
R8073 a_22576_5966.n9 a_22576_5966.n8 9
R8074 a_22576_5966.n13 a_22576_5966.n12 7.729
R8075 a_22576_5966.n13 a_22576_5966.n10 6.296
R8076 a_22576_5966.n16 a_22576_5966.n1 4.508
R8077 a_22576_5966.n15 a_22576_5966.n14 4.501
R8078 a_22576_5966.n15 a_22576_5966.n9 4.501
R8079 a_22576_5966.n16 a_22576_5966.n3 4.494
R8080 a_22576_5966.n18 a_22576_5966.t2 1.259
R8081 a_22576_5966.n12 a_22576_5966.n11 0.536
R8082 a_22576_5966.n18 a_22576_5966.n17 0.415
R8083 a_22576_5966.n14 a_22576_5966.n13 0.151
R8084 a_22576_5966.n7 a_22576_5966.n5 0.028
R8085 a_22576_5966.n3 a_22576_5966.n2 0.025
R8086 a_22576_5966.n17 a_22576_5966.n16 0.021
R8087 a_22576_5966.n9 a_22576_5966.n7 0.012
R8088 a_22576_5966.n16 a_22576_5966.n15 0.006
R8089 a_22866_6042.n26 a_22866_6042.t1 10.181
R8090 a_22866_6042.n18 a_22866_6042.t0 10.181
R8091 a_22866_6042.t2 a_22866_6042.n39 9.68
R8092 a_22866_6042.n3 a_22866_6042.n2 9.302
R8093 a_22866_6042.n13 a_22866_6042.n12 9.302
R8094 a_22866_6042.n32 a_22866_6042.n31 9.3
R8095 a_22866_6042.n34 a_22866_6042.n33 9.3
R8096 a_22866_6042.n7 a_22866_6042.n6 9.3
R8097 a_22866_6042.n5 a_22866_6042.n4 9.3
R8098 a_22866_6042.n36 a_22866_6042.n35 9
R8099 a_22866_6042.n9 a_22866_6042.n8 9
R8100 a_22866_6042.n27 a_22866_6042.n25 7.729
R8101 a_22866_6042.n19 a_22866_6042.n17 7.729
R8102 a_22866_6042.n27 a_22866_6042.n26 6.296
R8103 a_22866_6042.n19 a_22866_6042.n18 6.296
R8104 a_22866_6042.n30 a_22866_6042.n3 4.508
R8105 a_22866_6042.n14 a_22866_6042.n13 4.508
R8106 a_22866_6042.n37 a_22866_6042.n36 4.496
R8107 a_22866_6042.n21 a_22866_6042.n20 4.496
R8108 a_22866_6042.n29 a_22866_6042.n28 4.495
R8109 a_22866_6042.n10 a_22866_6042.n9 4.495
R8110 a_22866_6042.n14 a_22866_6042.n11 4.494
R8111 a_22866_6042.n30 a_22866_6042.n1 4.494
R8112 a_22866_6042.n39 a_22866_6042.t3 1.087
R8113 a_22866_6042.n25 a_22866_6042.n24 0.536
R8114 a_22866_6042.n17 a_22866_6042.n16 0.536
R8115 a_22866_6042.n39 a_22866_6042.n38 0.255
R8116 a_22866_6042.n28 a_22866_6042.n27 0.151
R8117 a_22866_6042.n20 a_22866_6042.n19 0.151
R8118 a_22866_6042.n23 a_22866_6042.n22 0.125
R8119 a_22866_6042.n34 a_22866_6042.n32 0.028
R8120 a_22866_6042.n7 a_22866_6042.n5 0.028
R8121 a_22866_6042.n1 a_22866_6042.n0 0.025
R8122 a_22866_6042.n20 a_22866_6042.n15 0.024
R8123 a_22866_6042.n36 a_22866_6042.n34 0.012
R8124 a_22866_6042.n9 a_22866_6042.n7 0.012
R8125 a_22866_6042.n29 a_22866_6042.n23 0.011
R8126 a_22866_6042.n30 a_22866_6042.n29 0.011
R8127 a_22866_6042.n14 a_22866_6042.n10 0.011
R8128 a_22866_6042.n38 a_22866_6042.n37 0.01
R8129 a_22866_6042.n22 a_22866_6042.n21 0.01
R8130 a_22866_6042.n21 a_22866_6042.n14 0.01
R8131 a_22866_6042.n37 a_22866_6042.n30 0.01
R8132 a_13666_65322.n26 a_13666_65322.t0 10.181
R8133 a_13666_65322.n18 a_13666_65322.t3 10.181
R8134 a_13666_65322.t1 a_13666_65322.n39 9.68
R8135 a_13666_65322.n3 a_13666_65322.n2 9.302
R8136 a_13666_65322.n13 a_13666_65322.n12 9.302
R8137 a_13666_65322.n32 a_13666_65322.n31 9.3
R8138 a_13666_65322.n34 a_13666_65322.n33 9.3
R8139 a_13666_65322.n7 a_13666_65322.n6 9.3
R8140 a_13666_65322.n5 a_13666_65322.n4 9.3
R8141 a_13666_65322.n36 a_13666_65322.n35 9
R8142 a_13666_65322.n9 a_13666_65322.n8 9
R8143 a_13666_65322.n27 a_13666_65322.n25 7.729
R8144 a_13666_65322.n19 a_13666_65322.n17 7.729
R8145 a_13666_65322.n27 a_13666_65322.n26 6.296
R8146 a_13666_65322.n19 a_13666_65322.n18 6.296
R8147 a_13666_65322.n30 a_13666_65322.n3 4.508
R8148 a_13666_65322.n14 a_13666_65322.n13 4.508
R8149 a_13666_65322.n37 a_13666_65322.n36 4.496
R8150 a_13666_65322.n21 a_13666_65322.n20 4.496
R8151 a_13666_65322.n29 a_13666_65322.n28 4.495
R8152 a_13666_65322.n10 a_13666_65322.n9 4.495
R8153 a_13666_65322.n14 a_13666_65322.n11 4.494
R8154 a_13666_65322.n30 a_13666_65322.n1 4.494
R8155 a_13666_65322.n39 a_13666_65322.t2 1.087
R8156 a_13666_65322.n25 a_13666_65322.n24 0.536
R8157 a_13666_65322.n17 a_13666_65322.n16 0.536
R8158 a_13666_65322.n39 a_13666_65322.n38 0.255
R8159 a_13666_65322.n28 a_13666_65322.n27 0.151
R8160 a_13666_65322.n20 a_13666_65322.n19 0.151
R8161 a_13666_65322.n23 a_13666_65322.n22 0.125
R8162 a_13666_65322.n34 a_13666_65322.n32 0.028
R8163 a_13666_65322.n7 a_13666_65322.n5 0.028
R8164 a_13666_65322.n1 a_13666_65322.n0 0.025
R8165 a_13666_65322.n20 a_13666_65322.n15 0.024
R8166 a_13666_65322.n36 a_13666_65322.n34 0.012
R8167 a_13666_65322.n9 a_13666_65322.n7 0.012
R8168 a_13666_65322.n29 a_13666_65322.n23 0.011
R8169 a_13666_65322.n30 a_13666_65322.n29 0.011
R8170 a_13666_65322.n14 a_13666_65322.n10 0.011
R8171 a_13666_65322.n38 a_13666_65322.n37 0.01
R8172 a_13666_65322.n22 a_13666_65322.n21 0.01
R8173 a_13666_65322.n21 a_13666_65322.n14 0.01
R8174 a_13666_65322.n37 a_13666_65322.n30 0.01
R8175 a_22866_15922.n26 a_22866_15922.t0 10.181
R8176 a_22866_15922.n18 a_22866_15922.t1 10.181
R8177 a_22866_15922.t2 a_22866_15922.n39 9.68
R8178 a_22866_15922.n3 a_22866_15922.n2 9.302
R8179 a_22866_15922.n13 a_22866_15922.n12 9.302
R8180 a_22866_15922.n32 a_22866_15922.n31 9.3
R8181 a_22866_15922.n34 a_22866_15922.n33 9.3
R8182 a_22866_15922.n7 a_22866_15922.n6 9.3
R8183 a_22866_15922.n5 a_22866_15922.n4 9.3
R8184 a_22866_15922.n36 a_22866_15922.n35 9
R8185 a_22866_15922.n9 a_22866_15922.n8 9
R8186 a_22866_15922.n27 a_22866_15922.n25 7.729
R8187 a_22866_15922.n19 a_22866_15922.n17 7.729
R8188 a_22866_15922.n27 a_22866_15922.n26 6.296
R8189 a_22866_15922.n19 a_22866_15922.n18 6.296
R8190 a_22866_15922.n30 a_22866_15922.n3 4.508
R8191 a_22866_15922.n14 a_22866_15922.n13 4.508
R8192 a_22866_15922.n37 a_22866_15922.n36 4.496
R8193 a_22866_15922.n21 a_22866_15922.n20 4.496
R8194 a_22866_15922.n29 a_22866_15922.n28 4.495
R8195 a_22866_15922.n10 a_22866_15922.n9 4.495
R8196 a_22866_15922.n14 a_22866_15922.n11 4.494
R8197 a_22866_15922.n30 a_22866_15922.n1 4.494
R8198 a_22866_15922.n39 a_22866_15922.t3 1.087
R8199 a_22866_15922.n25 a_22866_15922.n24 0.536
R8200 a_22866_15922.n17 a_22866_15922.n16 0.536
R8201 a_22866_15922.n39 a_22866_15922.n38 0.255
R8202 a_22866_15922.n28 a_22866_15922.n27 0.151
R8203 a_22866_15922.n20 a_22866_15922.n19 0.151
R8204 a_22866_15922.n23 a_22866_15922.n22 0.125
R8205 a_22866_15922.n34 a_22866_15922.n32 0.028
R8206 a_22866_15922.n7 a_22866_15922.n5 0.028
R8207 a_22866_15922.n1 a_22866_15922.n0 0.025
R8208 a_22866_15922.n20 a_22866_15922.n15 0.024
R8209 a_22866_15922.n36 a_22866_15922.n34 0.012
R8210 a_22866_15922.n9 a_22866_15922.n7 0.012
R8211 a_22866_15922.n29 a_22866_15922.n23 0.011
R8212 a_22866_15922.n30 a_22866_15922.n29 0.011
R8213 a_22866_15922.n14 a_22866_15922.n10 0.011
R8214 a_22866_15922.n38 a_22866_15922.n37 0.01
R8215 a_22866_15922.n22 a_22866_15922.n21 0.01
R8216 a_22866_15922.n21 a_22866_15922.n14 0.01
R8217 a_22866_15922.n37 a_22866_15922.n30 0.01
R8218 a_32066_25802.n26 a_32066_25802.t1 10.181
R8219 a_32066_25802.n18 a_32066_25802.t0 10.181
R8220 a_32066_25802.t3 a_32066_25802.n39 9.68
R8221 a_32066_25802.n3 a_32066_25802.n2 9.302
R8222 a_32066_25802.n13 a_32066_25802.n12 9.302
R8223 a_32066_25802.n32 a_32066_25802.n31 9.3
R8224 a_32066_25802.n34 a_32066_25802.n33 9.3
R8225 a_32066_25802.n7 a_32066_25802.n6 9.3
R8226 a_32066_25802.n5 a_32066_25802.n4 9.3
R8227 a_32066_25802.n36 a_32066_25802.n35 9
R8228 a_32066_25802.n9 a_32066_25802.n8 9
R8229 a_32066_25802.n27 a_32066_25802.n25 7.729
R8230 a_32066_25802.n19 a_32066_25802.n17 7.729
R8231 a_32066_25802.n27 a_32066_25802.n26 6.296
R8232 a_32066_25802.n19 a_32066_25802.n18 6.296
R8233 a_32066_25802.n30 a_32066_25802.n3 4.508
R8234 a_32066_25802.n14 a_32066_25802.n13 4.508
R8235 a_32066_25802.n37 a_32066_25802.n36 4.496
R8236 a_32066_25802.n21 a_32066_25802.n20 4.496
R8237 a_32066_25802.n29 a_32066_25802.n28 4.495
R8238 a_32066_25802.n10 a_32066_25802.n9 4.495
R8239 a_32066_25802.n14 a_32066_25802.n11 4.494
R8240 a_32066_25802.n30 a_32066_25802.n1 4.494
R8241 a_32066_25802.n39 a_32066_25802.t2 1.087
R8242 a_32066_25802.n25 a_32066_25802.n24 0.536
R8243 a_32066_25802.n17 a_32066_25802.n16 0.536
R8244 a_32066_25802.n39 a_32066_25802.n38 0.255
R8245 a_32066_25802.n28 a_32066_25802.n27 0.151
R8246 a_32066_25802.n20 a_32066_25802.n19 0.151
R8247 a_32066_25802.n23 a_32066_25802.n22 0.125
R8248 a_32066_25802.n34 a_32066_25802.n32 0.028
R8249 a_32066_25802.n7 a_32066_25802.n5 0.028
R8250 a_32066_25802.n1 a_32066_25802.n0 0.025
R8251 a_32066_25802.n20 a_32066_25802.n15 0.024
R8252 a_32066_25802.n36 a_32066_25802.n34 0.012
R8253 a_32066_25802.n9 a_32066_25802.n7 0.012
R8254 a_32066_25802.n29 a_32066_25802.n23 0.011
R8255 a_32066_25802.n30 a_32066_25802.n29 0.011
R8256 a_32066_25802.n14 a_32066_25802.n10 0.011
R8257 a_32066_25802.n38 a_32066_25802.n37 0.01
R8258 a_32066_25802.n22 a_32066_25802.n21 0.01
R8259 a_32066_25802.n21 a_32066_25802.n14 0.01
R8260 a_32066_25802.n37 a_32066_25802.n30 0.01
R8261 a_50176_35606.n10 a_50176_35606.t1 10.181
R8262 a_50176_35606.n10 a_50176_35606.t0 10.181
R8263 a_50176_35606.t3 a_50176_35606.n18 9.68
R8264 a_50176_35606.n1 a_50176_35606.n0 9.302
R8265 a_50176_35606.n7 a_50176_35606.n6 9.3
R8266 a_50176_35606.n5 a_50176_35606.n4 9.3
R8267 a_50176_35606.n9 a_50176_35606.n8 9
R8268 a_50176_35606.n13 a_50176_35606.n12 7.729
R8269 a_50176_35606.n13 a_50176_35606.n10 6.296
R8270 a_50176_35606.n16 a_50176_35606.n1 4.508
R8271 a_50176_35606.n15 a_50176_35606.n14 4.501
R8272 a_50176_35606.n15 a_50176_35606.n9 4.501
R8273 a_50176_35606.n16 a_50176_35606.n3 4.494
R8274 a_50176_35606.n18 a_50176_35606.t2 1.259
R8275 a_50176_35606.n12 a_50176_35606.n11 0.536
R8276 a_50176_35606.n18 a_50176_35606.n17 0.415
R8277 a_50176_35606.n14 a_50176_35606.n13 0.151
R8278 a_50176_35606.n7 a_50176_35606.n5 0.028
R8279 a_50176_35606.n3 a_50176_35606.n2 0.025
R8280 a_50176_35606.n17 a_50176_35606.n16 0.021
R8281 a_50176_35606.n9 a_50176_35606.n7 0.012
R8282 a_50176_35606.n16 a_50176_35606.n15 0.006
R8283 a_59666_15922.n26 a_59666_15922.t1 10.181
R8284 a_59666_15922.n18 a_59666_15922.t2 10.181
R8285 a_59666_15922.t0 a_59666_15922.n39 9.68
R8286 a_59666_15922.n3 a_59666_15922.n2 9.302
R8287 a_59666_15922.n13 a_59666_15922.n12 9.302
R8288 a_59666_15922.n32 a_59666_15922.n31 9.3
R8289 a_59666_15922.n34 a_59666_15922.n33 9.3
R8290 a_59666_15922.n7 a_59666_15922.n6 9.3
R8291 a_59666_15922.n5 a_59666_15922.n4 9.3
R8292 a_59666_15922.n36 a_59666_15922.n35 9
R8293 a_59666_15922.n9 a_59666_15922.n8 9
R8294 a_59666_15922.n27 a_59666_15922.n25 7.729
R8295 a_59666_15922.n19 a_59666_15922.n17 7.729
R8296 a_59666_15922.n27 a_59666_15922.n26 6.296
R8297 a_59666_15922.n19 a_59666_15922.n18 6.296
R8298 a_59666_15922.n30 a_59666_15922.n3 4.508
R8299 a_59666_15922.n14 a_59666_15922.n13 4.508
R8300 a_59666_15922.n37 a_59666_15922.n36 4.496
R8301 a_59666_15922.n21 a_59666_15922.n20 4.496
R8302 a_59666_15922.n29 a_59666_15922.n28 4.495
R8303 a_59666_15922.n10 a_59666_15922.n9 4.495
R8304 a_59666_15922.n14 a_59666_15922.n11 4.494
R8305 a_59666_15922.n30 a_59666_15922.n1 4.494
R8306 a_59666_15922.n39 a_59666_15922.t3 1.087
R8307 a_59666_15922.n25 a_59666_15922.n24 0.536
R8308 a_59666_15922.n17 a_59666_15922.n16 0.536
R8309 a_59666_15922.n39 a_59666_15922.n38 0.255
R8310 a_59666_15922.n28 a_59666_15922.n27 0.151
R8311 a_59666_15922.n20 a_59666_15922.n19 0.151
R8312 a_59666_15922.n23 a_59666_15922.n22 0.125
R8313 a_59666_15922.n34 a_59666_15922.n32 0.028
R8314 a_59666_15922.n7 a_59666_15922.n5 0.028
R8315 a_59666_15922.n1 a_59666_15922.n0 0.025
R8316 a_59666_15922.n20 a_59666_15922.n15 0.024
R8317 a_59666_15922.n36 a_59666_15922.n34 0.012
R8318 a_59666_15922.n9 a_59666_15922.n7 0.012
R8319 a_59666_15922.n29 a_59666_15922.n23 0.011
R8320 a_59666_15922.n30 a_59666_15922.n29 0.011
R8321 a_59666_15922.n14 a_59666_15922.n10 0.011
R8322 a_59666_15922.n38 a_59666_15922.n37 0.01
R8323 a_59666_15922.n22 a_59666_15922.n21 0.01
R8324 a_59666_15922.n21 a_59666_15922.n14 0.01
R8325 a_59666_15922.n37 a_59666_15922.n30 0.01
R8326 a_59376_15846.n10 a_59376_15846.t0 10.181
R8327 a_59376_15846.n10 a_59376_15846.t1 10.181
R8328 a_59376_15846.t2 a_59376_15846.n18 9.68
R8329 a_59376_15846.n1 a_59376_15846.n0 9.302
R8330 a_59376_15846.n7 a_59376_15846.n6 9.3
R8331 a_59376_15846.n5 a_59376_15846.n4 9.3
R8332 a_59376_15846.n9 a_59376_15846.n8 9
R8333 a_59376_15846.n13 a_59376_15846.n12 7.729
R8334 a_59376_15846.n13 a_59376_15846.n10 6.296
R8335 a_59376_15846.n16 a_59376_15846.n1 4.508
R8336 a_59376_15846.n15 a_59376_15846.n14 4.501
R8337 a_59376_15846.n15 a_59376_15846.n9 4.501
R8338 a_59376_15846.n16 a_59376_15846.n3 4.494
R8339 a_59376_15846.n18 a_59376_15846.t3 1.259
R8340 a_59376_15846.n12 a_59376_15846.n11 0.536
R8341 a_59376_15846.n18 a_59376_15846.n17 0.415
R8342 a_59376_15846.n14 a_59376_15846.n13 0.151
R8343 a_59376_15846.n7 a_59376_15846.n5 0.028
R8344 a_59376_15846.n3 a_59376_15846.n2 0.025
R8345 a_59376_15846.n17 a_59376_15846.n16 0.021
R8346 a_59376_15846.n9 a_59376_15846.n7 0.012
R8347 a_59376_15846.n16 a_59376_15846.n15 0.006
R8348 a_59376_55366.n10 a_59376_55366.t1 10.181
R8349 a_59376_55366.n10 a_59376_55366.t0 10.181
R8350 a_59376_55366.t3 a_59376_55366.n18 9.68
R8351 a_59376_55366.n1 a_59376_55366.n0 9.302
R8352 a_59376_55366.n7 a_59376_55366.n6 9.3
R8353 a_59376_55366.n5 a_59376_55366.n4 9.3
R8354 a_59376_55366.n9 a_59376_55366.n8 9
R8355 a_59376_55366.n13 a_59376_55366.n12 7.729
R8356 a_59376_55366.n13 a_59376_55366.n10 6.296
R8357 a_59376_55366.n16 a_59376_55366.n1 4.508
R8358 a_59376_55366.n15 a_59376_55366.n14 4.501
R8359 a_59376_55366.n15 a_59376_55366.n9 4.501
R8360 a_59376_55366.n16 a_59376_55366.n3 4.494
R8361 a_59376_55366.n18 a_59376_55366.t2 1.259
R8362 a_59376_55366.n12 a_59376_55366.n11 0.536
R8363 a_59376_55366.n18 a_59376_55366.n17 0.415
R8364 a_59376_55366.n14 a_59376_55366.n13 0.151
R8365 a_59376_55366.n7 a_59376_55366.n5 0.028
R8366 a_59376_55366.n3 a_59376_55366.n2 0.025
R8367 a_59376_55366.n17 a_59376_55366.n16 0.021
R8368 a_59376_55366.n9 a_59376_55366.n7 0.012
R8369 a_59376_55366.n16 a_59376_55366.n15 0.006
R8370 a_13376_25726.n10 a_13376_25726.t1 10.181
R8371 a_13376_25726.n10 a_13376_25726.t0 10.181
R8372 a_13376_25726.t3 a_13376_25726.n18 9.68
R8373 a_13376_25726.n1 a_13376_25726.n0 9.302
R8374 a_13376_25726.n7 a_13376_25726.n6 9.3
R8375 a_13376_25726.n5 a_13376_25726.n4 9.3
R8376 a_13376_25726.n9 a_13376_25726.n8 9
R8377 a_13376_25726.n13 a_13376_25726.n12 7.729
R8378 a_13376_25726.n13 a_13376_25726.n10 6.296
R8379 a_13376_25726.n16 a_13376_25726.n1 4.508
R8380 a_13376_25726.n15 a_13376_25726.n14 4.501
R8381 a_13376_25726.n15 a_13376_25726.n9 4.501
R8382 a_13376_25726.n16 a_13376_25726.n3 4.494
R8383 a_13376_25726.n18 a_13376_25726.t2 1.259
R8384 a_13376_25726.n12 a_13376_25726.n11 0.536
R8385 a_13376_25726.n18 a_13376_25726.n17 0.415
R8386 a_13376_25726.n14 a_13376_25726.n13 0.151
R8387 a_13376_25726.n7 a_13376_25726.n5 0.028
R8388 a_13376_25726.n3 a_13376_25726.n2 0.025
R8389 a_13376_25726.n17 a_13376_25726.n16 0.021
R8390 a_13376_25726.n9 a_13376_25726.n7 0.012
R8391 a_13376_25726.n16 a_13376_25726.n15 0.006
R8392 a_13666_25802.n26 a_13666_25802.t1 10.181
R8393 a_13666_25802.n18 a_13666_25802.t0 10.181
R8394 a_13666_25802.t3 a_13666_25802.n39 9.68
R8395 a_13666_25802.n3 a_13666_25802.n2 9.302
R8396 a_13666_25802.n13 a_13666_25802.n12 9.302
R8397 a_13666_25802.n32 a_13666_25802.n31 9.3
R8398 a_13666_25802.n34 a_13666_25802.n33 9.3
R8399 a_13666_25802.n7 a_13666_25802.n6 9.3
R8400 a_13666_25802.n5 a_13666_25802.n4 9.3
R8401 a_13666_25802.n36 a_13666_25802.n35 9
R8402 a_13666_25802.n9 a_13666_25802.n8 9
R8403 a_13666_25802.n27 a_13666_25802.n25 7.729
R8404 a_13666_25802.n19 a_13666_25802.n17 7.729
R8405 a_13666_25802.n27 a_13666_25802.n26 6.296
R8406 a_13666_25802.n19 a_13666_25802.n18 6.296
R8407 a_13666_25802.n30 a_13666_25802.n3 4.508
R8408 a_13666_25802.n14 a_13666_25802.n13 4.508
R8409 a_13666_25802.n37 a_13666_25802.n36 4.496
R8410 a_13666_25802.n21 a_13666_25802.n20 4.496
R8411 a_13666_25802.n29 a_13666_25802.n28 4.495
R8412 a_13666_25802.n10 a_13666_25802.n9 4.495
R8413 a_13666_25802.n14 a_13666_25802.n11 4.494
R8414 a_13666_25802.n30 a_13666_25802.n1 4.494
R8415 a_13666_25802.n39 a_13666_25802.t2 1.087
R8416 a_13666_25802.n25 a_13666_25802.n24 0.536
R8417 a_13666_25802.n17 a_13666_25802.n16 0.536
R8418 a_13666_25802.n39 a_13666_25802.n38 0.255
R8419 a_13666_25802.n28 a_13666_25802.n27 0.151
R8420 a_13666_25802.n20 a_13666_25802.n19 0.151
R8421 a_13666_25802.n23 a_13666_25802.n22 0.125
R8422 a_13666_25802.n34 a_13666_25802.n32 0.028
R8423 a_13666_25802.n7 a_13666_25802.n5 0.028
R8424 a_13666_25802.n1 a_13666_25802.n0 0.025
R8425 a_13666_25802.n20 a_13666_25802.n15 0.024
R8426 a_13666_25802.n36 a_13666_25802.n34 0.012
R8427 a_13666_25802.n9 a_13666_25802.n7 0.012
R8428 a_13666_25802.n29 a_13666_25802.n23 0.011
R8429 a_13666_25802.n30 a_13666_25802.n29 0.011
R8430 a_13666_25802.n14 a_13666_25802.n10 0.011
R8431 a_13666_25802.n38 a_13666_25802.n37 0.01
R8432 a_13666_25802.n22 a_13666_25802.n21 0.01
R8433 a_13666_25802.n21 a_13666_25802.n14 0.01
R8434 a_13666_25802.n37 a_13666_25802.n30 0.01
R8435 a_4176_25726.n10 a_4176_25726.t0 10.181
R8436 a_4176_25726.n10 a_4176_25726.t1 10.181
R8437 a_4176_25726.t3 a_4176_25726.n18 9.68
R8438 a_4176_25726.n1 a_4176_25726.n0 9.302
R8439 a_4176_25726.n7 a_4176_25726.n6 9.3
R8440 a_4176_25726.n5 a_4176_25726.n4 9.3
R8441 a_4176_25726.n9 a_4176_25726.n8 9
R8442 a_4176_25726.n13 a_4176_25726.n12 7.729
R8443 a_4176_25726.n13 a_4176_25726.n10 6.296
R8444 a_4176_25726.n16 a_4176_25726.n1 4.508
R8445 a_4176_25726.n15 a_4176_25726.n14 4.501
R8446 a_4176_25726.n15 a_4176_25726.n9 4.501
R8447 a_4176_25726.n16 a_4176_25726.n3 4.494
R8448 a_4176_25726.n18 a_4176_25726.t2 1.259
R8449 a_4176_25726.n12 a_4176_25726.n11 0.536
R8450 a_4176_25726.n18 a_4176_25726.n17 0.415
R8451 a_4176_25726.n14 a_4176_25726.n13 0.151
R8452 a_4176_25726.n7 a_4176_25726.n5 0.028
R8453 a_4176_25726.n3 a_4176_25726.n2 0.025
R8454 a_4176_25726.n17 a_4176_25726.n16 0.021
R8455 a_4176_25726.n9 a_4176_25726.n7 0.012
R8456 a_4176_25726.n16 a_4176_25726.n15 0.006
R8457 a_31776_35606.n10 a_31776_35606.t1 10.181
R8458 a_31776_35606.n10 a_31776_35606.t0 10.181
R8459 a_31776_35606.t3 a_31776_35606.n18 9.68
R8460 a_31776_35606.n1 a_31776_35606.n0 9.302
R8461 a_31776_35606.n7 a_31776_35606.n6 9.3
R8462 a_31776_35606.n5 a_31776_35606.n4 9.3
R8463 a_31776_35606.n9 a_31776_35606.n8 9
R8464 a_31776_35606.n13 a_31776_35606.n12 7.729
R8465 a_31776_35606.n13 a_31776_35606.n10 6.296
R8466 a_31776_35606.n16 a_31776_35606.n1 4.508
R8467 a_31776_35606.n15 a_31776_35606.n14 4.501
R8468 a_31776_35606.n15 a_31776_35606.n9 4.501
R8469 a_31776_35606.n16 a_31776_35606.n3 4.494
R8470 a_31776_35606.n18 a_31776_35606.t2 1.259
R8471 a_31776_35606.n12 a_31776_35606.n11 0.536
R8472 a_31776_35606.n18 a_31776_35606.n17 0.415
R8473 a_31776_35606.n14 a_31776_35606.n13 0.151
R8474 a_31776_35606.n7 a_31776_35606.n5 0.028
R8475 a_31776_35606.n3 a_31776_35606.n2 0.025
R8476 a_31776_35606.n17 a_31776_35606.n16 0.021
R8477 a_31776_35606.n9 a_31776_35606.n7 0.012
R8478 a_31776_35606.n16 a_31776_35606.n15 0.006
R8479 a_68866_6042.n26 a_68866_6042.t1 10.181
R8480 a_68866_6042.n18 a_68866_6042.t2 10.181
R8481 a_68866_6042.t0 a_68866_6042.n39 9.68
R8482 a_68866_6042.n3 a_68866_6042.n2 9.302
R8483 a_68866_6042.n13 a_68866_6042.n12 9.302
R8484 a_68866_6042.n32 a_68866_6042.n31 9.3
R8485 a_68866_6042.n34 a_68866_6042.n33 9.3
R8486 a_68866_6042.n7 a_68866_6042.n6 9.3
R8487 a_68866_6042.n5 a_68866_6042.n4 9.3
R8488 a_68866_6042.n36 a_68866_6042.n35 9
R8489 a_68866_6042.n9 a_68866_6042.n8 9
R8490 a_68866_6042.n27 a_68866_6042.n25 7.729
R8491 a_68866_6042.n19 a_68866_6042.n17 7.729
R8492 a_68866_6042.n27 a_68866_6042.n26 6.296
R8493 a_68866_6042.n19 a_68866_6042.n18 6.296
R8494 a_68866_6042.n30 a_68866_6042.n3 4.508
R8495 a_68866_6042.n14 a_68866_6042.n13 4.508
R8496 a_68866_6042.n37 a_68866_6042.n36 4.496
R8497 a_68866_6042.n21 a_68866_6042.n20 4.496
R8498 a_68866_6042.n29 a_68866_6042.n28 4.495
R8499 a_68866_6042.n10 a_68866_6042.n9 4.495
R8500 a_68866_6042.n14 a_68866_6042.n11 4.494
R8501 a_68866_6042.n30 a_68866_6042.n1 4.494
R8502 a_68866_6042.n39 a_68866_6042.t3 1.087
R8503 a_68866_6042.n25 a_68866_6042.n24 0.536
R8504 a_68866_6042.n17 a_68866_6042.n16 0.536
R8505 a_68866_6042.n39 a_68866_6042.n38 0.255
R8506 a_68866_6042.n28 a_68866_6042.n27 0.151
R8507 a_68866_6042.n20 a_68866_6042.n19 0.151
R8508 a_68866_6042.n23 a_68866_6042.n22 0.125
R8509 a_68866_6042.n34 a_68866_6042.n32 0.028
R8510 a_68866_6042.n7 a_68866_6042.n5 0.028
R8511 a_68866_6042.n1 a_68866_6042.n0 0.025
R8512 a_68866_6042.n20 a_68866_6042.n15 0.024
R8513 a_68866_6042.n36 a_68866_6042.n34 0.012
R8514 a_68866_6042.n9 a_68866_6042.n7 0.012
R8515 a_68866_6042.n29 a_68866_6042.n23 0.011
R8516 a_68866_6042.n30 a_68866_6042.n29 0.011
R8517 a_68866_6042.n14 a_68866_6042.n10 0.011
R8518 a_68866_6042.n38 a_68866_6042.n37 0.01
R8519 a_68866_6042.n22 a_68866_6042.n21 0.01
R8520 a_68866_6042.n21 a_68866_6042.n14 0.01
R8521 a_68866_6042.n37 a_68866_6042.n30 0.01
R8522 a_50466_55442.n26 a_50466_55442.t0 10.181
R8523 a_50466_55442.n18 a_50466_55442.t1 10.181
R8524 a_50466_55442.t3 a_50466_55442.n39 9.68
R8525 a_50466_55442.n3 a_50466_55442.n2 9.302
R8526 a_50466_55442.n13 a_50466_55442.n12 9.302
R8527 a_50466_55442.n32 a_50466_55442.n31 9.3
R8528 a_50466_55442.n34 a_50466_55442.n33 9.3
R8529 a_50466_55442.n7 a_50466_55442.n6 9.3
R8530 a_50466_55442.n5 a_50466_55442.n4 9.3
R8531 a_50466_55442.n36 a_50466_55442.n35 9
R8532 a_50466_55442.n9 a_50466_55442.n8 9
R8533 a_50466_55442.n27 a_50466_55442.n25 7.729
R8534 a_50466_55442.n19 a_50466_55442.n17 7.729
R8535 a_50466_55442.n27 a_50466_55442.n26 6.296
R8536 a_50466_55442.n19 a_50466_55442.n18 6.296
R8537 a_50466_55442.n30 a_50466_55442.n3 4.508
R8538 a_50466_55442.n14 a_50466_55442.n13 4.508
R8539 a_50466_55442.n37 a_50466_55442.n36 4.496
R8540 a_50466_55442.n21 a_50466_55442.n20 4.496
R8541 a_50466_55442.n29 a_50466_55442.n28 4.495
R8542 a_50466_55442.n10 a_50466_55442.n9 4.495
R8543 a_50466_55442.n14 a_50466_55442.n11 4.494
R8544 a_50466_55442.n30 a_50466_55442.n1 4.494
R8545 a_50466_55442.n39 a_50466_55442.t2 1.087
R8546 a_50466_55442.n25 a_50466_55442.n24 0.536
R8547 a_50466_55442.n17 a_50466_55442.n16 0.536
R8548 a_50466_55442.n39 a_50466_55442.n38 0.255
R8549 a_50466_55442.n28 a_50466_55442.n27 0.151
R8550 a_50466_55442.n20 a_50466_55442.n19 0.151
R8551 a_50466_55442.n23 a_50466_55442.n22 0.125
R8552 a_50466_55442.n34 a_50466_55442.n32 0.028
R8553 a_50466_55442.n7 a_50466_55442.n5 0.028
R8554 a_50466_55442.n1 a_50466_55442.n0 0.025
R8555 a_50466_55442.n20 a_50466_55442.n15 0.024
R8556 a_50466_55442.n36 a_50466_55442.n34 0.012
R8557 a_50466_55442.n9 a_50466_55442.n7 0.012
R8558 a_50466_55442.n29 a_50466_55442.n23 0.011
R8559 a_50466_55442.n30 a_50466_55442.n29 0.011
R8560 a_50466_55442.n14 a_50466_55442.n10 0.011
R8561 a_50466_55442.n38 a_50466_55442.n37 0.01
R8562 a_50466_55442.n22 a_50466_55442.n21 0.01
R8563 a_50466_55442.n21 a_50466_55442.n14 0.01
R8564 a_50466_55442.n37 a_50466_55442.n30 0.01
R8565 a_41266_25802.n26 a_41266_25802.t1 10.181
R8566 a_41266_25802.n18 a_41266_25802.t0 10.181
R8567 a_41266_25802.t2 a_41266_25802.n39 9.68
R8568 a_41266_25802.n3 a_41266_25802.n2 9.302
R8569 a_41266_25802.n13 a_41266_25802.n12 9.302
R8570 a_41266_25802.n32 a_41266_25802.n31 9.3
R8571 a_41266_25802.n34 a_41266_25802.n33 9.3
R8572 a_41266_25802.n7 a_41266_25802.n6 9.3
R8573 a_41266_25802.n5 a_41266_25802.n4 9.3
R8574 a_41266_25802.n36 a_41266_25802.n35 9
R8575 a_41266_25802.n9 a_41266_25802.n8 9
R8576 a_41266_25802.n27 a_41266_25802.n25 7.729
R8577 a_41266_25802.n19 a_41266_25802.n17 7.729
R8578 a_41266_25802.n27 a_41266_25802.n26 6.296
R8579 a_41266_25802.n19 a_41266_25802.n18 6.296
R8580 a_41266_25802.n30 a_41266_25802.n3 4.508
R8581 a_41266_25802.n14 a_41266_25802.n13 4.508
R8582 a_41266_25802.n37 a_41266_25802.n36 4.496
R8583 a_41266_25802.n21 a_41266_25802.n20 4.496
R8584 a_41266_25802.n29 a_41266_25802.n28 4.495
R8585 a_41266_25802.n10 a_41266_25802.n9 4.495
R8586 a_41266_25802.n14 a_41266_25802.n11 4.494
R8587 a_41266_25802.n30 a_41266_25802.n1 4.494
R8588 a_41266_25802.n39 a_41266_25802.t3 1.087
R8589 a_41266_25802.n25 a_41266_25802.n24 0.536
R8590 a_41266_25802.n17 a_41266_25802.n16 0.536
R8591 a_41266_25802.n39 a_41266_25802.n38 0.255
R8592 a_41266_25802.n28 a_41266_25802.n27 0.151
R8593 a_41266_25802.n20 a_41266_25802.n19 0.151
R8594 a_41266_25802.n23 a_41266_25802.n22 0.125
R8595 a_41266_25802.n34 a_41266_25802.n32 0.028
R8596 a_41266_25802.n7 a_41266_25802.n5 0.028
R8597 a_41266_25802.n1 a_41266_25802.n0 0.025
R8598 a_41266_25802.n20 a_41266_25802.n15 0.024
R8599 a_41266_25802.n36 a_41266_25802.n34 0.012
R8600 a_41266_25802.n9 a_41266_25802.n7 0.012
R8601 a_41266_25802.n29 a_41266_25802.n23 0.011
R8602 a_41266_25802.n30 a_41266_25802.n29 0.011
R8603 a_41266_25802.n14 a_41266_25802.n10 0.011
R8604 a_41266_25802.n38 a_41266_25802.n37 0.01
R8605 a_41266_25802.n22 a_41266_25802.n21 0.01
R8606 a_41266_25802.n21 a_41266_25802.n14 0.01
R8607 a_41266_25802.n37 a_41266_25802.n30 0.01
R8608 a_32066_15922.n26 a_32066_15922.t1 10.181
R8609 a_32066_15922.n18 a_32066_15922.t2 10.181
R8610 a_32066_15922.t0 a_32066_15922.n39 9.68
R8611 a_32066_15922.n3 a_32066_15922.n2 9.302
R8612 a_32066_15922.n13 a_32066_15922.n12 9.302
R8613 a_32066_15922.n32 a_32066_15922.n31 9.3
R8614 a_32066_15922.n34 a_32066_15922.n33 9.3
R8615 a_32066_15922.n7 a_32066_15922.n6 9.3
R8616 a_32066_15922.n5 a_32066_15922.n4 9.3
R8617 a_32066_15922.n36 a_32066_15922.n35 9
R8618 a_32066_15922.n9 a_32066_15922.n8 9
R8619 a_32066_15922.n27 a_32066_15922.n25 7.729
R8620 a_32066_15922.n19 a_32066_15922.n17 7.729
R8621 a_32066_15922.n27 a_32066_15922.n26 6.296
R8622 a_32066_15922.n19 a_32066_15922.n18 6.296
R8623 a_32066_15922.n30 a_32066_15922.n3 4.508
R8624 a_32066_15922.n14 a_32066_15922.n13 4.508
R8625 a_32066_15922.n37 a_32066_15922.n36 4.496
R8626 a_32066_15922.n21 a_32066_15922.n20 4.496
R8627 a_32066_15922.n29 a_32066_15922.n28 4.495
R8628 a_32066_15922.n10 a_32066_15922.n9 4.495
R8629 a_32066_15922.n14 a_32066_15922.n11 4.494
R8630 a_32066_15922.n30 a_32066_15922.n1 4.494
R8631 a_32066_15922.n39 a_32066_15922.t3 1.087
R8632 a_32066_15922.n25 a_32066_15922.n24 0.536
R8633 a_32066_15922.n17 a_32066_15922.n16 0.536
R8634 a_32066_15922.n39 a_32066_15922.n38 0.255
R8635 a_32066_15922.n28 a_32066_15922.n27 0.151
R8636 a_32066_15922.n20 a_32066_15922.n19 0.151
R8637 a_32066_15922.n23 a_32066_15922.n22 0.125
R8638 a_32066_15922.n34 a_32066_15922.n32 0.028
R8639 a_32066_15922.n7 a_32066_15922.n5 0.028
R8640 a_32066_15922.n1 a_32066_15922.n0 0.025
R8641 a_32066_15922.n20 a_32066_15922.n15 0.024
R8642 a_32066_15922.n36 a_32066_15922.n34 0.012
R8643 a_32066_15922.n9 a_32066_15922.n7 0.012
R8644 a_32066_15922.n29 a_32066_15922.n23 0.011
R8645 a_32066_15922.n30 a_32066_15922.n29 0.011
R8646 a_32066_15922.n14 a_32066_15922.n10 0.011
R8647 a_32066_15922.n38 a_32066_15922.n37 0.01
R8648 a_32066_15922.n22 a_32066_15922.n21 0.01
R8649 a_32066_15922.n21 a_32066_15922.n14 0.01
R8650 a_32066_15922.n37 a_32066_15922.n30 0.01
R8651 bit3.n56 bit3.t14 552.693
R8652 bit3.n2 bit3.t7 300.446
R8653 bit3.n0 bit3.t16 300.446
R8654 bit3.n9 bit3.t8 300.446
R8655 bit3.n7 bit3.t15 300.446
R8656 bit3.n16 bit3.t13 300.446
R8657 bit3.n14 bit3.t5 300.446
R8658 bit3.n23 bit3.t12 300.446
R8659 bit3.n21 bit3.t3 300.446
R8660 bit3.n30 bit3.t10 300.446
R8661 bit3.n28 bit3.t1 300.446
R8662 bit3.n37 bit3.t9 300.446
R8663 bit3.n35 bit3.t4 300.446
R8664 bit3.n44 bit3.t11 300.446
R8665 bit3.n42 bit3.t2 300.446
R8666 bit3.n53 bit3.t17 300.446
R8667 bit3.n51 bit3.t6 300.446
R8668 bit3.n56 bit3.t0 279.56
R8669 bit3.n57 bit3.n56 120.317
R8670 bit3.n52 bit3.n51 27.537
R8671 bit3.n5 bit3.n2 27.536
R8672 bit3.n12 bit3.n9 27.536
R8673 bit3.n19 bit3.n16 27.536
R8674 bit3.n26 bit3.n23 27.536
R8675 bit3.n33 bit3.n30 27.536
R8676 bit3.n40 bit3.n37 27.536
R8677 bit3.n47 bit3.n44 27.536
R8678 bit3.n1 bit3.n0 24.127
R8679 bit3.n8 bit3.n7 24.127
R8680 bit3.n15 bit3.n14 24.127
R8681 bit3.n22 bit3.n21 24.127
R8682 bit3.n29 bit3.n28 24.127
R8683 bit3.n36 bit3.n35 24.127
R8684 bit3.n43 bit3.n42 24.127
R8685 bit3.n54 bit3.n53 24.127
R8686 bit3.n4 bit3.n3 8.764
R8687 bit3.n11 bit3.n10 8.764
R8688 bit3.n18 bit3.n17 8.764
R8689 bit3.n25 bit3.n24 8.764
R8690 bit3.n32 bit3.n31 8.764
R8691 bit3.n39 bit3.n38 8.764
R8692 bit3.n46 bit3.n45 8.764
R8693 bit3.n50 bit3.n49 8.764
R8694 bit3.n6 bit3.n1 4.662
R8695 bit3.n13 bit3.n8 4.662
R8696 bit3.n20 bit3.n15 4.662
R8697 bit3.n27 bit3.n22 4.662
R8698 bit3.n34 bit3.n29 4.662
R8699 bit3.n41 bit3.n36 4.662
R8700 bit3.n48 bit3.n43 4.662
R8701 bit3.n55 bit3.n54 4.661
R8702 bit3.n5 bit3.n4 3.401
R8703 bit3.n12 bit3.n11 3.401
R8704 bit3.n19 bit3.n18 3.401
R8705 bit3.n26 bit3.n25 3.401
R8706 bit3.n33 bit3.n32 3.401
R8707 bit3.n40 bit3.n39 3.401
R8708 bit3.n47 bit3.n46 3.401
R8709 bit3.n52 bit3.n50 3.401
R8710 bit3 bit3.n64 0.851
R8711 bit3.n55 bit3.n52 0.626
R8712 bit3.n6 bit3.n5 0.626
R8713 bit3.n13 bit3.n12 0.626
R8714 bit3.n20 bit3.n19 0.626
R8715 bit3.n27 bit3.n26 0.626
R8716 bit3.n34 bit3.n33 0.626
R8717 bit3.n41 bit3.n40 0.626
R8718 bit3.n48 bit3.n47 0.626
R8719 bit3.n64 bit3.n63 0.575
R8720 bit3.n63 bit3.n62 0.575
R8721 bit3.n62 bit3.n61 0.575
R8722 bit3.n61 bit3.n60 0.575
R8723 bit3.n60 bit3.n59 0.575
R8724 bit3.n59 bit3.n58 0.575
R8725 bit3.n58 bit3.n57 0.575
R8726 bit3.n64 bit3.n6 0.298
R8727 bit3.n63 bit3.n13 0.298
R8728 bit3.n62 bit3.n20 0.298
R8729 bit3.n61 bit3.n27 0.298
R8730 bit3.n60 bit3.n34 0.298
R8731 bit3.n59 bit3.n41 0.298
R8732 bit3.n58 bit3.n48 0.298
R8733 bit3.n57 bit3.n55 0.298
R8734 a_32066_65322.n26 a_32066_65322.t0 10.181
R8735 a_32066_65322.n18 a_32066_65322.t1 10.181
R8736 a_32066_65322.t3 a_32066_65322.n39 9.68
R8737 a_32066_65322.n3 a_32066_65322.n2 9.302
R8738 a_32066_65322.n13 a_32066_65322.n12 9.302
R8739 a_32066_65322.n32 a_32066_65322.n31 9.3
R8740 a_32066_65322.n34 a_32066_65322.n33 9.3
R8741 a_32066_65322.n7 a_32066_65322.n6 9.3
R8742 a_32066_65322.n5 a_32066_65322.n4 9.3
R8743 a_32066_65322.n36 a_32066_65322.n35 9
R8744 a_32066_65322.n9 a_32066_65322.n8 9
R8745 a_32066_65322.n27 a_32066_65322.n25 7.729
R8746 a_32066_65322.n19 a_32066_65322.n17 7.729
R8747 a_32066_65322.n27 a_32066_65322.n26 6.296
R8748 a_32066_65322.n19 a_32066_65322.n18 6.296
R8749 a_32066_65322.n30 a_32066_65322.n3 4.508
R8750 a_32066_65322.n14 a_32066_65322.n13 4.508
R8751 a_32066_65322.n37 a_32066_65322.n36 4.496
R8752 a_32066_65322.n21 a_32066_65322.n20 4.496
R8753 a_32066_65322.n29 a_32066_65322.n28 4.495
R8754 a_32066_65322.n10 a_32066_65322.n9 4.495
R8755 a_32066_65322.n14 a_32066_65322.n11 4.494
R8756 a_32066_65322.n30 a_32066_65322.n1 4.494
R8757 a_32066_65322.n39 a_32066_65322.t2 1.087
R8758 a_32066_65322.n25 a_32066_65322.n24 0.536
R8759 a_32066_65322.n17 a_32066_65322.n16 0.536
R8760 a_32066_65322.n39 a_32066_65322.n38 0.255
R8761 a_32066_65322.n28 a_32066_65322.n27 0.151
R8762 a_32066_65322.n20 a_32066_65322.n19 0.151
R8763 a_32066_65322.n23 a_32066_65322.n22 0.125
R8764 a_32066_65322.n34 a_32066_65322.n32 0.028
R8765 a_32066_65322.n7 a_32066_65322.n5 0.028
R8766 a_32066_65322.n1 a_32066_65322.n0 0.025
R8767 a_32066_65322.n20 a_32066_65322.n15 0.024
R8768 a_32066_65322.n36 a_32066_65322.n34 0.012
R8769 a_32066_65322.n9 a_32066_65322.n7 0.012
R8770 a_32066_65322.n29 a_32066_65322.n23 0.011
R8771 a_32066_65322.n30 a_32066_65322.n29 0.011
R8772 a_32066_65322.n14 a_32066_65322.n10 0.011
R8773 a_32066_65322.n38 a_32066_65322.n37 0.01
R8774 a_32066_65322.n22 a_32066_65322.n21 0.01
R8775 a_32066_65322.n21 a_32066_65322.n14 0.01
R8776 a_32066_65322.n37 a_32066_65322.n30 0.01
R8777 a_31776_65246.n10 a_31776_65246.t0 10.181
R8778 a_31776_65246.n10 a_31776_65246.t1 10.181
R8779 a_31776_65246.t3 a_31776_65246.n18 9.68
R8780 a_31776_65246.n1 a_31776_65246.n0 9.302
R8781 a_31776_65246.n7 a_31776_65246.n6 9.3
R8782 a_31776_65246.n5 a_31776_65246.n4 9.3
R8783 a_31776_65246.n9 a_31776_65246.n8 9
R8784 a_31776_65246.n13 a_31776_65246.n12 7.729
R8785 a_31776_65246.n13 a_31776_65246.n10 6.296
R8786 a_31776_65246.n16 a_31776_65246.n1 4.508
R8787 a_31776_65246.n15 a_31776_65246.n14 4.501
R8788 a_31776_65246.n15 a_31776_65246.n9 4.501
R8789 a_31776_65246.n16 a_31776_65246.n3 4.494
R8790 a_31776_65246.n18 a_31776_65246.t2 1.259
R8791 a_31776_65246.n12 a_31776_65246.n11 0.536
R8792 a_31776_65246.n18 a_31776_65246.n17 0.415
R8793 a_31776_65246.n14 a_31776_65246.n13 0.151
R8794 a_31776_65246.n7 a_31776_65246.n5 0.028
R8795 a_31776_65246.n3 a_31776_65246.n2 0.025
R8796 a_31776_65246.n17 a_31776_65246.n16 0.021
R8797 a_31776_65246.n9 a_31776_65246.n7 0.012
R8798 a_31776_65246.n16 a_31776_65246.n15 0.006
R8799 a_59376_35606.n10 a_59376_35606.t2 10.181
R8800 a_59376_35606.n10 a_59376_35606.t1 10.181
R8801 a_59376_35606.t0 a_59376_35606.n18 9.68
R8802 a_59376_35606.n1 a_59376_35606.n0 9.302
R8803 a_59376_35606.n7 a_59376_35606.n6 9.3
R8804 a_59376_35606.n5 a_59376_35606.n4 9.3
R8805 a_59376_35606.n9 a_59376_35606.n8 9
R8806 a_59376_35606.n13 a_59376_35606.n12 7.729
R8807 a_59376_35606.n13 a_59376_35606.n10 6.296
R8808 a_59376_35606.n16 a_59376_35606.n1 4.508
R8809 a_59376_35606.n15 a_59376_35606.n14 4.501
R8810 a_59376_35606.n15 a_59376_35606.n9 4.501
R8811 a_59376_35606.n16 a_59376_35606.n3 4.494
R8812 a_59376_35606.n18 a_59376_35606.t3 1.259
R8813 a_59376_35606.n12 a_59376_35606.n11 0.536
R8814 a_59376_35606.n18 a_59376_35606.n17 0.415
R8815 a_59376_35606.n14 a_59376_35606.n13 0.151
R8816 a_59376_35606.n7 a_59376_35606.n5 0.028
R8817 a_59376_35606.n3 a_59376_35606.n2 0.025
R8818 a_59376_35606.n17 a_59376_35606.n16 0.021
R8819 a_59376_35606.n9 a_59376_35606.n7 0.012
R8820 a_59376_35606.n16 a_59376_35606.n15 0.006
R8821 a_59666_35682.n26 a_59666_35682.t2 10.181
R8822 a_59666_35682.n18 a_59666_35682.t1 10.181
R8823 a_59666_35682.t0 a_59666_35682.n39 9.68
R8824 a_59666_35682.n3 a_59666_35682.n2 9.302
R8825 a_59666_35682.n13 a_59666_35682.n12 9.302
R8826 a_59666_35682.n32 a_59666_35682.n31 9.3
R8827 a_59666_35682.n34 a_59666_35682.n33 9.3
R8828 a_59666_35682.n7 a_59666_35682.n6 9.3
R8829 a_59666_35682.n5 a_59666_35682.n4 9.3
R8830 a_59666_35682.n36 a_59666_35682.n35 9
R8831 a_59666_35682.n9 a_59666_35682.n8 9
R8832 a_59666_35682.n27 a_59666_35682.n25 7.729
R8833 a_59666_35682.n19 a_59666_35682.n17 7.729
R8834 a_59666_35682.n27 a_59666_35682.n26 6.296
R8835 a_59666_35682.n19 a_59666_35682.n18 6.296
R8836 a_59666_35682.n30 a_59666_35682.n3 4.508
R8837 a_59666_35682.n14 a_59666_35682.n13 4.508
R8838 a_59666_35682.n37 a_59666_35682.n36 4.496
R8839 a_59666_35682.n21 a_59666_35682.n20 4.496
R8840 a_59666_35682.n29 a_59666_35682.n28 4.495
R8841 a_59666_35682.n10 a_59666_35682.n9 4.495
R8842 a_59666_35682.n14 a_59666_35682.n11 4.494
R8843 a_59666_35682.n30 a_59666_35682.n1 4.494
R8844 a_59666_35682.n39 a_59666_35682.t3 1.087
R8845 a_59666_35682.n25 a_59666_35682.n24 0.536
R8846 a_59666_35682.n17 a_59666_35682.n16 0.536
R8847 a_59666_35682.n39 a_59666_35682.n38 0.255
R8848 a_59666_35682.n28 a_59666_35682.n27 0.151
R8849 a_59666_35682.n20 a_59666_35682.n19 0.151
R8850 a_59666_35682.n23 a_59666_35682.n22 0.125
R8851 a_59666_35682.n34 a_59666_35682.n32 0.028
R8852 a_59666_35682.n7 a_59666_35682.n5 0.028
R8853 a_59666_35682.n1 a_59666_35682.n0 0.025
R8854 a_59666_35682.n20 a_59666_35682.n15 0.024
R8855 a_59666_35682.n36 a_59666_35682.n34 0.012
R8856 a_59666_35682.n9 a_59666_35682.n7 0.012
R8857 a_59666_35682.n29 a_59666_35682.n23 0.011
R8858 a_59666_35682.n30 a_59666_35682.n29 0.011
R8859 a_59666_35682.n14 a_59666_35682.n10 0.011
R8860 a_59666_35682.n38 a_59666_35682.n37 0.01
R8861 a_59666_35682.n22 a_59666_35682.n21 0.01
R8862 a_59666_35682.n21 a_59666_35682.n14 0.01
R8863 a_59666_35682.n37 a_59666_35682.n30 0.01
R8864 a_68866_15922.n26 a_68866_15922.t1 10.181
R8865 a_68866_15922.n18 a_68866_15922.t0 10.181
R8866 a_68866_15922.t3 a_68866_15922.n39 9.68
R8867 a_68866_15922.n3 a_68866_15922.n2 9.302
R8868 a_68866_15922.n13 a_68866_15922.n12 9.302
R8869 a_68866_15922.n32 a_68866_15922.n31 9.3
R8870 a_68866_15922.n34 a_68866_15922.n33 9.3
R8871 a_68866_15922.n7 a_68866_15922.n6 9.3
R8872 a_68866_15922.n5 a_68866_15922.n4 9.3
R8873 a_68866_15922.n36 a_68866_15922.n35 9
R8874 a_68866_15922.n9 a_68866_15922.n8 9
R8875 a_68866_15922.n27 a_68866_15922.n25 7.729
R8876 a_68866_15922.n19 a_68866_15922.n17 7.729
R8877 a_68866_15922.n27 a_68866_15922.n26 6.296
R8878 a_68866_15922.n19 a_68866_15922.n18 6.296
R8879 a_68866_15922.n30 a_68866_15922.n3 4.508
R8880 a_68866_15922.n14 a_68866_15922.n13 4.508
R8881 a_68866_15922.n37 a_68866_15922.n36 4.496
R8882 a_68866_15922.n21 a_68866_15922.n20 4.496
R8883 a_68866_15922.n29 a_68866_15922.n28 4.495
R8884 a_68866_15922.n10 a_68866_15922.n9 4.495
R8885 a_68866_15922.n14 a_68866_15922.n11 4.494
R8886 a_68866_15922.n30 a_68866_15922.n1 4.494
R8887 a_68866_15922.n39 a_68866_15922.t2 1.087
R8888 a_68866_15922.n25 a_68866_15922.n24 0.536
R8889 a_68866_15922.n17 a_68866_15922.n16 0.536
R8890 a_68866_15922.n39 a_68866_15922.n38 0.255
R8891 a_68866_15922.n28 a_68866_15922.n27 0.151
R8892 a_68866_15922.n20 a_68866_15922.n19 0.151
R8893 a_68866_15922.n23 a_68866_15922.n22 0.125
R8894 a_68866_15922.n34 a_68866_15922.n32 0.028
R8895 a_68866_15922.n7 a_68866_15922.n5 0.028
R8896 a_68866_15922.n1 a_68866_15922.n0 0.025
R8897 a_68866_15922.n20 a_68866_15922.n15 0.024
R8898 a_68866_15922.n36 a_68866_15922.n34 0.012
R8899 a_68866_15922.n9 a_68866_15922.n7 0.012
R8900 a_68866_15922.n29 a_68866_15922.n23 0.011
R8901 a_68866_15922.n30 a_68866_15922.n29 0.011
R8902 a_68866_15922.n14 a_68866_15922.n10 0.011
R8903 a_68866_15922.n38 a_68866_15922.n37 0.01
R8904 a_68866_15922.n22 a_68866_15922.n21 0.01
R8905 a_68866_15922.n21 a_68866_15922.n14 0.01
R8906 a_68866_15922.n37 a_68866_15922.n30 0.01
R8907 a_68576_15846.n10 a_68576_15846.t0 10.181
R8908 a_68576_15846.n10 a_68576_15846.t1 10.181
R8909 a_68576_15846.t2 a_68576_15846.n18 9.68
R8910 a_68576_15846.n1 a_68576_15846.n0 9.302
R8911 a_68576_15846.n7 a_68576_15846.n6 9.3
R8912 a_68576_15846.n5 a_68576_15846.n4 9.3
R8913 a_68576_15846.n9 a_68576_15846.n8 9
R8914 a_68576_15846.n13 a_68576_15846.n12 7.729
R8915 a_68576_15846.n13 a_68576_15846.n10 6.296
R8916 a_68576_15846.n16 a_68576_15846.n1 4.508
R8917 a_68576_15846.n15 a_68576_15846.n14 4.501
R8918 a_68576_15846.n15 a_68576_15846.n9 4.501
R8919 a_68576_15846.n16 a_68576_15846.n3 4.494
R8920 a_68576_15846.n18 a_68576_15846.t3 1.259
R8921 a_68576_15846.n12 a_68576_15846.n11 0.536
R8922 a_68576_15846.n18 a_68576_15846.n17 0.415
R8923 a_68576_15846.n14 a_68576_15846.n13 0.151
R8924 a_68576_15846.n7 a_68576_15846.n5 0.028
R8925 a_68576_15846.n3 a_68576_15846.n2 0.025
R8926 a_68576_15846.n17 a_68576_15846.n16 0.021
R8927 a_68576_15846.n9 a_68576_15846.n7 0.012
R8928 a_68576_15846.n16 a_68576_15846.n15 0.006
R8929 a_n436_74606.t4 a_n436_74606.n7 139.026
R8930 a_n436_74606.n7 a_n436_74606.t3 85.389
R8931 a_n436_74606.n7 a_n436_74606.n6 54.371
R8932 a_n436_74606.n0 a_n436_74606.t8 9.633
R8933 a_n436_74606.n6 a_n436_74606.t6 9.587
R8934 a_n436_74606.n5 a_n436_74606.t9 9.587
R8935 a_n436_74606.n4 a_n436_74606.t5 9.587
R8936 a_n436_74606.n3 a_n436_74606.t0 9.587
R8937 a_n436_74606.n2 a_n436_74606.t2 9.587
R8938 a_n436_74606.n1 a_n436_74606.t7 9.587
R8939 a_n436_74606.n0 a_n436_74606.t1 9.587
R8940 a_n436_74606.n1 a_n436_74606.n0 0.528
R8941 a_n436_74606.n3 a_n436_74606.n2 0.528
R8942 a_n436_74606.n5 a_n436_74606.n4 0.528
R8943 a_n436_74606.n2 a_n436_74606.n1 0.046
R8944 a_n436_74606.n4 a_n436_74606.n3 0.046
R8945 a_n436_74606.n6 a_n436_74606.n5 0.046
R8946 a_4466_45562.n26 a_4466_45562.t0 10.181
R8947 a_4466_45562.n18 a_4466_45562.t1 10.181
R8948 a_4466_45562.t3 a_4466_45562.n39 9.68
R8949 a_4466_45562.n3 a_4466_45562.n2 9.302
R8950 a_4466_45562.n13 a_4466_45562.n12 9.302
R8951 a_4466_45562.n32 a_4466_45562.n31 9.3
R8952 a_4466_45562.n34 a_4466_45562.n33 9.3
R8953 a_4466_45562.n7 a_4466_45562.n6 9.3
R8954 a_4466_45562.n5 a_4466_45562.n4 9.3
R8955 a_4466_45562.n36 a_4466_45562.n35 9
R8956 a_4466_45562.n9 a_4466_45562.n8 9
R8957 a_4466_45562.n27 a_4466_45562.n25 7.729
R8958 a_4466_45562.n19 a_4466_45562.n17 7.729
R8959 a_4466_45562.n27 a_4466_45562.n26 6.296
R8960 a_4466_45562.n19 a_4466_45562.n18 6.296
R8961 a_4466_45562.n30 a_4466_45562.n3 4.508
R8962 a_4466_45562.n14 a_4466_45562.n13 4.508
R8963 a_4466_45562.n37 a_4466_45562.n36 4.496
R8964 a_4466_45562.n21 a_4466_45562.n20 4.496
R8965 a_4466_45562.n29 a_4466_45562.n28 4.495
R8966 a_4466_45562.n10 a_4466_45562.n9 4.495
R8967 a_4466_45562.n14 a_4466_45562.n11 4.494
R8968 a_4466_45562.n30 a_4466_45562.n1 4.494
R8969 a_4466_45562.n39 a_4466_45562.t2 1.087
R8970 a_4466_45562.n25 a_4466_45562.n24 0.536
R8971 a_4466_45562.n17 a_4466_45562.n16 0.536
R8972 a_4466_45562.n39 a_4466_45562.n38 0.255
R8973 a_4466_45562.n28 a_4466_45562.n27 0.151
R8974 a_4466_45562.n20 a_4466_45562.n19 0.151
R8975 a_4466_45562.n23 a_4466_45562.n22 0.125
R8976 a_4466_45562.n34 a_4466_45562.n32 0.028
R8977 a_4466_45562.n7 a_4466_45562.n5 0.028
R8978 a_4466_45562.n1 a_4466_45562.n0 0.025
R8979 a_4466_45562.n20 a_4466_45562.n15 0.024
R8980 a_4466_45562.n36 a_4466_45562.n34 0.012
R8981 a_4466_45562.n9 a_4466_45562.n7 0.012
R8982 a_4466_45562.n29 a_4466_45562.n23 0.011
R8983 a_4466_45562.n30 a_4466_45562.n29 0.011
R8984 a_4466_45562.n14 a_4466_45562.n10 0.011
R8985 a_4466_45562.n38 a_4466_45562.n37 0.01
R8986 a_4466_45562.n22 a_4466_45562.n21 0.01
R8987 a_4466_45562.n21 a_4466_45562.n14 0.01
R8988 a_4466_45562.n37 a_4466_45562.n30 0.01
R8989 a_4176_45486.n10 a_4176_45486.t0 10.181
R8990 a_4176_45486.n10 a_4176_45486.t1 10.181
R8991 a_4176_45486.t2 a_4176_45486.n18 9.68
R8992 a_4176_45486.n1 a_4176_45486.n0 9.302
R8993 a_4176_45486.n7 a_4176_45486.n6 9.3
R8994 a_4176_45486.n5 a_4176_45486.n4 9.3
R8995 a_4176_45486.n9 a_4176_45486.n8 9
R8996 a_4176_45486.n13 a_4176_45486.n12 7.729
R8997 a_4176_45486.n13 a_4176_45486.n10 6.296
R8998 a_4176_45486.n16 a_4176_45486.n1 4.508
R8999 a_4176_45486.n15 a_4176_45486.n14 4.501
R9000 a_4176_45486.n15 a_4176_45486.n9 4.501
R9001 a_4176_45486.n16 a_4176_45486.n3 4.494
R9002 a_4176_45486.n18 a_4176_45486.t3 1.259
R9003 a_4176_45486.n12 a_4176_45486.n11 0.536
R9004 a_4176_45486.n18 a_4176_45486.n17 0.415
R9005 a_4176_45486.n14 a_4176_45486.n13 0.151
R9006 a_4176_45486.n7 a_4176_45486.n5 0.028
R9007 a_4176_45486.n3 a_4176_45486.n2 0.025
R9008 a_4176_45486.n17 a_4176_45486.n16 0.021
R9009 a_4176_45486.n9 a_4176_45486.n7 0.012
R9010 a_4176_45486.n16 a_4176_45486.n15 0.006
R9011 a_68576_55366.n10 a_68576_55366.t1 10.181
R9012 a_68576_55366.n10 a_68576_55366.t0 10.181
R9013 a_68576_55366.t3 a_68576_55366.n18 9.68
R9014 a_68576_55366.n1 a_68576_55366.n0 9.302
R9015 a_68576_55366.n7 a_68576_55366.n6 9.3
R9016 a_68576_55366.n5 a_68576_55366.n4 9.3
R9017 a_68576_55366.n9 a_68576_55366.n8 9
R9018 a_68576_55366.n13 a_68576_55366.n12 7.729
R9019 a_68576_55366.n13 a_68576_55366.n10 6.296
R9020 a_68576_55366.n16 a_68576_55366.n1 4.508
R9021 a_68576_55366.n15 a_68576_55366.n14 4.501
R9022 a_68576_55366.n15 a_68576_55366.n9 4.501
R9023 a_68576_55366.n16 a_68576_55366.n3 4.494
R9024 a_68576_55366.n18 a_68576_55366.t2 1.259
R9025 a_68576_55366.n12 a_68576_55366.n11 0.536
R9026 a_68576_55366.n18 a_68576_55366.n17 0.415
R9027 a_68576_55366.n14 a_68576_55366.n13 0.151
R9028 a_68576_55366.n7 a_68576_55366.n5 0.028
R9029 a_68576_55366.n3 a_68576_55366.n2 0.025
R9030 a_68576_55366.n17 a_68576_55366.n16 0.021
R9031 a_68576_55366.n9 a_68576_55366.n7 0.012
R9032 a_68576_55366.n16 a_68576_55366.n15 0.006
R9033 a_68576_5966.n10 a_68576_5966.t1 10.181
R9034 a_68576_5966.n10 a_68576_5966.t2 10.181
R9035 a_68576_5966.t0 a_68576_5966.n18 9.68
R9036 a_68576_5966.n1 a_68576_5966.n0 9.302
R9037 a_68576_5966.n7 a_68576_5966.n6 9.3
R9038 a_68576_5966.n5 a_68576_5966.n4 9.3
R9039 a_68576_5966.n9 a_68576_5966.n8 9
R9040 a_68576_5966.n13 a_68576_5966.n12 7.729
R9041 a_68576_5966.n13 a_68576_5966.n10 6.296
R9042 a_68576_5966.n16 a_68576_5966.n1 4.508
R9043 a_68576_5966.n15 a_68576_5966.n14 4.501
R9044 a_68576_5966.n15 a_68576_5966.n9 4.501
R9045 a_68576_5966.n16 a_68576_5966.n3 4.494
R9046 a_68576_5966.n18 a_68576_5966.t3 1.259
R9047 a_68576_5966.n12 a_68576_5966.n11 0.536
R9048 a_68576_5966.n18 a_68576_5966.n17 0.415
R9049 a_68576_5966.n14 a_68576_5966.n13 0.151
R9050 a_68576_5966.n7 a_68576_5966.n5 0.028
R9051 a_68576_5966.n3 a_68576_5966.n2 0.025
R9052 a_68576_5966.n17 a_68576_5966.n16 0.021
R9053 a_68576_5966.n9 a_68576_5966.n7 0.012
R9054 a_68576_5966.n16 a_68576_5966.n15 0.006
R9055 a_4176_85006.n10 a_4176_85006.t2 10.181
R9056 a_4176_85006.n10 a_4176_85006.t3 10.181
R9057 a_4176_85006.t1 a_4176_85006.n18 9.68
R9058 a_4176_85006.n1 a_4176_85006.n0 9.302
R9059 a_4176_85006.n7 a_4176_85006.n6 9.3
R9060 a_4176_85006.n5 a_4176_85006.n4 9.3
R9061 a_4176_85006.n9 a_4176_85006.n8 9
R9062 a_4176_85006.n13 a_4176_85006.n12 7.729
R9063 a_4176_85006.n13 a_4176_85006.n10 6.296
R9064 a_4176_85006.n16 a_4176_85006.n1 4.508
R9065 a_4176_85006.n15 a_4176_85006.n14 4.501
R9066 a_4176_85006.n15 a_4176_85006.n9 4.501
R9067 a_4176_85006.n16 a_4176_85006.n3 4.494
R9068 a_4176_85006.n18 a_4176_85006.t0 1.259
R9069 a_4176_85006.n12 a_4176_85006.n11 0.536
R9070 a_4176_85006.n18 a_4176_85006.n17 0.415
R9071 a_4176_85006.n14 a_4176_85006.n13 0.151
R9072 a_4176_85006.n7 a_4176_85006.n5 0.028
R9073 a_4176_85006.n3 a_4176_85006.n2 0.025
R9074 a_4176_85006.n17 a_4176_85006.n16 0.021
R9075 a_4176_85006.n9 a_4176_85006.n7 0.012
R9076 a_4176_85006.n16 a_4176_85006.n15 0.006
R9077 a_59666_6042.n26 a_59666_6042.t2 10.181
R9078 a_59666_6042.n18 a_59666_6042.t1 10.181
R9079 a_59666_6042.t0 a_59666_6042.n39 9.68
R9080 a_59666_6042.n3 a_59666_6042.n2 9.302
R9081 a_59666_6042.n13 a_59666_6042.n12 9.302
R9082 a_59666_6042.n32 a_59666_6042.n31 9.3
R9083 a_59666_6042.n34 a_59666_6042.n33 9.3
R9084 a_59666_6042.n7 a_59666_6042.n6 9.3
R9085 a_59666_6042.n5 a_59666_6042.n4 9.3
R9086 a_59666_6042.n36 a_59666_6042.n35 9
R9087 a_59666_6042.n9 a_59666_6042.n8 9
R9088 a_59666_6042.n27 a_59666_6042.n25 7.729
R9089 a_59666_6042.n19 a_59666_6042.n17 7.729
R9090 a_59666_6042.n27 a_59666_6042.n26 6.296
R9091 a_59666_6042.n19 a_59666_6042.n18 6.296
R9092 a_59666_6042.n30 a_59666_6042.n3 4.508
R9093 a_59666_6042.n14 a_59666_6042.n13 4.508
R9094 a_59666_6042.n37 a_59666_6042.n36 4.496
R9095 a_59666_6042.n21 a_59666_6042.n20 4.496
R9096 a_59666_6042.n29 a_59666_6042.n28 4.495
R9097 a_59666_6042.n10 a_59666_6042.n9 4.495
R9098 a_59666_6042.n14 a_59666_6042.n11 4.494
R9099 a_59666_6042.n30 a_59666_6042.n1 4.494
R9100 a_59666_6042.n39 a_59666_6042.t3 1.087
R9101 a_59666_6042.n25 a_59666_6042.n24 0.536
R9102 a_59666_6042.n17 a_59666_6042.n16 0.536
R9103 a_59666_6042.n39 a_59666_6042.n38 0.255
R9104 a_59666_6042.n28 a_59666_6042.n27 0.151
R9105 a_59666_6042.n20 a_59666_6042.n19 0.151
R9106 a_59666_6042.n23 a_59666_6042.n22 0.125
R9107 a_59666_6042.n34 a_59666_6042.n32 0.028
R9108 a_59666_6042.n7 a_59666_6042.n5 0.028
R9109 a_59666_6042.n1 a_59666_6042.n0 0.025
R9110 a_59666_6042.n20 a_59666_6042.n15 0.024
R9111 a_59666_6042.n36 a_59666_6042.n34 0.012
R9112 a_59666_6042.n9 a_59666_6042.n7 0.012
R9113 a_59666_6042.n29 a_59666_6042.n23 0.011
R9114 a_59666_6042.n30 a_59666_6042.n29 0.011
R9115 a_59666_6042.n14 a_59666_6042.n10 0.011
R9116 a_59666_6042.n38 a_59666_6042.n37 0.01
R9117 a_59666_6042.n22 a_59666_6042.n21 0.01
R9118 a_59666_6042.n21 a_59666_6042.n14 0.01
R9119 a_59666_6042.n37 a_59666_6042.n30 0.01
R9120 a_13376_5966.n10 a_13376_5966.t1 10.181
R9121 a_13376_5966.n10 a_13376_5966.t0 10.181
R9122 a_13376_5966.t3 a_13376_5966.n18 9.68
R9123 a_13376_5966.n1 a_13376_5966.n0 9.302
R9124 a_13376_5966.n7 a_13376_5966.n6 9.3
R9125 a_13376_5966.n5 a_13376_5966.n4 9.3
R9126 a_13376_5966.n9 a_13376_5966.n8 9
R9127 a_13376_5966.n13 a_13376_5966.n12 7.729
R9128 a_13376_5966.n13 a_13376_5966.n10 6.296
R9129 a_13376_5966.n16 a_13376_5966.n1 4.508
R9130 a_13376_5966.n15 a_13376_5966.n14 4.501
R9131 a_13376_5966.n15 a_13376_5966.n9 4.501
R9132 a_13376_5966.n16 a_13376_5966.n3 4.494
R9133 a_13376_5966.n18 a_13376_5966.t2 1.259
R9134 a_13376_5966.n12 a_13376_5966.n11 0.536
R9135 a_13376_5966.n18 a_13376_5966.n17 0.415
R9136 a_13376_5966.n14 a_13376_5966.n13 0.151
R9137 a_13376_5966.n7 a_13376_5966.n5 0.028
R9138 a_13376_5966.n3 a_13376_5966.n2 0.025
R9139 a_13376_5966.n17 a_13376_5966.n16 0.021
R9140 a_13376_5966.n9 a_13376_5966.n7 0.012
R9141 a_13376_5966.n16 a_13376_5966.n15 0.006
R9142 a_13666_6042.n26 a_13666_6042.t1 10.181
R9143 a_13666_6042.n18 a_13666_6042.t0 10.181
R9144 a_13666_6042.t3 a_13666_6042.n39 9.68
R9145 a_13666_6042.n3 a_13666_6042.n2 9.302
R9146 a_13666_6042.n13 a_13666_6042.n12 9.302
R9147 a_13666_6042.n32 a_13666_6042.n31 9.3
R9148 a_13666_6042.n34 a_13666_6042.n33 9.3
R9149 a_13666_6042.n7 a_13666_6042.n6 9.3
R9150 a_13666_6042.n5 a_13666_6042.n4 9.3
R9151 a_13666_6042.n36 a_13666_6042.n35 9
R9152 a_13666_6042.n9 a_13666_6042.n8 9
R9153 a_13666_6042.n27 a_13666_6042.n25 7.729
R9154 a_13666_6042.n19 a_13666_6042.n17 7.729
R9155 a_13666_6042.n27 a_13666_6042.n26 6.296
R9156 a_13666_6042.n19 a_13666_6042.n18 6.296
R9157 a_13666_6042.n30 a_13666_6042.n3 4.508
R9158 a_13666_6042.n14 a_13666_6042.n13 4.508
R9159 a_13666_6042.n37 a_13666_6042.n36 4.496
R9160 a_13666_6042.n21 a_13666_6042.n20 4.496
R9161 a_13666_6042.n29 a_13666_6042.n28 4.495
R9162 a_13666_6042.n10 a_13666_6042.n9 4.495
R9163 a_13666_6042.n14 a_13666_6042.n11 4.494
R9164 a_13666_6042.n30 a_13666_6042.n1 4.494
R9165 a_13666_6042.n39 a_13666_6042.t2 1.087
R9166 a_13666_6042.n25 a_13666_6042.n24 0.536
R9167 a_13666_6042.n17 a_13666_6042.n16 0.536
R9168 a_13666_6042.n39 a_13666_6042.n38 0.255
R9169 a_13666_6042.n28 a_13666_6042.n27 0.151
R9170 a_13666_6042.n20 a_13666_6042.n19 0.151
R9171 a_13666_6042.n23 a_13666_6042.n22 0.125
R9172 a_13666_6042.n34 a_13666_6042.n32 0.028
R9173 a_13666_6042.n7 a_13666_6042.n5 0.028
R9174 a_13666_6042.n1 a_13666_6042.n0 0.025
R9175 a_13666_6042.n20 a_13666_6042.n15 0.024
R9176 a_13666_6042.n36 a_13666_6042.n34 0.012
R9177 a_13666_6042.n9 a_13666_6042.n7 0.012
R9178 a_13666_6042.n29 a_13666_6042.n23 0.011
R9179 a_13666_6042.n30 a_13666_6042.n29 0.011
R9180 a_13666_6042.n14 a_13666_6042.n10 0.011
R9181 a_13666_6042.n38 a_13666_6042.n37 0.01
R9182 a_13666_6042.n22 a_13666_6042.n21 0.01
R9183 a_13666_6042.n21 a_13666_6042.n14 0.01
R9184 a_13666_6042.n37 a_13666_6042.n30 0.01
R9185 a_40976_35606.n10 a_40976_35606.t2 10.181
R9186 a_40976_35606.n10 a_40976_35606.t1 10.181
R9187 a_40976_35606.t0 a_40976_35606.n18 9.68
R9188 a_40976_35606.n1 a_40976_35606.n0 9.302
R9189 a_40976_35606.n7 a_40976_35606.n6 9.3
R9190 a_40976_35606.n5 a_40976_35606.n4 9.3
R9191 a_40976_35606.n9 a_40976_35606.n8 9
R9192 a_40976_35606.n13 a_40976_35606.n12 7.729
R9193 a_40976_35606.n13 a_40976_35606.n10 6.296
R9194 a_40976_35606.n16 a_40976_35606.n1 4.508
R9195 a_40976_35606.n15 a_40976_35606.n14 4.501
R9196 a_40976_35606.n15 a_40976_35606.n9 4.501
R9197 a_40976_35606.n16 a_40976_35606.n3 4.494
R9198 a_40976_35606.n18 a_40976_35606.t3 1.259
R9199 a_40976_35606.n12 a_40976_35606.n11 0.536
R9200 a_40976_35606.n18 a_40976_35606.n17 0.415
R9201 a_40976_35606.n14 a_40976_35606.n13 0.151
R9202 a_40976_35606.n7 a_40976_35606.n5 0.028
R9203 a_40976_35606.n3 a_40976_35606.n2 0.025
R9204 a_40976_35606.n17 a_40976_35606.n16 0.021
R9205 a_40976_35606.n9 a_40976_35606.n7 0.012
R9206 a_40976_35606.n16 a_40976_35606.n15 0.006
R9207 a_68576_45486.n10 a_68576_45486.t1 10.181
R9208 a_68576_45486.n10 a_68576_45486.t0 10.181
R9209 a_68576_45486.t3 a_68576_45486.n18 9.68
R9210 a_68576_45486.n1 a_68576_45486.n0 9.302
R9211 a_68576_45486.n7 a_68576_45486.n6 9.3
R9212 a_68576_45486.n5 a_68576_45486.n4 9.3
R9213 a_68576_45486.n9 a_68576_45486.n8 9
R9214 a_68576_45486.n13 a_68576_45486.n12 7.729
R9215 a_68576_45486.n13 a_68576_45486.n10 6.296
R9216 a_68576_45486.n16 a_68576_45486.n1 4.508
R9217 a_68576_45486.n15 a_68576_45486.n14 4.501
R9218 a_68576_45486.n15 a_68576_45486.n9 4.501
R9219 a_68576_45486.n16 a_68576_45486.n3 4.494
R9220 a_68576_45486.n18 a_68576_45486.t2 1.259
R9221 a_68576_45486.n12 a_68576_45486.n11 0.536
R9222 a_68576_45486.n18 a_68576_45486.n17 0.415
R9223 a_68576_45486.n14 a_68576_45486.n13 0.151
R9224 a_68576_45486.n7 a_68576_45486.n5 0.028
R9225 a_68576_45486.n3 a_68576_45486.n2 0.025
R9226 a_68576_45486.n17 a_68576_45486.n16 0.021
R9227 a_68576_45486.n9 a_68576_45486.n7 0.012
R9228 a_68576_45486.n16 a_68576_45486.n15 0.006
R9229 a_50176_25726.n10 a_50176_25726.t1 10.181
R9230 a_50176_25726.n10 a_50176_25726.t0 10.181
R9231 a_50176_25726.t3 a_50176_25726.n18 9.68
R9232 a_50176_25726.n1 a_50176_25726.n0 9.302
R9233 a_50176_25726.n7 a_50176_25726.n6 9.3
R9234 a_50176_25726.n5 a_50176_25726.n4 9.3
R9235 a_50176_25726.n9 a_50176_25726.n8 9
R9236 a_50176_25726.n13 a_50176_25726.n12 7.729
R9237 a_50176_25726.n13 a_50176_25726.n10 6.296
R9238 a_50176_25726.n16 a_50176_25726.n1 4.508
R9239 a_50176_25726.n15 a_50176_25726.n14 4.501
R9240 a_50176_25726.n15 a_50176_25726.n9 4.501
R9241 a_50176_25726.n16 a_50176_25726.n3 4.494
R9242 a_50176_25726.n18 a_50176_25726.t2 1.259
R9243 a_50176_25726.n12 a_50176_25726.n11 0.536
R9244 a_50176_25726.n18 a_50176_25726.n17 0.415
R9245 a_50176_25726.n14 a_50176_25726.n13 0.151
R9246 a_50176_25726.n7 a_50176_25726.n5 0.028
R9247 a_50176_25726.n3 a_50176_25726.n2 0.025
R9248 a_50176_25726.n17 a_50176_25726.n16 0.021
R9249 a_50176_25726.n9 a_50176_25726.n7 0.012
R9250 a_50176_25726.n16 a_50176_25726.n15 0.006
R9251 a_50466_25802.n26 a_50466_25802.t1 10.181
R9252 a_50466_25802.n18 a_50466_25802.t0 10.181
R9253 a_50466_25802.t3 a_50466_25802.n39 9.68
R9254 a_50466_25802.n3 a_50466_25802.n2 9.302
R9255 a_50466_25802.n13 a_50466_25802.n12 9.302
R9256 a_50466_25802.n32 a_50466_25802.n31 9.3
R9257 a_50466_25802.n34 a_50466_25802.n33 9.3
R9258 a_50466_25802.n7 a_50466_25802.n6 9.3
R9259 a_50466_25802.n5 a_50466_25802.n4 9.3
R9260 a_50466_25802.n36 a_50466_25802.n35 9
R9261 a_50466_25802.n9 a_50466_25802.n8 9
R9262 a_50466_25802.n27 a_50466_25802.n25 7.729
R9263 a_50466_25802.n19 a_50466_25802.n17 7.729
R9264 a_50466_25802.n27 a_50466_25802.n26 6.296
R9265 a_50466_25802.n19 a_50466_25802.n18 6.296
R9266 a_50466_25802.n30 a_50466_25802.n3 4.508
R9267 a_50466_25802.n14 a_50466_25802.n13 4.508
R9268 a_50466_25802.n37 a_50466_25802.n36 4.496
R9269 a_50466_25802.n21 a_50466_25802.n20 4.496
R9270 a_50466_25802.n29 a_50466_25802.n28 4.495
R9271 a_50466_25802.n10 a_50466_25802.n9 4.495
R9272 a_50466_25802.n14 a_50466_25802.n11 4.494
R9273 a_50466_25802.n30 a_50466_25802.n1 4.494
R9274 a_50466_25802.n39 a_50466_25802.t2 1.087
R9275 a_50466_25802.n25 a_50466_25802.n24 0.536
R9276 a_50466_25802.n17 a_50466_25802.n16 0.536
R9277 a_50466_25802.n39 a_50466_25802.n38 0.255
R9278 a_50466_25802.n28 a_50466_25802.n27 0.151
R9279 a_50466_25802.n20 a_50466_25802.n19 0.151
R9280 a_50466_25802.n23 a_50466_25802.n22 0.125
R9281 a_50466_25802.n34 a_50466_25802.n32 0.028
R9282 a_50466_25802.n7 a_50466_25802.n5 0.028
R9283 a_50466_25802.n1 a_50466_25802.n0 0.025
R9284 a_50466_25802.n20 a_50466_25802.n15 0.024
R9285 a_50466_25802.n36 a_50466_25802.n34 0.012
R9286 a_50466_25802.n9 a_50466_25802.n7 0.012
R9287 a_50466_25802.n29 a_50466_25802.n23 0.011
R9288 a_50466_25802.n30 a_50466_25802.n29 0.011
R9289 a_50466_25802.n14 a_50466_25802.n10 0.011
R9290 a_50466_25802.n38 a_50466_25802.n37 0.01
R9291 a_50466_25802.n22 a_50466_25802.n21 0.01
R9292 a_50466_25802.n21 a_50466_25802.n14 0.01
R9293 a_50466_25802.n37 a_50466_25802.n30 0.01
R9294 a_41266_65322.n26 a_41266_65322.t1 10.181
R9295 a_41266_65322.n18 a_41266_65322.t2 10.181
R9296 a_41266_65322.t0 a_41266_65322.n39 9.68
R9297 a_41266_65322.n3 a_41266_65322.n2 9.302
R9298 a_41266_65322.n13 a_41266_65322.n12 9.302
R9299 a_41266_65322.n32 a_41266_65322.n31 9.3
R9300 a_41266_65322.n34 a_41266_65322.n33 9.3
R9301 a_41266_65322.n7 a_41266_65322.n6 9.3
R9302 a_41266_65322.n5 a_41266_65322.n4 9.3
R9303 a_41266_65322.n36 a_41266_65322.n35 9
R9304 a_41266_65322.n9 a_41266_65322.n8 9
R9305 a_41266_65322.n27 a_41266_65322.n25 7.729
R9306 a_41266_65322.n19 a_41266_65322.n17 7.729
R9307 a_41266_65322.n27 a_41266_65322.n26 6.296
R9308 a_41266_65322.n19 a_41266_65322.n18 6.296
R9309 a_41266_65322.n30 a_41266_65322.n3 4.508
R9310 a_41266_65322.n14 a_41266_65322.n13 4.508
R9311 a_41266_65322.n37 a_41266_65322.n36 4.496
R9312 a_41266_65322.n21 a_41266_65322.n20 4.496
R9313 a_41266_65322.n29 a_41266_65322.n28 4.495
R9314 a_41266_65322.n10 a_41266_65322.n9 4.495
R9315 a_41266_65322.n14 a_41266_65322.n11 4.494
R9316 a_41266_65322.n30 a_41266_65322.n1 4.494
R9317 a_41266_65322.n39 a_41266_65322.t3 1.087
R9318 a_41266_65322.n25 a_41266_65322.n24 0.536
R9319 a_41266_65322.n17 a_41266_65322.n16 0.536
R9320 a_41266_65322.n39 a_41266_65322.n38 0.255
R9321 a_41266_65322.n28 a_41266_65322.n27 0.151
R9322 a_41266_65322.n20 a_41266_65322.n19 0.151
R9323 a_41266_65322.n23 a_41266_65322.n22 0.125
R9324 a_41266_65322.n34 a_41266_65322.n32 0.028
R9325 a_41266_65322.n7 a_41266_65322.n5 0.028
R9326 a_41266_65322.n1 a_41266_65322.n0 0.025
R9327 a_41266_65322.n20 a_41266_65322.n15 0.024
R9328 a_41266_65322.n36 a_41266_65322.n34 0.012
R9329 a_41266_65322.n9 a_41266_65322.n7 0.012
R9330 a_41266_65322.n29 a_41266_65322.n23 0.011
R9331 a_41266_65322.n30 a_41266_65322.n29 0.011
R9332 a_41266_65322.n14 a_41266_65322.n10 0.011
R9333 a_41266_65322.n38 a_41266_65322.n37 0.01
R9334 a_41266_65322.n22 a_41266_65322.n21 0.01
R9335 a_41266_65322.n21 a_41266_65322.n14 0.01
R9336 a_41266_65322.n37 a_41266_65322.n30 0.01
R9337 a_40976_65246.n10 a_40976_65246.t0 10.181
R9338 a_40976_65246.n10 a_40976_65246.t1 10.181
R9339 a_40976_65246.t2 a_40976_65246.n18 9.68
R9340 a_40976_65246.n1 a_40976_65246.n0 9.302
R9341 a_40976_65246.n7 a_40976_65246.n6 9.3
R9342 a_40976_65246.n5 a_40976_65246.n4 9.3
R9343 a_40976_65246.n9 a_40976_65246.n8 9
R9344 a_40976_65246.n13 a_40976_65246.n12 7.729
R9345 a_40976_65246.n13 a_40976_65246.n10 6.296
R9346 a_40976_65246.n16 a_40976_65246.n1 4.508
R9347 a_40976_65246.n15 a_40976_65246.n14 4.501
R9348 a_40976_65246.n15 a_40976_65246.n9 4.501
R9349 a_40976_65246.n16 a_40976_65246.n3 4.494
R9350 a_40976_65246.n18 a_40976_65246.t3 1.259
R9351 a_40976_65246.n12 a_40976_65246.n11 0.536
R9352 a_40976_65246.n18 a_40976_65246.n17 0.415
R9353 a_40976_65246.n14 a_40976_65246.n13 0.151
R9354 a_40976_65246.n7 a_40976_65246.n5 0.028
R9355 a_40976_65246.n3 a_40976_65246.n2 0.025
R9356 a_40976_65246.n17 a_40976_65246.n16 0.021
R9357 a_40976_65246.n9 a_40976_65246.n7 0.012
R9358 a_40976_65246.n16 a_40976_65246.n15 0.006
R9359 a_68576_65246.n10 a_68576_65246.t1 10.181
R9360 a_68576_65246.n10 a_68576_65246.t0 10.181
R9361 a_68576_65246.t3 a_68576_65246.n18 9.68
R9362 a_68576_65246.n1 a_68576_65246.n0 9.302
R9363 a_68576_65246.n7 a_68576_65246.n6 9.3
R9364 a_68576_65246.n5 a_68576_65246.n4 9.3
R9365 a_68576_65246.n9 a_68576_65246.n8 9
R9366 a_68576_65246.n13 a_68576_65246.n12 7.729
R9367 a_68576_65246.n13 a_68576_65246.n10 6.296
R9368 a_68576_65246.n16 a_68576_65246.n1 4.508
R9369 a_68576_65246.n15 a_68576_65246.n14 4.501
R9370 a_68576_65246.n15 a_68576_65246.n9 4.501
R9371 a_68576_65246.n16 a_68576_65246.n3 4.494
R9372 a_68576_65246.n18 a_68576_65246.t2 1.259
R9373 a_68576_65246.n12 a_68576_65246.n11 0.536
R9374 a_68576_65246.n18 a_68576_65246.n17 0.415
R9375 a_68576_65246.n14 a_68576_65246.n13 0.151
R9376 a_68576_65246.n7 a_68576_65246.n5 0.028
R9377 a_68576_65246.n3 a_68576_65246.n2 0.025
R9378 a_68576_65246.n17 a_68576_65246.n16 0.021
R9379 a_68576_65246.n9 a_68576_65246.n7 0.012
R9380 a_68576_65246.n16 a_68576_65246.n15 0.006
R9381 a_4466_85082.n26 a_4466_85082.t2 10.181
R9382 a_4466_85082.n18 a_4466_85082.t3 10.181
R9383 a_4466_85082.t1 a_4466_85082.n39 9.68
R9384 a_4466_85082.n3 a_4466_85082.n2 9.302
R9385 a_4466_85082.n13 a_4466_85082.n12 9.302
R9386 a_4466_85082.n32 a_4466_85082.n31 9.3
R9387 a_4466_85082.n34 a_4466_85082.n33 9.3
R9388 a_4466_85082.n7 a_4466_85082.n6 9.3
R9389 a_4466_85082.n5 a_4466_85082.n4 9.3
R9390 a_4466_85082.n36 a_4466_85082.n35 9
R9391 a_4466_85082.n9 a_4466_85082.n8 9
R9392 a_4466_85082.n27 a_4466_85082.n25 7.729
R9393 a_4466_85082.n19 a_4466_85082.n17 7.729
R9394 a_4466_85082.n27 a_4466_85082.n26 6.296
R9395 a_4466_85082.n19 a_4466_85082.n18 6.296
R9396 a_4466_85082.n30 a_4466_85082.n3 4.508
R9397 a_4466_85082.n14 a_4466_85082.n13 4.508
R9398 a_4466_85082.n37 a_4466_85082.n36 4.496
R9399 a_4466_85082.n21 a_4466_85082.n20 4.496
R9400 a_4466_85082.n29 a_4466_85082.n28 4.495
R9401 a_4466_85082.n10 a_4466_85082.n9 4.495
R9402 a_4466_85082.n14 a_4466_85082.n11 4.494
R9403 a_4466_85082.n30 a_4466_85082.n1 4.494
R9404 a_4466_85082.n39 a_4466_85082.t0 1.087
R9405 a_4466_85082.n25 a_4466_85082.n24 0.536
R9406 a_4466_85082.n17 a_4466_85082.n16 0.536
R9407 a_4466_85082.n39 a_4466_85082.n38 0.255
R9408 a_4466_85082.n28 a_4466_85082.n27 0.151
R9409 a_4466_85082.n20 a_4466_85082.n19 0.151
R9410 a_4466_85082.n23 a_4466_85082.n22 0.125
R9411 a_4466_85082.n34 a_4466_85082.n32 0.028
R9412 a_4466_85082.n7 a_4466_85082.n5 0.028
R9413 a_4466_85082.n1 a_4466_85082.n0 0.025
R9414 a_4466_85082.n20 a_4466_85082.n15 0.024
R9415 a_4466_85082.n36 a_4466_85082.n34 0.012
R9416 a_4466_85082.n9 a_4466_85082.n7 0.012
R9417 a_4466_85082.n29 a_4466_85082.n23 0.011
R9418 a_4466_85082.n30 a_4466_85082.n29 0.011
R9419 a_4466_85082.n14 a_4466_85082.n10 0.011
R9420 a_4466_85082.n38 a_4466_85082.n37 0.01
R9421 a_4466_85082.n22 a_4466_85082.n21 0.01
R9422 a_4466_85082.n21 a_4466_85082.n14 0.01
R9423 a_4466_85082.n37 a_4466_85082.n30 0.01
R9424 a_59666_25802.n26 a_59666_25802.t1 10.181
R9425 a_59666_25802.n18 a_59666_25802.t0 10.181
R9426 a_59666_25802.t2 a_59666_25802.n39 9.68
R9427 a_59666_25802.n3 a_59666_25802.n2 9.302
R9428 a_59666_25802.n13 a_59666_25802.n12 9.302
R9429 a_59666_25802.n32 a_59666_25802.n31 9.3
R9430 a_59666_25802.n34 a_59666_25802.n33 9.3
R9431 a_59666_25802.n7 a_59666_25802.n6 9.3
R9432 a_59666_25802.n5 a_59666_25802.n4 9.3
R9433 a_59666_25802.n36 a_59666_25802.n35 9
R9434 a_59666_25802.n9 a_59666_25802.n8 9
R9435 a_59666_25802.n27 a_59666_25802.n25 7.729
R9436 a_59666_25802.n19 a_59666_25802.n17 7.729
R9437 a_59666_25802.n27 a_59666_25802.n26 6.296
R9438 a_59666_25802.n19 a_59666_25802.n18 6.296
R9439 a_59666_25802.n30 a_59666_25802.n3 4.508
R9440 a_59666_25802.n14 a_59666_25802.n13 4.508
R9441 a_59666_25802.n37 a_59666_25802.n36 4.496
R9442 a_59666_25802.n21 a_59666_25802.n20 4.496
R9443 a_59666_25802.n29 a_59666_25802.n28 4.495
R9444 a_59666_25802.n10 a_59666_25802.n9 4.495
R9445 a_59666_25802.n14 a_59666_25802.n11 4.494
R9446 a_59666_25802.n30 a_59666_25802.n1 4.494
R9447 a_59666_25802.n39 a_59666_25802.t3 1.087
R9448 a_59666_25802.n25 a_59666_25802.n24 0.536
R9449 a_59666_25802.n17 a_59666_25802.n16 0.536
R9450 a_59666_25802.n39 a_59666_25802.n38 0.255
R9451 a_59666_25802.n28 a_59666_25802.n27 0.151
R9452 a_59666_25802.n20 a_59666_25802.n19 0.151
R9453 a_59666_25802.n23 a_59666_25802.n22 0.125
R9454 a_59666_25802.n34 a_59666_25802.n32 0.028
R9455 a_59666_25802.n7 a_59666_25802.n5 0.028
R9456 a_59666_25802.n1 a_59666_25802.n0 0.025
R9457 a_59666_25802.n20 a_59666_25802.n15 0.024
R9458 a_59666_25802.n36 a_59666_25802.n34 0.012
R9459 a_59666_25802.n9 a_59666_25802.n7 0.012
R9460 a_59666_25802.n29 a_59666_25802.n23 0.011
R9461 a_59666_25802.n30 a_59666_25802.n29 0.011
R9462 a_59666_25802.n14 a_59666_25802.n10 0.011
R9463 a_59666_25802.n38 a_59666_25802.n37 0.01
R9464 a_59666_25802.n22 a_59666_25802.n21 0.01
R9465 a_59666_25802.n21 a_59666_25802.n14 0.01
R9466 a_59666_25802.n37 a_59666_25802.n30 0.01
R9467 a_59376_25726.n10 a_59376_25726.t0 10.181
R9468 a_59376_25726.n10 a_59376_25726.t1 10.181
R9469 a_59376_25726.t3 a_59376_25726.n18 9.68
R9470 a_59376_25726.n1 a_59376_25726.n0 9.302
R9471 a_59376_25726.n7 a_59376_25726.n6 9.3
R9472 a_59376_25726.n5 a_59376_25726.n4 9.3
R9473 a_59376_25726.n9 a_59376_25726.n8 9
R9474 a_59376_25726.n13 a_59376_25726.n12 7.729
R9475 a_59376_25726.n13 a_59376_25726.n10 6.296
R9476 a_59376_25726.n16 a_59376_25726.n1 4.508
R9477 a_59376_25726.n15 a_59376_25726.n14 4.501
R9478 a_59376_25726.n15 a_59376_25726.n9 4.501
R9479 a_59376_25726.n16 a_59376_25726.n3 4.494
R9480 a_59376_25726.n18 a_59376_25726.t2 1.259
R9481 a_59376_25726.n12 a_59376_25726.n11 0.536
R9482 a_59376_25726.n18 a_59376_25726.n17 0.415
R9483 a_59376_25726.n14 a_59376_25726.n13 0.151
R9484 a_59376_25726.n7 a_59376_25726.n5 0.028
R9485 a_59376_25726.n3 a_59376_25726.n2 0.025
R9486 a_59376_25726.n17 a_59376_25726.n16 0.021
R9487 a_59376_25726.n9 a_59376_25726.n7 0.012
R9488 a_59376_25726.n16 a_59376_25726.n15 0.006
R9489 bit1.n14 bit1.t5 552.693
R9490 bit1.n2 bit1.t0 300.446
R9491 bit1.n0 bit1.t3 300.446
R9492 bit1.n11 bit1.t1 300.446
R9493 bit1.n9 bit1.t4 300.446
R9494 bit1.n14 bit1.t2 279.56
R9495 bit1.n15 bit1.n14 120.317
R9496 bit1.n10 bit1.n9 27.537
R9497 bit1.n5 bit1.n2 27.536
R9498 bit1.n1 bit1.n0 24.127
R9499 bit1.n12 bit1.n11 24.127
R9500 bit1.n4 bit1.n3 8.764
R9501 bit1.n8 bit1.n7 8.764
R9502 bit1.n6 bit1.n1 4.662
R9503 bit1.n13 bit1.n12 4.661
R9504 bit1 bit1.n16 4.301
R9505 bit1.n5 bit1.n4 3.401
R9506 bit1.n10 bit1.n8 3.401
R9507 bit1.n13 bit1.n10 0.626
R9508 bit1.n6 bit1.n5 0.626
R9509 bit1.n16 bit1.n15 0.575
R9510 bit1.n16 bit1.n6 0.298
R9511 bit1.n15 bit1.n13 0.298
R9512 a_13376_85006.n10 a_13376_85006.t3 10.181
R9513 a_13376_85006.n10 a_13376_85006.t2 10.181
R9514 a_13376_85006.t0 a_13376_85006.n18 9.68
R9515 a_13376_85006.n1 a_13376_85006.n0 9.302
R9516 a_13376_85006.n7 a_13376_85006.n6 9.3
R9517 a_13376_85006.n5 a_13376_85006.n4 9.3
R9518 a_13376_85006.n9 a_13376_85006.n8 9
R9519 a_13376_85006.n13 a_13376_85006.n12 7.729
R9520 a_13376_85006.n13 a_13376_85006.n10 6.296
R9521 a_13376_85006.n16 a_13376_85006.n1 4.508
R9522 a_13376_85006.n15 a_13376_85006.n14 4.501
R9523 a_13376_85006.n15 a_13376_85006.n9 4.501
R9524 a_13376_85006.n16 a_13376_85006.n3 4.494
R9525 a_13376_85006.n18 a_13376_85006.t1 1.259
R9526 a_13376_85006.n12 a_13376_85006.n11 0.536
R9527 a_13376_85006.n18 a_13376_85006.n17 0.415
R9528 a_13376_85006.n14 a_13376_85006.n13 0.151
R9529 a_13376_85006.n7 a_13376_85006.n5 0.028
R9530 a_13376_85006.n3 a_13376_85006.n2 0.025
R9531 a_13376_85006.n17 a_13376_85006.n16 0.021
R9532 a_13376_85006.n9 a_13376_85006.n7 0.012
R9533 a_13376_85006.n16 a_13376_85006.n15 0.006
R9534 a_13666_85082.n26 a_13666_85082.t2 10.181
R9535 a_13666_85082.n18 a_13666_85082.t1 10.181
R9536 a_13666_85082.t3 a_13666_85082.n39 9.68
R9537 a_13666_85082.n3 a_13666_85082.n2 9.302
R9538 a_13666_85082.n13 a_13666_85082.n12 9.302
R9539 a_13666_85082.n32 a_13666_85082.n31 9.3
R9540 a_13666_85082.n34 a_13666_85082.n33 9.3
R9541 a_13666_85082.n7 a_13666_85082.n6 9.3
R9542 a_13666_85082.n5 a_13666_85082.n4 9.3
R9543 a_13666_85082.n36 a_13666_85082.n35 9
R9544 a_13666_85082.n9 a_13666_85082.n8 9
R9545 a_13666_85082.n27 a_13666_85082.n25 7.729
R9546 a_13666_85082.n19 a_13666_85082.n17 7.729
R9547 a_13666_85082.n27 a_13666_85082.n26 6.296
R9548 a_13666_85082.n19 a_13666_85082.n18 6.296
R9549 a_13666_85082.n30 a_13666_85082.n3 4.508
R9550 a_13666_85082.n14 a_13666_85082.n13 4.508
R9551 a_13666_85082.n37 a_13666_85082.n36 4.496
R9552 a_13666_85082.n21 a_13666_85082.n20 4.496
R9553 a_13666_85082.n29 a_13666_85082.n28 4.495
R9554 a_13666_85082.n10 a_13666_85082.n9 4.495
R9555 a_13666_85082.n14 a_13666_85082.n11 4.494
R9556 a_13666_85082.n30 a_13666_85082.n1 4.494
R9557 a_13666_85082.n39 a_13666_85082.t0 1.087
R9558 a_13666_85082.n25 a_13666_85082.n24 0.536
R9559 a_13666_85082.n17 a_13666_85082.n16 0.536
R9560 a_13666_85082.n39 a_13666_85082.n38 0.255
R9561 a_13666_85082.n28 a_13666_85082.n27 0.151
R9562 a_13666_85082.n20 a_13666_85082.n19 0.151
R9563 a_13666_85082.n23 a_13666_85082.n22 0.125
R9564 a_13666_85082.n34 a_13666_85082.n32 0.028
R9565 a_13666_85082.n7 a_13666_85082.n5 0.028
R9566 a_13666_85082.n1 a_13666_85082.n0 0.025
R9567 a_13666_85082.n20 a_13666_85082.n15 0.024
R9568 a_13666_85082.n36 a_13666_85082.n34 0.012
R9569 a_13666_85082.n9 a_13666_85082.n7 0.012
R9570 a_13666_85082.n29 a_13666_85082.n23 0.011
R9571 a_13666_85082.n30 a_13666_85082.n29 0.011
R9572 a_13666_85082.n14 a_13666_85082.n10 0.011
R9573 a_13666_85082.n38 a_13666_85082.n37 0.01
R9574 a_13666_85082.n22 a_13666_85082.n21 0.01
R9575 a_13666_85082.n21 a_13666_85082.n14 0.01
R9576 a_13666_85082.n37 a_13666_85082.n30 0.01
R9577 a_59376_65246.n10 a_59376_65246.t1 10.181
R9578 a_59376_65246.n10 a_59376_65246.t0 10.181
R9579 a_59376_65246.t3 a_59376_65246.n18 9.68
R9580 a_59376_65246.n1 a_59376_65246.n0 9.302
R9581 a_59376_65246.n7 a_59376_65246.n6 9.3
R9582 a_59376_65246.n5 a_59376_65246.n4 9.3
R9583 a_59376_65246.n9 a_59376_65246.n8 9
R9584 a_59376_65246.n13 a_59376_65246.n12 7.729
R9585 a_59376_65246.n13 a_59376_65246.n10 6.296
R9586 a_59376_65246.n16 a_59376_65246.n1 4.508
R9587 a_59376_65246.n15 a_59376_65246.n14 4.501
R9588 a_59376_65246.n15 a_59376_65246.n9 4.501
R9589 a_59376_65246.n16 a_59376_65246.n3 4.494
R9590 a_59376_65246.n18 a_59376_65246.t2 1.259
R9591 a_59376_65246.n12 a_59376_65246.n11 0.536
R9592 a_59376_65246.n18 a_59376_65246.n17 0.415
R9593 a_59376_65246.n14 a_59376_65246.n13 0.151
R9594 a_59376_65246.n7 a_59376_65246.n5 0.028
R9595 a_59376_65246.n3 a_59376_65246.n2 0.025
R9596 a_59376_65246.n17 a_59376_65246.n16 0.021
R9597 a_59376_65246.n9 a_59376_65246.n7 0.012
R9598 a_59376_65246.n16 a_59376_65246.n15 0.006
R9599 a_4466_15922.n26 a_4466_15922.t2 10.181
R9600 a_4466_15922.n18 a_4466_15922.t1 10.181
R9601 a_4466_15922.t0 a_4466_15922.n39 9.68
R9602 a_4466_15922.n3 a_4466_15922.n2 9.302
R9603 a_4466_15922.n13 a_4466_15922.n12 9.302
R9604 a_4466_15922.n32 a_4466_15922.n31 9.3
R9605 a_4466_15922.n34 a_4466_15922.n33 9.3
R9606 a_4466_15922.n7 a_4466_15922.n6 9.3
R9607 a_4466_15922.n5 a_4466_15922.n4 9.3
R9608 a_4466_15922.n36 a_4466_15922.n35 9
R9609 a_4466_15922.n9 a_4466_15922.n8 9
R9610 a_4466_15922.n27 a_4466_15922.n25 7.729
R9611 a_4466_15922.n19 a_4466_15922.n17 7.729
R9612 a_4466_15922.n27 a_4466_15922.n26 6.296
R9613 a_4466_15922.n19 a_4466_15922.n18 6.296
R9614 a_4466_15922.n30 a_4466_15922.n3 4.508
R9615 a_4466_15922.n14 a_4466_15922.n13 4.508
R9616 a_4466_15922.n37 a_4466_15922.n36 4.496
R9617 a_4466_15922.n21 a_4466_15922.n20 4.496
R9618 a_4466_15922.n29 a_4466_15922.n28 4.495
R9619 a_4466_15922.n10 a_4466_15922.n9 4.495
R9620 a_4466_15922.n14 a_4466_15922.n11 4.494
R9621 a_4466_15922.n30 a_4466_15922.n1 4.494
R9622 a_4466_15922.n39 a_4466_15922.t3 1.087
R9623 a_4466_15922.n25 a_4466_15922.n24 0.536
R9624 a_4466_15922.n17 a_4466_15922.n16 0.536
R9625 a_4466_15922.n39 a_4466_15922.n38 0.255
R9626 a_4466_15922.n28 a_4466_15922.n27 0.151
R9627 a_4466_15922.n20 a_4466_15922.n19 0.151
R9628 a_4466_15922.n23 a_4466_15922.n22 0.125
R9629 a_4466_15922.n34 a_4466_15922.n32 0.028
R9630 a_4466_15922.n7 a_4466_15922.n5 0.028
R9631 a_4466_15922.n1 a_4466_15922.n0 0.025
R9632 a_4466_15922.n20 a_4466_15922.n15 0.024
R9633 a_4466_15922.n36 a_4466_15922.n34 0.012
R9634 a_4466_15922.n9 a_4466_15922.n7 0.012
R9635 a_4466_15922.n29 a_4466_15922.n23 0.011
R9636 a_4466_15922.n30 a_4466_15922.n29 0.011
R9637 a_4466_15922.n14 a_4466_15922.n10 0.011
R9638 a_4466_15922.n38 a_4466_15922.n37 0.01
R9639 a_4466_15922.n22 a_4466_15922.n21 0.01
R9640 a_4466_15922.n21 a_4466_15922.n14 0.01
R9641 a_4466_15922.n37 a_4466_15922.n30 0.01
R9642 a_22866_65322.n26 a_22866_65322.t0 10.181
R9643 a_22866_65322.n18 a_22866_65322.t1 10.181
R9644 a_22866_65322.t3 a_22866_65322.n39 9.68
R9645 a_22866_65322.n3 a_22866_65322.n2 9.302
R9646 a_22866_65322.n13 a_22866_65322.n12 9.302
R9647 a_22866_65322.n32 a_22866_65322.n31 9.3
R9648 a_22866_65322.n34 a_22866_65322.n33 9.3
R9649 a_22866_65322.n7 a_22866_65322.n6 9.3
R9650 a_22866_65322.n5 a_22866_65322.n4 9.3
R9651 a_22866_65322.n36 a_22866_65322.n35 9
R9652 a_22866_65322.n9 a_22866_65322.n8 9
R9653 a_22866_65322.n27 a_22866_65322.n25 7.729
R9654 a_22866_65322.n19 a_22866_65322.n17 7.729
R9655 a_22866_65322.n27 a_22866_65322.n26 6.296
R9656 a_22866_65322.n19 a_22866_65322.n18 6.296
R9657 a_22866_65322.n30 a_22866_65322.n3 4.508
R9658 a_22866_65322.n14 a_22866_65322.n13 4.508
R9659 a_22866_65322.n37 a_22866_65322.n36 4.496
R9660 a_22866_65322.n21 a_22866_65322.n20 4.496
R9661 a_22866_65322.n29 a_22866_65322.n28 4.495
R9662 a_22866_65322.n10 a_22866_65322.n9 4.495
R9663 a_22866_65322.n14 a_22866_65322.n11 4.494
R9664 a_22866_65322.n30 a_22866_65322.n1 4.494
R9665 a_22866_65322.n39 a_22866_65322.t2 1.087
R9666 a_22866_65322.n25 a_22866_65322.n24 0.536
R9667 a_22866_65322.n17 a_22866_65322.n16 0.536
R9668 a_22866_65322.n39 a_22866_65322.n38 0.255
R9669 a_22866_65322.n28 a_22866_65322.n27 0.151
R9670 a_22866_65322.n20 a_22866_65322.n19 0.151
R9671 a_22866_65322.n23 a_22866_65322.n22 0.125
R9672 a_22866_65322.n34 a_22866_65322.n32 0.028
R9673 a_22866_65322.n7 a_22866_65322.n5 0.028
R9674 a_22866_65322.n1 a_22866_65322.n0 0.025
R9675 a_22866_65322.n20 a_22866_65322.n15 0.024
R9676 a_22866_65322.n36 a_22866_65322.n34 0.012
R9677 a_22866_65322.n9 a_22866_65322.n7 0.012
R9678 a_22866_65322.n29 a_22866_65322.n23 0.011
R9679 a_22866_65322.n30 a_22866_65322.n29 0.011
R9680 a_22866_65322.n14 a_22866_65322.n10 0.011
R9681 a_22866_65322.n38 a_22866_65322.n37 0.01
R9682 a_22866_65322.n22 a_22866_65322.n21 0.01
R9683 a_22866_65322.n21 a_22866_65322.n14 0.01
R9684 a_22866_65322.n37 a_22866_65322.n30 0.01
R9685 a_22576_65246.n10 a_22576_65246.t0 10.181
R9686 a_22576_65246.n10 a_22576_65246.t1 10.181
R9687 a_22576_65246.t3 a_22576_65246.n18 9.68
R9688 a_22576_65246.n1 a_22576_65246.n0 9.302
R9689 a_22576_65246.n7 a_22576_65246.n6 9.3
R9690 a_22576_65246.n5 a_22576_65246.n4 9.3
R9691 a_22576_65246.n9 a_22576_65246.n8 9
R9692 a_22576_65246.n13 a_22576_65246.n12 7.729
R9693 a_22576_65246.n13 a_22576_65246.n10 6.296
R9694 a_22576_65246.n16 a_22576_65246.n1 4.508
R9695 a_22576_65246.n15 a_22576_65246.n14 4.501
R9696 a_22576_65246.n15 a_22576_65246.n9 4.501
R9697 a_22576_65246.n16 a_22576_65246.n3 4.494
R9698 a_22576_65246.n18 a_22576_65246.t2 1.259
R9699 a_22576_65246.n12 a_22576_65246.n11 0.536
R9700 a_22576_65246.n18 a_22576_65246.n17 0.415
R9701 a_22576_65246.n14 a_22576_65246.n13 0.151
R9702 a_22576_65246.n7 a_22576_65246.n5 0.028
R9703 a_22576_65246.n3 a_22576_65246.n2 0.025
R9704 a_22576_65246.n17 a_22576_65246.n16 0.021
R9705 a_22576_65246.n9 a_22576_65246.n7 0.012
R9706 a_22576_65246.n16 a_22576_65246.n15 0.006
R9707 a_68866_65322.n26 a_68866_65322.t1 10.181
R9708 a_68866_65322.n18 a_68866_65322.t0 10.181
R9709 a_68866_65322.t2 a_68866_65322.n39 9.68
R9710 a_68866_65322.n3 a_68866_65322.n2 9.302
R9711 a_68866_65322.n13 a_68866_65322.n12 9.302
R9712 a_68866_65322.n32 a_68866_65322.n31 9.3
R9713 a_68866_65322.n34 a_68866_65322.n33 9.3
R9714 a_68866_65322.n7 a_68866_65322.n6 9.3
R9715 a_68866_65322.n5 a_68866_65322.n4 9.3
R9716 a_68866_65322.n36 a_68866_65322.n35 9
R9717 a_68866_65322.n9 a_68866_65322.n8 9
R9718 a_68866_65322.n27 a_68866_65322.n25 7.729
R9719 a_68866_65322.n19 a_68866_65322.n17 7.729
R9720 a_68866_65322.n27 a_68866_65322.n26 6.296
R9721 a_68866_65322.n19 a_68866_65322.n18 6.296
R9722 a_68866_65322.n30 a_68866_65322.n3 4.508
R9723 a_68866_65322.n14 a_68866_65322.n13 4.508
R9724 a_68866_65322.n37 a_68866_65322.n36 4.496
R9725 a_68866_65322.n21 a_68866_65322.n20 4.496
R9726 a_68866_65322.n29 a_68866_65322.n28 4.495
R9727 a_68866_65322.n10 a_68866_65322.n9 4.495
R9728 a_68866_65322.n14 a_68866_65322.n11 4.494
R9729 a_68866_65322.n30 a_68866_65322.n1 4.494
R9730 a_68866_65322.n39 a_68866_65322.t3 1.087
R9731 a_68866_65322.n25 a_68866_65322.n24 0.536
R9732 a_68866_65322.n17 a_68866_65322.n16 0.536
R9733 a_68866_65322.n39 a_68866_65322.n38 0.255
R9734 a_68866_65322.n28 a_68866_65322.n27 0.151
R9735 a_68866_65322.n20 a_68866_65322.n19 0.151
R9736 a_68866_65322.n23 a_68866_65322.n22 0.125
R9737 a_68866_65322.n34 a_68866_65322.n32 0.028
R9738 a_68866_65322.n7 a_68866_65322.n5 0.028
R9739 a_68866_65322.n1 a_68866_65322.n0 0.025
R9740 a_68866_65322.n20 a_68866_65322.n15 0.024
R9741 a_68866_65322.n36 a_68866_65322.n34 0.012
R9742 a_68866_65322.n9 a_68866_65322.n7 0.012
R9743 a_68866_65322.n29 a_68866_65322.n23 0.011
R9744 a_68866_65322.n30 a_68866_65322.n29 0.011
R9745 a_68866_65322.n14 a_68866_65322.n10 0.011
R9746 a_68866_65322.n38 a_68866_65322.n37 0.01
R9747 a_68866_65322.n22 a_68866_65322.n21 0.01
R9748 a_68866_65322.n21 a_68866_65322.n14 0.01
R9749 a_68866_65322.n37 a_68866_65322.n30 0.01
R9750 a_40976_45486.n10 a_40976_45486.t1 10.181
R9751 a_40976_45486.n10 a_40976_45486.t0 10.181
R9752 a_40976_45486.t3 a_40976_45486.n18 9.68
R9753 a_40976_45486.n1 a_40976_45486.n0 9.302
R9754 a_40976_45486.n7 a_40976_45486.n6 9.3
R9755 a_40976_45486.n5 a_40976_45486.n4 9.3
R9756 a_40976_45486.n9 a_40976_45486.n8 9
R9757 a_40976_45486.n13 a_40976_45486.n12 7.729
R9758 a_40976_45486.n13 a_40976_45486.n10 6.296
R9759 a_40976_45486.n16 a_40976_45486.n1 4.508
R9760 a_40976_45486.n15 a_40976_45486.n14 4.501
R9761 a_40976_45486.n15 a_40976_45486.n9 4.501
R9762 a_40976_45486.n16 a_40976_45486.n3 4.494
R9763 a_40976_45486.n18 a_40976_45486.t2 1.259
R9764 a_40976_45486.n12 a_40976_45486.n11 0.536
R9765 a_40976_45486.n18 a_40976_45486.n17 0.415
R9766 a_40976_45486.n14 a_40976_45486.n13 0.151
R9767 a_40976_45486.n7 a_40976_45486.n5 0.028
R9768 a_40976_45486.n3 a_40976_45486.n2 0.025
R9769 a_40976_45486.n17 a_40976_45486.n16 0.021
R9770 a_40976_45486.n9 a_40976_45486.n7 0.012
R9771 a_40976_45486.n16 a_40976_45486.n15 0.006
R9772 a_59376_5966.n10 a_59376_5966.t1 10.181
R9773 a_59376_5966.n10 a_59376_5966.t0 10.181
R9774 a_59376_5966.t3 a_59376_5966.n18 9.68
R9775 a_59376_5966.n1 a_59376_5966.n0 9.302
R9776 a_59376_5966.n7 a_59376_5966.n6 9.3
R9777 a_59376_5966.n5 a_59376_5966.n4 9.3
R9778 a_59376_5966.n9 a_59376_5966.n8 9
R9779 a_59376_5966.n13 a_59376_5966.n12 7.729
R9780 a_59376_5966.n13 a_59376_5966.n10 6.296
R9781 a_59376_5966.n16 a_59376_5966.n1 4.508
R9782 a_59376_5966.n15 a_59376_5966.n14 4.501
R9783 a_59376_5966.n15 a_59376_5966.n9 4.501
R9784 a_59376_5966.n16 a_59376_5966.n3 4.494
R9785 a_59376_5966.n18 a_59376_5966.t2 1.259
R9786 a_59376_5966.n12 a_59376_5966.n11 0.536
R9787 a_59376_5966.n18 a_59376_5966.n17 0.415
R9788 a_59376_5966.n14 a_59376_5966.n13 0.151
R9789 a_59376_5966.n7 a_59376_5966.n5 0.028
R9790 a_59376_5966.n3 a_59376_5966.n2 0.025
R9791 a_59376_5966.n17 a_59376_5966.n16 0.021
R9792 a_59376_5966.n9 a_59376_5966.n7 0.012
R9793 a_59376_5966.n16 a_59376_5966.n15 0.006
R9794 a_31776_75126.n10 a_31776_75126.t1 10.181
R9795 a_31776_75126.n10 a_31776_75126.t2 10.181
R9796 a_31776_75126.t0 a_31776_75126.n18 9.68
R9797 a_31776_75126.n1 a_31776_75126.n0 9.302
R9798 a_31776_75126.n7 a_31776_75126.n6 9.3
R9799 a_31776_75126.n5 a_31776_75126.n4 9.3
R9800 a_31776_75126.n9 a_31776_75126.n8 9
R9801 a_31776_75126.n13 a_31776_75126.n12 7.729
R9802 a_31776_75126.n13 a_31776_75126.n10 6.296
R9803 a_31776_75126.n16 a_31776_75126.n1 4.508
R9804 a_31776_75126.n15 a_31776_75126.n14 4.501
R9805 a_31776_75126.n15 a_31776_75126.n9 4.501
R9806 a_31776_75126.n16 a_31776_75126.n3 4.494
R9807 a_31776_75126.n18 a_31776_75126.t3 1.259
R9808 a_31776_75126.n12 a_31776_75126.n11 0.536
R9809 a_31776_75126.n18 a_31776_75126.n17 0.415
R9810 a_31776_75126.n14 a_31776_75126.n13 0.151
R9811 a_31776_75126.n7 a_31776_75126.n5 0.028
R9812 a_31776_75126.n3 a_31776_75126.n2 0.025
R9813 a_31776_75126.n17 a_31776_75126.n16 0.021
R9814 a_31776_75126.n9 a_31776_75126.n7 0.012
R9815 a_31776_75126.n16 a_31776_75126.n15 0.006
R9816 a_50176_65246.n10 a_50176_65246.t0 10.181
R9817 a_50176_65246.n10 a_50176_65246.t1 10.181
R9818 a_50176_65246.t3 a_50176_65246.n18 9.68
R9819 a_50176_65246.n1 a_50176_65246.n0 9.302
R9820 a_50176_65246.n7 a_50176_65246.n6 9.3
R9821 a_50176_65246.n5 a_50176_65246.n4 9.3
R9822 a_50176_65246.n9 a_50176_65246.n8 9
R9823 a_50176_65246.n13 a_50176_65246.n12 7.729
R9824 a_50176_65246.n13 a_50176_65246.n10 6.296
R9825 a_50176_65246.n16 a_50176_65246.n1 4.508
R9826 a_50176_65246.n15 a_50176_65246.n14 4.501
R9827 a_50176_65246.n15 a_50176_65246.n9 4.501
R9828 a_50176_65246.n16 a_50176_65246.n3 4.494
R9829 a_50176_65246.n18 a_50176_65246.t2 1.259
R9830 a_50176_65246.n12 a_50176_65246.n11 0.536
R9831 a_50176_65246.n18 a_50176_65246.n17 0.415
R9832 a_50176_65246.n14 a_50176_65246.n13 0.151
R9833 a_50176_65246.n7 a_50176_65246.n5 0.028
R9834 a_50176_65246.n3 a_50176_65246.n2 0.025
R9835 a_50176_65246.n17 a_50176_65246.n16 0.021
R9836 a_50176_65246.n9 a_50176_65246.n7 0.012
R9837 a_50176_65246.n16 a_50176_65246.n15 0.006
R9838 a_32066_75202.n26 a_32066_75202.t0 10.181
R9839 a_32066_75202.n18 a_32066_75202.t1 10.181
R9840 a_32066_75202.t3 a_32066_75202.n39 9.68
R9841 a_32066_75202.n3 a_32066_75202.n2 9.302
R9842 a_32066_75202.n13 a_32066_75202.n12 9.302
R9843 a_32066_75202.n32 a_32066_75202.n31 9.3
R9844 a_32066_75202.n34 a_32066_75202.n33 9.3
R9845 a_32066_75202.n7 a_32066_75202.n6 9.3
R9846 a_32066_75202.n5 a_32066_75202.n4 9.3
R9847 a_32066_75202.n36 a_32066_75202.n35 9
R9848 a_32066_75202.n9 a_32066_75202.n8 9
R9849 a_32066_75202.n27 a_32066_75202.n25 7.729
R9850 a_32066_75202.n19 a_32066_75202.n17 7.729
R9851 a_32066_75202.n27 a_32066_75202.n26 6.296
R9852 a_32066_75202.n19 a_32066_75202.n18 6.296
R9853 a_32066_75202.n30 a_32066_75202.n3 4.508
R9854 a_32066_75202.n14 a_32066_75202.n13 4.508
R9855 a_32066_75202.n37 a_32066_75202.n36 4.496
R9856 a_32066_75202.n21 a_32066_75202.n20 4.496
R9857 a_32066_75202.n29 a_32066_75202.n28 4.495
R9858 a_32066_75202.n10 a_32066_75202.n9 4.495
R9859 a_32066_75202.n14 a_32066_75202.n11 4.494
R9860 a_32066_75202.n30 a_32066_75202.n1 4.494
R9861 a_32066_75202.n39 a_32066_75202.t2 1.087
R9862 a_32066_75202.n25 a_32066_75202.n24 0.536
R9863 a_32066_75202.n17 a_32066_75202.n16 0.536
R9864 a_32066_75202.n39 a_32066_75202.n38 0.255
R9865 a_32066_75202.n28 a_32066_75202.n27 0.151
R9866 a_32066_75202.n20 a_32066_75202.n19 0.151
R9867 a_32066_75202.n23 a_32066_75202.n22 0.125
R9868 a_32066_75202.n34 a_32066_75202.n32 0.028
R9869 a_32066_75202.n7 a_32066_75202.n5 0.028
R9870 a_32066_75202.n1 a_32066_75202.n0 0.025
R9871 a_32066_75202.n20 a_32066_75202.n15 0.024
R9872 a_32066_75202.n36 a_32066_75202.n34 0.012
R9873 a_32066_75202.n9 a_32066_75202.n7 0.012
R9874 a_32066_75202.n29 a_32066_75202.n23 0.011
R9875 a_32066_75202.n30 a_32066_75202.n29 0.011
R9876 a_32066_75202.n14 a_32066_75202.n10 0.011
R9877 a_32066_75202.n38 a_32066_75202.n37 0.01
R9878 a_32066_75202.n22 a_32066_75202.n21 0.01
R9879 a_32066_75202.n21 a_32066_75202.n14 0.01
R9880 a_32066_75202.n37 a_32066_75202.n30 0.01
R9881 a_59666_45562.n26 a_59666_45562.t1 10.181
R9882 a_59666_45562.n18 a_59666_45562.t0 10.181
R9883 a_59666_45562.t2 a_59666_45562.n39 9.68
R9884 a_59666_45562.n3 a_59666_45562.n2 9.302
R9885 a_59666_45562.n13 a_59666_45562.n12 9.302
R9886 a_59666_45562.n32 a_59666_45562.n31 9.3
R9887 a_59666_45562.n34 a_59666_45562.n33 9.3
R9888 a_59666_45562.n7 a_59666_45562.n6 9.3
R9889 a_59666_45562.n5 a_59666_45562.n4 9.3
R9890 a_59666_45562.n36 a_59666_45562.n35 9
R9891 a_59666_45562.n9 a_59666_45562.n8 9
R9892 a_59666_45562.n27 a_59666_45562.n25 7.729
R9893 a_59666_45562.n19 a_59666_45562.n17 7.729
R9894 a_59666_45562.n27 a_59666_45562.n26 6.296
R9895 a_59666_45562.n19 a_59666_45562.n18 6.296
R9896 a_59666_45562.n30 a_59666_45562.n3 4.508
R9897 a_59666_45562.n14 a_59666_45562.n13 4.508
R9898 a_59666_45562.n37 a_59666_45562.n36 4.496
R9899 a_59666_45562.n21 a_59666_45562.n20 4.496
R9900 a_59666_45562.n29 a_59666_45562.n28 4.495
R9901 a_59666_45562.n10 a_59666_45562.n9 4.495
R9902 a_59666_45562.n14 a_59666_45562.n11 4.494
R9903 a_59666_45562.n30 a_59666_45562.n1 4.494
R9904 a_59666_45562.n39 a_59666_45562.t3 1.087
R9905 a_59666_45562.n25 a_59666_45562.n24 0.536
R9906 a_59666_45562.n17 a_59666_45562.n16 0.536
R9907 a_59666_45562.n39 a_59666_45562.n38 0.255
R9908 a_59666_45562.n28 a_59666_45562.n27 0.151
R9909 a_59666_45562.n20 a_59666_45562.n19 0.151
R9910 a_59666_45562.n23 a_59666_45562.n22 0.125
R9911 a_59666_45562.n34 a_59666_45562.n32 0.028
R9912 a_59666_45562.n7 a_59666_45562.n5 0.028
R9913 a_59666_45562.n1 a_59666_45562.n0 0.025
R9914 a_59666_45562.n20 a_59666_45562.n15 0.024
R9915 a_59666_45562.n36 a_59666_45562.n34 0.012
R9916 a_59666_45562.n9 a_59666_45562.n7 0.012
R9917 a_59666_45562.n29 a_59666_45562.n23 0.011
R9918 a_59666_45562.n30 a_59666_45562.n29 0.011
R9919 a_59666_45562.n14 a_59666_45562.n10 0.011
R9920 a_59666_45562.n38 a_59666_45562.n37 0.01
R9921 a_59666_45562.n22 a_59666_45562.n21 0.01
R9922 a_59666_45562.n21 a_59666_45562.n14 0.01
R9923 a_59666_45562.n37 a_59666_45562.n30 0.01
R9924 a_68866_25802.n26 a_68866_25802.t1 10.181
R9925 a_68866_25802.n18 a_68866_25802.t2 10.181
R9926 a_68866_25802.t0 a_68866_25802.n39 9.68
R9927 a_68866_25802.n3 a_68866_25802.n2 9.302
R9928 a_68866_25802.n13 a_68866_25802.n12 9.302
R9929 a_68866_25802.n32 a_68866_25802.n31 9.3
R9930 a_68866_25802.n34 a_68866_25802.n33 9.3
R9931 a_68866_25802.n7 a_68866_25802.n6 9.3
R9932 a_68866_25802.n5 a_68866_25802.n4 9.3
R9933 a_68866_25802.n36 a_68866_25802.n35 9
R9934 a_68866_25802.n9 a_68866_25802.n8 9
R9935 a_68866_25802.n27 a_68866_25802.n25 7.729
R9936 a_68866_25802.n19 a_68866_25802.n17 7.729
R9937 a_68866_25802.n27 a_68866_25802.n26 6.296
R9938 a_68866_25802.n19 a_68866_25802.n18 6.296
R9939 a_68866_25802.n30 a_68866_25802.n3 4.508
R9940 a_68866_25802.n14 a_68866_25802.n13 4.508
R9941 a_68866_25802.n37 a_68866_25802.n36 4.496
R9942 a_68866_25802.n21 a_68866_25802.n20 4.496
R9943 a_68866_25802.n29 a_68866_25802.n28 4.495
R9944 a_68866_25802.n10 a_68866_25802.n9 4.495
R9945 a_68866_25802.n14 a_68866_25802.n11 4.494
R9946 a_68866_25802.n30 a_68866_25802.n1 4.494
R9947 a_68866_25802.n39 a_68866_25802.t3 1.087
R9948 a_68866_25802.n25 a_68866_25802.n24 0.536
R9949 a_68866_25802.n17 a_68866_25802.n16 0.536
R9950 a_68866_25802.n39 a_68866_25802.n38 0.255
R9951 a_68866_25802.n28 a_68866_25802.n27 0.151
R9952 a_68866_25802.n20 a_68866_25802.n19 0.151
R9953 a_68866_25802.n23 a_68866_25802.n22 0.125
R9954 a_68866_25802.n34 a_68866_25802.n32 0.028
R9955 a_68866_25802.n7 a_68866_25802.n5 0.028
R9956 a_68866_25802.n1 a_68866_25802.n0 0.025
R9957 a_68866_25802.n20 a_68866_25802.n15 0.024
R9958 a_68866_25802.n36 a_68866_25802.n34 0.012
R9959 a_68866_25802.n9 a_68866_25802.n7 0.012
R9960 a_68866_25802.n29 a_68866_25802.n23 0.011
R9961 a_68866_25802.n30 a_68866_25802.n29 0.011
R9962 a_68866_25802.n14 a_68866_25802.n10 0.011
R9963 a_68866_25802.n38 a_68866_25802.n37 0.01
R9964 a_68866_25802.n22 a_68866_25802.n21 0.01
R9965 a_68866_25802.n21 a_68866_25802.n14 0.01
R9966 a_68866_25802.n37 a_68866_25802.n30 0.01
R9967 a_68576_25726.n10 a_68576_25726.t1 10.181
R9968 a_68576_25726.n10 a_68576_25726.t2 10.181
R9969 a_68576_25726.t0 a_68576_25726.n18 9.68
R9970 a_68576_25726.n1 a_68576_25726.n0 9.302
R9971 a_68576_25726.n7 a_68576_25726.n6 9.3
R9972 a_68576_25726.n5 a_68576_25726.n4 9.3
R9973 a_68576_25726.n9 a_68576_25726.n8 9
R9974 a_68576_25726.n13 a_68576_25726.n12 7.729
R9975 a_68576_25726.n13 a_68576_25726.n10 6.296
R9976 a_68576_25726.n16 a_68576_25726.n1 4.508
R9977 a_68576_25726.n15 a_68576_25726.n14 4.501
R9978 a_68576_25726.n15 a_68576_25726.n9 4.501
R9979 a_68576_25726.n16 a_68576_25726.n3 4.494
R9980 a_68576_25726.n18 a_68576_25726.t3 1.259
R9981 a_68576_25726.n12 a_68576_25726.n11 0.536
R9982 a_68576_25726.n18 a_68576_25726.n17 0.415
R9983 a_68576_25726.n14 a_68576_25726.n13 0.151
R9984 a_68576_25726.n7 a_68576_25726.n5 0.028
R9985 a_68576_25726.n3 a_68576_25726.n2 0.025
R9986 a_68576_25726.n17 a_68576_25726.n16 0.021
R9987 a_68576_25726.n9 a_68576_25726.n7 0.012
R9988 a_68576_25726.n16 a_68576_25726.n15 0.006
R9989 a_n436_84486.t3 a_n436_84486.n3 139.026
R9990 a_n436_84486.n3 a_n436_84486.t2 85.389
R9991 a_n436_84486.n3 a_n436_84486.n2 54.371
R9992 a_n436_84486.n0 a_n436_84486.t5 9.633
R9993 a_n436_84486.n2 a_n436_84486.t1 9.587
R9994 a_n436_84486.n1 a_n436_84486.t4 9.587
R9995 a_n436_84486.n0 a_n436_84486.t0 9.587
R9996 a_n436_84486.n1 a_n436_84486.n0 0.528
R9997 a_n436_84486.n2 a_n436_84486.n1 0.046
R9998 a_40976_5966.n10 a_40976_5966.t1 10.181
R9999 a_40976_5966.n10 a_40976_5966.t0 10.181
R10000 a_40976_5966.t3 a_40976_5966.n18 9.68
R10001 a_40976_5966.n1 a_40976_5966.n0 9.302
R10002 a_40976_5966.n7 a_40976_5966.n6 9.3
R10003 a_40976_5966.n5 a_40976_5966.n4 9.3
R10004 a_40976_5966.n9 a_40976_5966.n8 9
R10005 a_40976_5966.n13 a_40976_5966.n12 7.729
R10006 a_40976_5966.n13 a_40976_5966.n10 6.296
R10007 a_40976_5966.n16 a_40976_5966.n1 4.508
R10008 a_40976_5966.n15 a_40976_5966.n14 4.501
R10009 a_40976_5966.n15 a_40976_5966.n9 4.501
R10010 a_40976_5966.n16 a_40976_5966.n3 4.494
R10011 a_40976_5966.n18 a_40976_5966.t2 1.259
R10012 a_40976_5966.n12 a_40976_5966.n11 0.536
R10013 a_40976_5966.n18 a_40976_5966.n17 0.415
R10014 a_40976_5966.n14 a_40976_5966.n13 0.151
R10015 a_40976_5966.n7 a_40976_5966.n5 0.028
R10016 a_40976_5966.n3 a_40976_5966.n2 0.025
R10017 a_40976_5966.n17 a_40976_5966.n16 0.021
R10018 a_40976_5966.n9 a_40976_5966.n7 0.012
R10019 a_40976_5966.n16 a_40976_5966.n15 0.006
R10020 a_13666_35682.n26 a_13666_35682.t1 10.181
R10021 a_13666_35682.n18 a_13666_35682.t0 10.181
R10022 a_13666_35682.t3 a_13666_35682.n39 9.68
R10023 a_13666_35682.n3 a_13666_35682.n2 9.302
R10024 a_13666_35682.n13 a_13666_35682.n12 9.302
R10025 a_13666_35682.n32 a_13666_35682.n31 9.3
R10026 a_13666_35682.n34 a_13666_35682.n33 9.3
R10027 a_13666_35682.n7 a_13666_35682.n6 9.3
R10028 a_13666_35682.n5 a_13666_35682.n4 9.3
R10029 a_13666_35682.n36 a_13666_35682.n35 9
R10030 a_13666_35682.n9 a_13666_35682.n8 9
R10031 a_13666_35682.n27 a_13666_35682.n25 7.729
R10032 a_13666_35682.n19 a_13666_35682.n17 7.729
R10033 a_13666_35682.n27 a_13666_35682.n26 6.296
R10034 a_13666_35682.n19 a_13666_35682.n18 6.296
R10035 a_13666_35682.n30 a_13666_35682.n3 4.508
R10036 a_13666_35682.n14 a_13666_35682.n13 4.508
R10037 a_13666_35682.n37 a_13666_35682.n36 4.496
R10038 a_13666_35682.n21 a_13666_35682.n20 4.496
R10039 a_13666_35682.n29 a_13666_35682.n28 4.495
R10040 a_13666_35682.n10 a_13666_35682.n9 4.495
R10041 a_13666_35682.n14 a_13666_35682.n11 4.494
R10042 a_13666_35682.n30 a_13666_35682.n1 4.494
R10043 a_13666_35682.n39 a_13666_35682.t2 1.087
R10044 a_13666_35682.n25 a_13666_35682.n24 0.536
R10045 a_13666_35682.n17 a_13666_35682.n16 0.536
R10046 a_13666_35682.n39 a_13666_35682.n38 0.255
R10047 a_13666_35682.n28 a_13666_35682.n27 0.151
R10048 a_13666_35682.n20 a_13666_35682.n19 0.151
R10049 a_13666_35682.n23 a_13666_35682.n22 0.125
R10050 a_13666_35682.n34 a_13666_35682.n32 0.028
R10051 a_13666_35682.n7 a_13666_35682.n5 0.028
R10052 a_13666_35682.n1 a_13666_35682.n0 0.025
R10053 a_13666_35682.n20 a_13666_35682.n15 0.024
R10054 a_13666_35682.n36 a_13666_35682.n34 0.012
R10055 a_13666_35682.n9 a_13666_35682.n7 0.012
R10056 a_13666_35682.n29 a_13666_35682.n23 0.011
R10057 a_13666_35682.n30 a_13666_35682.n29 0.011
R10058 a_13666_35682.n14 a_13666_35682.n10 0.011
R10059 a_13666_35682.n38 a_13666_35682.n37 0.01
R10060 a_13666_35682.n22 a_13666_35682.n21 0.01
R10061 a_13666_35682.n21 a_13666_35682.n14 0.01
R10062 a_13666_35682.n37 a_13666_35682.n30 0.01
R10063 a_41266_6042.n26 a_41266_6042.t2 10.181
R10064 a_41266_6042.n18 a_41266_6042.t1 10.181
R10065 a_41266_6042.t0 a_41266_6042.n39 9.68
R10066 a_41266_6042.n3 a_41266_6042.n2 9.302
R10067 a_41266_6042.n13 a_41266_6042.n12 9.302
R10068 a_41266_6042.n32 a_41266_6042.n31 9.3
R10069 a_41266_6042.n34 a_41266_6042.n33 9.3
R10070 a_41266_6042.n7 a_41266_6042.n6 9.3
R10071 a_41266_6042.n5 a_41266_6042.n4 9.3
R10072 a_41266_6042.n36 a_41266_6042.n35 9
R10073 a_41266_6042.n9 a_41266_6042.n8 9
R10074 a_41266_6042.n27 a_41266_6042.n25 7.729
R10075 a_41266_6042.n19 a_41266_6042.n17 7.729
R10076 a_41266_6042.n27 a_41266_6042.n26 6.296
R10077 a_41266_6042.n19 a_41266_6042.n18 6.296
R10078 a_41266_6042.n30 a_41266_6042.n3 4.508
R10079 a_41266_6042.n14 a_41266_6042.n13 4.508
R10080 a_41266_6042.n37 a_41266_6042.n36 4.496
R10081 a_41266_6042.n21 a_41266_6042.n20 4.496
R10082 a_41266_6042.n29 a_41266_6042.n28 4.495
R10083 a_41266_6042.n10 a_41266_6042.n9 4.495
R10084 a_41266_6042.n14 a_41266_6042.n11 4.494
R10085 a_41266_6042.n30 a_41266_6042.n1 4.494
R10086 a_41266_6042.n39 a_41266_6042.t3 1.087
R10087 a_41266_6042.n25 a_41266_6042.n24 0.536
R10088 a_41266_6042.n17 a_41266_6042.n16 0.536
R10089 a_41266_6042.n39 a_41266_6042.n38 0.255
R10090 a_41266_6042.n28 a_41266_6042.n27 0.151
R10091 a_41266_6042.n20 a_41266_6042.n19 0.151
R10092 a_41266_6042.n23 a_41266_6042.n22 0.125
R10093 a_41266_6042.n34 a_41266_6042.n32 0.028
R10094 a_41266_6042.n7 a_41266_6042.n5 0.028
R10095 a_41266_6042.n1 a_41266_6042.n0 0.025
R10096 a_41266_6042.n20 a_41266_6042.n15 0.024
R10097 a_41266_6042.n36 a_41266_6042.n34 0.012
R10098 a_41266_6042.n9 a_41266_6042.n7 0.012
R10099 a_41266_6042.n29 a_41266_6042.n23 0.011
R10100 a_41266_6042.n30 a_41266_6042.n29 0.011
R10101 a_41266_6042.n14 a_41266_6042.n10 0.011
R10102 a_41266_6042.n38 a_41266_6042.n37 0.01
R10103 a_41266_6042.n22 a_41266_6042.n21 0.01
R10104 a_41266_6042.n21 a_41266_6042.n14 0.01
R10105 a_41266_6042.n37 a_41266_6042.n30 0.01
R10106 a_13666_75202.n26 a_13666_75202.t1 10.181
R10107 a_13666_75202.n18 a_13666_75202.t2 10.181
R10108 a_13666_75202.t0 a_13666_75202.n39 9.68
R10109 a_13666_75202.n3 a_13666_75202.n2 9.302
R10110 a_13666_75202.n13 a_13666_75202.n12 9.302
R10111 a_13666_75202.n32 a_13666_75202.n31 9.3
R10112 a_13666_75202.n34 a_13666_75202.n33 9.3
R10113 a_13666_75202.n7 a_13666_75202.n6 9.3
R10114 a_13666_75202.n5 a_13666_75202.n4 9.3
R10115 a_13666_75202.n36 a_13666_75202.n35 9
R10116 a_13666_75202.n9 a_13666_75202.n8 9
R10117 a_13666_75202.n27 a_13666_75202.n25 7.729
R10118 a_13666_75202.n19 a_13666_75202.n17 7.729
R10119 a_13666_75202.n27 a_13666_75202.n26 6.296
R10120 a_13666_75202.n19 a_13666_75202.n18 6.296
R10121 a_13666_75202.n30 a_13666_75202.n3 4.508
R10122 a_13666_75202.n14 a_13666_75202.n13 4.508
R10123 a_13666_75202.n37 a_13666_75202.n36 4.496
R10124 a_13666_75202.n21 a_13666_75202.n20 4.496
R10125 a_13666_75202.n29 a_13666_75202.n28 4.495
R10126 a_13666_75202.n10 a_13666_75202.n9 4.495
R10127 a_13666_75202.n14 a_13666_75202.n11 4.494
R10128 a_13666_75202.n30 a_13666_75202.n1 4.494
R10129 a_13666_75202.n39 a_13666_75202.t3 1.087
R10130 a_13666_75202.n25 a_13666_75202.n24 0.536
R10131 a_13666_75202.n17 a_13666_75202.n16 0.536
R10132 a_13666_75202.n39 a_13666_75202.n38 0.255
R10133 a_13666_75202.n28 a_13666_75202.n27 0.151
R10134 a_13666_75202.n20 a_13666_75202.n19 0.151
R10135 a_13666_75202.n23 a_13666_75202.n22 0.125
R10136 a_13666_75202.n34 a_13666_75202.n32 0.028
R10137 a_13666_75202.n7 a_13666_75202.n5 0.028
R10138 a_13666_75202.n1 a_13666_75202.n0 0.025
R10139 a_13666_75202.n20 a_13666_75202.n15 0.024
R10140 a_13666_75202.n36 a_13666_75202.n34 0.012
R10141 a_13666_75202.n9 a_13666_75202.n7 0.012
R10142 a_13666_75202.n29 a_13666_75202.n23 0.011
R10143 a_13666_75202.n30 a_13666_75202.n29 0.011
R10144 a_13666_75202.n14 a_13666_75202.n10 0.011
R10145 a_13666_75202.n38 a_13666_75202.n37 0.01
R10146 a_13666_75202.n22 a_13666_75202.n21 0.01
R10147 a_13666_75202.n21 a_13666_75202.n14 0.01
R10148 a_13666_75202.n37 a_13666_75202.n30 0.01
R10149 a_13376_75126.n10 a_13376_75126.t0 10.181
R10150 a_13376_75126.n10 a_13376_75126.t1 10.181
R10151 a_13376_75126.t3 a_13376_75126.n18 9.68
R10152 a_13376_75126.n1 a_13376_75126.n0 9.302
R10153 a_13376_75126.n7 a_13376_75126.n6 9.3
R10154 a_13376_75126.n5 a_13376_75126.n4 9.3
R10155 a_13376_75126.n9 a_13376_75126.n8 9
R10156 a_13376_75126.n13 a_13376_75126.n12 7.729
R10157 a_13376_75126.n13 a_13376_75126.n10 6.296
R10158 a_13376_75126.n16 a_13376_75126.n1 4.508
R10159 a_13376_75126.n15 a_13376_75126.n14 4.501
R10160 a_13376_75126.n15 a_13376_75126.n9 4.501
R10161 a_13376_75126.n16 a_13376_75126.n3 4.494
R10162 a_13376_75126.n18 a_13376_75126.t2 1.259
R10163 a_13376_75126.n12 a_13376_75126.n11 0.536
R10164 a_13376_75126.n18 a_13376_75126.n17 0.415
R10165 a_13376_75126.n14 a_13376_75126.n13 0.151
R10166 a_13376_75126.n7 a_13376_75126.n5 0.028
R10167 a_13376_75126.n3 a_13376_75126.n2 0.025
R10168 a_13376_75126.n17 a_13376_75126.n16 0.021
R10169 a_13376_75126.n9 a_13376_75126.n7 0.012
R10170 a_13376_75126.n16 a_13376_75126.n15 0.006
R10171 a_68866_55442.n26 a_68866_55442.t2 10.181
R10172 a_68866_55442.n18 a_68866_55442.t1 10.181
R10173 a_68866_55442.t0 a_68866_55442.n39 9.68
R10174 a_68866_55442.n3 a_68866_55442.n2 9.302
R10175 a_68866_55442.n13 a_68866_55442.n12 9.302
R10176 a_68866_55442.n32 a_68866_55442.n31 9.3
R10177 a_68866_55442.n34 a_68866_55442.n33 9.3
R10178 a_68866_55442.n7 a_68866_55442.n6 9.3
R10179 a_68866_55442.n5 a_68866_55442.n4 9.3
R10180 a_68866_55442.n36 a_68866_55442.n35 9
R10181 a_68866_55442.n9 a_68866_55442.n8 9
R10182 a_68866_55442.n27 a_68866_55442.n25 7.729
R10183 a_68866_55442.n19 a_68866_55442.n17 7.729
R10184 a_68866_55442.n27 a_68866_55442.n26 6.296
R10185 a_68866_55442.n19 a_68866_55442.n18 6.296
R10186 a_68866_55442.n30 a_68866_55442.n3 4.508
R10187 a_68866_55442.n14 a_68866_55442.n13 4.508
R10188 a_68866_55442.n37 a_68866_55442.n36 4.496
R10189 a_68866_55442.n21 a_68866_55442.n20 4.496
R10190 a_68866_55442.n29 a_68866_55442.n28 4.495
R10191 a_68866_55442.n10 a_68866_55442.n9 4.495
R10192 a_68866_55442.n14 a_68866_55442.n11 4.494
R10193 a_68866_55442.n30 a_68866_55442.n1 4.494
R10194 a_68866_55442.n39 a_68866_55442.t3 1.087
R10195 a_68866_55442.n25 a_68866_55442.n24 0.536
R10196 a_68866_55442.n17 a_68866_55442.n16 0.536
R10197 a_68866_55442.n39 a_68866_55442.n38 0.255
R10198 a_68866_55442.n28 a_68866_55442.n27 0.151
R10199 a_68866_55442.n20 a_68866_55442.n19 0.151
R10200 a_68866_55442.n23 a_68866_55442.n22 0.125
R10201 a_68866_55442.n34 a_68866_55442.n32 0.028
R10202 a_68866_55442.n7 a_68866_55442.n5 0.028
R10203 a_68866_55442.n1 a_68866_55442.n0 0.025
R10204 a_68866_55442.n20 a_68866_55442.n15 0.024
R10205 a_68866_55442.n36 a_68866_55442.n34 0.012
R10206 a_68866_55442.n9 a_68866_55442.n7 0.012
R10207 a_68866_55442.n29 a_68866_55442.n23 0.011
R10208 a_68866_55442.n30 a_68866_55442.n29 0.011
R10209 a_68866_55442.n14 a_68866_55442.n10 0.011
R10210 a_68866_55442.n38 a_68866_55442.n37 0.01
R10211 a_68866_55442.n22 a_68866_55442.n21 0.01
R10212 a_68866_55442.n21 a_68866_55442.n14 0.01
R10213 a_68866_55442.n37 a_68866_55442.n30 0.01
R10214 a_22866_35682.n26 a_22866_35682.t1 10.181
R10215 a_22866_35682.n18 a_22866_35682.t0 10.181
R10216 a_22866_35682.t3 a_22866_35682.n39 9.68
R10217 a_22866_35682.n3 a_22866_35682.n2 9.302
R10218 a_22866_35682.n13 a_22866_35682.n12 9.302
R10219 a_22866_35682.n32 a_22866_35682.n31 9.3
R10220 a_22866_35682.n34 a_22866_35682.n33 9.3
R10221 a_22866_35682.n7 a_22866_35682.n6 9.3
R10222 a_22866_35682.n5 a_22866_35682.n4 9.3
R10223 a_22866_35682.n36 a_22866_35682.n35 9
R10224 a_22866_35682.n9 a_22866_35682.n8 9
R10225 a_22866_35682.n27 a_22866_35682.n25 7.729
R10226 a_22866_35682.n19 a_22866_35682.n17 7.729
R10227 a_22866_35682.n27 a_22866_35682.n26 6.296
R10228 a_22866_35682.n19 a_22866_35682.n18 6.296
R10229 a_22866_35682.n30 a_22866_35682.n3 4.508
R10230 a_22866_35682.n14 a_22866_35682.n13 4.508
R10231 a_22866_35682.n37 a_22866_35682.n36 4.496
R10232 a_22866_35682.n21 a_22866_35682.n20 4.496
R10233 a_22866_35682.n29 a_22866_35682.n28 4.495
R10234 a_22866_35682.n10 a_22866_35682.n9 4.495
R10235 a_22866_35682.n14 a_22866_35682.n11 4.494
R10236 a_22866_35682.n30 a_22866_35682.n1 4.494
R10237 a_22866_35682.n39 a_22866_35682.t2 1.087
R10238 a_22866_35682.n25 a_22866_35682.n24 0.536
R10239 a_22866_35682.n17 a_22866_35682.n16 0.536
R10240 a_22866_35682.n39 a_22866_35682.n38 0.255
R10241 a_22866_35682.n28 a_22866_35682.n27 0.151
R10242 a_22866_35682.n20 a_22866_35682.n19 0.151
R10243 a_22866_35682.n23 a_22866_35682.n22 0.125
R10244 a_22866_35682.n34 a_22866_35682.n32 0.028
R10245 a_22866_35682.n7 a_22866_35682.n5 0.028
R10246 a_22866_35682.n1 a_22866_35682.n0 0.025
R10247 a_22866_35682.n20 a_22866_35682.n15 0.024
R10248 a_22866_35682.n36 a_22866_35682.n34 0.012
R10249 a_22866_35682.n9 a_22866_35682.n7 0.012
R10250 a_22866_35682.n29 a_22866_35682.n23 0.011
R10251 a_22866_35682.n30 a_22866_35682.n29 0.011
R10252 a_22866_35682.n14 a_22866_35682.n10 0.011
R10253 a_22866_35682.n38 a_22866_35682.n37 0.01
R10254 a_22866_35682.n22 a_22866_35682.n21 0.01
R10255 a_22866_35682.n21 a_22866_35682.n14 0.01
R10256 a_22866_35682.n37 a_22866_35682.n30 0.01
R10257 a_13666_45562.n26 a_13666_45562.t1 10.181
R10258 a_13666_45562.n18 a_13666_45562.t0 10.181
R10259 a_13666_45562.t3 a_13666_45562.n39 9.68
R10260 a_13666_45562.n3 a_13666_45562.n2 9.302
R10261 a_13666_45562.n13 a_13666_45562.n12 9.302
R10262 a_13666_45562.n32 a_13666_45562.n31 9.3
R10263 a_13666_45562.n34 a_13666_45562.n33 9.3
R10264 a_13666_45562.n7 a_13666_45562.n6 9.3
R10265 a_13666_45562.n5 a_13666_45562.n4 9.3
R10266 a_13666_45562.n36 a_13666_45562.n35 9
R10267 a_13666_45562.n9 a_13666_45562.n8 9
R10268 a_13666_45562.n27 a_13666_45562.n25 7.729
R10269 a_13666_45562.n19 a_13666_45562.n17 7.729
R10270 a_13666_45562.n27 a_13666_45562.n26 6.296
R10271 a_13666_45562.n19 a_13666_45562.n18 6.296
R10272 a_13666_45562.n30 a_13666_45562.n3 4.508
R10273 a_13666_45562.n14 a_13666_45562.n13 4.508
R10274 a_13666_45562.n37 a_13666_45562.n36 4.496
R10275 a_13666_45562.n21 a_13666_45562.n20 4.496
R10276 a_13666_45562.n29 a_13666_45562.n28 4.495
R10277 a_13666_45562.n10 a_13666_45562.n9 4.495
R10278 a_13666_45562.n14 a_13666_45562.n11 4.494
R10279 a_13666_45562.n30 a_13666_45562.n1 4.494
R10280 a_13666_45562.n39 a_13666_45562.t2 1.087
R10281 a_13666_45562.n25 a_13666_45562.n24 0.536
R10282 a_13666_45562.n17 a_13666_45562.n16 0.536
R10283 a_13666_45562.n39 a_13666_45562.n38 0.255
R10284 a_13666_45562.n28 a_13666_45562.n27 0.151
R10285 a_13666_45562.n20 a_13666_45562.n19 0.151
R10286 a_13666_45562.n23 a_13666_45562.n22 0.125
R10287 a_13666_45562.n34 a_13666_45562.n32 0.028
R10288 a_13666_45562.n7 a_13666_45562.n5 0.028
R10289 a_13666_45562.n1 a_13666_45562.n0 0.025
R10290 a_13666_45562.n20 a_13666_45562.n15 0.024
R10291 a_13666_45562.n36 a_13666_45562.n34 0.012
R10292 a_13666_45562.n9 a_13666_45562.n7 0.012
R10293 a_13666_45562.n29 a_13666_45562.n23 0.011
R10294 a_13666_45562.n30 a_13666_45562.n29 0.011
R10295 a_13666_45562.n14 a_13666_45562.n10 0.011
R10296 a_13666_45562.n38 a_13666_45562.n37 0.01
R10297 a_13666_45562.n22 a_13666_45562.n21 0.01
R10298 a_13666_45562.n21 a_13666_45562.n14 0.01
R10299 a_13666_45562.n37 a_13666_45562.n30 0.01
R10300 a_4466_25802.n26 a_4466_25802.t1 10.181
R10301 a_4466_25802.n18 a_4466_25802.t0 10.181
R10302 a_4466_25802.t2 a_4466_25802.n39 9.68
R10303 a_4466_25802.n3 a_4466_25802.n2 9.302
R10304 a_4466_25802.n13 a_4466_25802.n12 9.302
R10305 a_4466_25802.n32 a_4466_25802.n31 9.3
R10306 a_4466_25802.n34 a_4466_25802.n33 9.3
R10307 a_4466_25802.n7 a_4466_25802.n6 9.3
R10308 a_4466_25802.n5 a_4466_25802.n4 9.3
R10309 a_4466_25802.n36 a_4466_25802.n35 9
R10310 a_4466_25802.n9 a_4466_25802.n8 9
R10311 a_4466_25802.n27 a_4466_25802.n25 7.729
R10312 a_4466_25802.n19 a_4466_25802.n17 7.729
R10313 a_4466_25802.n27 a_4466_25802.n26 6.296
R10314 a_4466_25802.n19 a_4466_25802.n18 6.296
R10315 a_4466_25802.n30 a_4466_25802.n3 4.508
R10316 a_4466_25802.n14 a_4466_25802.n13 4.508
R10317 a_4466_25802.n37 a_4466_25802.n36 4.496
R10318 a_4466_25802.n21 a_4466_25802.n20 4.496
R10319 a_4466_25802.n29 a_4466_25802.n28 4.495
R10320 a_4466_25802.n10 a_4466_25802.n9 4.495
R10321 a_4466_25802.n14 a_4466_25802.n11 4.494
R10322 a_4466_25802.n30 a_4466_25802.n1 4.494
R10323 a_4466_25802.n39 a_4466_25802.t3 1.087
R10324 a_4466_25802.n25 a_4466_25802.n24 0.536
R10325 a_4466_25802.n17 a_4466_25802.n16 0.536
R10326 a_4466_25802.n39 a_4466_25802.n38 0.255
R10327 a_4466_25802.n28 a_4466_25802.n27 0.151
R10328 a_4466_25802.n20 a_4466_25802.n19 0.151
R10329 a_4466_25802.n23 a_4466_25802.n22 0.125
R10330 a_4466_25802.n34 a_4466_25802.n32 0.028
R10331 a_4466_25802.n7 a_4466_25802.n5 0.028
R10332 a_4466_25802.n1 a_4466_25802.n0 0.025
R10333 a_4466_25802.n20 a_4466_25802.n15 0.024
R10334 a_4466_25802.n36 a_4466_25802.n34 0.012
R10335 a_4466_25802.n9 a_4466_25802.n7 0.012
R10336 a_4466_25802.n29 a_4466_25802.n23 0.011
R10337 a_4466_25802.n30 a_4466_25802.n29 0.011
R10338 a_4466_25802.n14 a_4466_25802.n10 0.011
R10339 a_4466_25802.n38 a_4466_25802.n37 0.01
R10340 a_4466_25802.n22 a_4466_25802.n21 0.01
R10341 a_4466_25802.n21 a_4466_25802.n14 0.01
R10342 a_4466_25802.n37 a_4466_25802.n30 0.01
R10343 a_22866_75202.n26 a_22866_75202.t0 10.181
R10344 a_22866_75202.n18 a_22866_75202.t1 10.181
R10345 a_22866_75202.t3 a_22866_75202.n39 9.68
R10346 a_22866_75202.n3 a_22866_75202.n2 9.302
R10347 a_22866_75202.n13 a_22866_75202.n12 9.302
R10348 a_22866_75202.n32 a_22866_75202.n31 9.3
R10349 a_22866_75202.n34 a_22866_75202.n33 9.3
R10350 a_22866_75202.n7 a_22866_75202.n6 9.3
R10351 a_22866_75202.n5 a_22866_75202.n4 9.3
R10352 a_22866_75202.n36 a_22866_75202.n35 9
R10353 a_22866_75202.n9 a_22866_75202.n8 9
R10354 a_22866_75202.n27 a_22866_75202.n25 7.729
R10355 a_22866_75202.n19 a_22866_75202.n17 7.729
R10356 a_22866_75202.n27 a_22866_75202.n26 6.296
R10357 a_22866_75202.n19 a_22866_75202.n18 6.296
R10358 a_22866_75202.n30 a_22866_75202.n3 4.508
R10359 a_22866_75202.n14 a_22866_75202.n13 4.508
R10360 a_22866_75202.n37 a_22866_75202.n36 4.496
R10361 a_22866_75202.n21 a_22866_75202.n20 4.496
R10362 a_22866_75202.n29 a_22866_75202.n28 4.495
R10363 a_22866_75202.n10 a_22866_75202.n9 4.495
R10364 a_22866_75202.n14 a_22866_75202.n11 4.494
R10365 a_22866_75202.n30 a_22866_75202.n1 4.494
R10366 a_22866_75202.n39 a_22866_75202.t2 1.087
R10367 a_22866_75202.n25 a_22866_75202.n24 0.536
R10368 a_22866_75202.n17 a_22866_75202.n16 0.536
R10369 a_22866_75202.n39 a_22866_75202.n38 0.255
R10370 a_22866_75202.n28 a_22866_75202.n27 0.151
R10371 a_22866_75202.n20 a_22866_75202.n19 0.151
R10372 a_22866_75202.n23 a_22866_75202.n22 0.125
R10373 a_22866_75202.n34 a_22866_75202.n32 0.028
R10374 a_22866_75202.n7 a_22866_75202.n5 0.028
R10375 a_22866_75202.n1 a_22866_75202.n0 0.025
R10376 a_22866_75202.n20 a_22866_75202.n15 0.024
R10377 a_22866_75202.n36 a_22866_75202.n34 0.012
R10378 a_22866_75202.n9 a_22866_75202.n7 0.012
R10379 a_22866_75202.n29 a_22866_75202.n23 0.011
R10380 a_22866_75202.n30 a_22866_75202.n29 0.011
R10381 a_22866_75202.n14 a_22866_75202.n10 0.011
R10382 a_22866_75202.n38 a_22866_75202.n37 0.01
R10383 a_22866_75202.n22 a_22866_75202.n21 0.01
R10384 a_22866_75202.n21 a_22866_75202.n14 0.01
R10385 a_22866_75202.n37 a_22866_75202.n30 0.01
R10386 a_22576_75126.n10 a_22576_75126.t1 10.181
R10387 a_22576_75126.n10 a_22576_75126.t2 10.181
R10388 a_22576_75126.t0 a_22576_75126.n18 9.68
R10389 a_22576_75126.n1 a_22576_75126.n0 9.302
R10390 a_22576_75126.n7 a_22576_75126.n6 9.3
R10391 a_22576_75126.n5 a_22576_75126.n4 9.3
R10392 a_22576_75126.n9 a_22576_75126.n8 9
R10393 a_22576_75126.n13 a_22576_75126.n12 7.729
R10394 a_22576_75126.n13 a_22576_75126.n10 6.296
R10395 a_22576_75126.n16 a_22576_75126.n1 4.508
R10396 a_22576_75126.n15 a_22576_75126.n14 4.501
R10397 a_22576_75126.n15 a_22576_75126.n9 4.501
R10398 a_22576_75126.n16 a_22576_75126.n3 4.494
R10399 a_22576_75126.n18 a_22576_75126.t3 1.259
R10400 a_22576_75126.n12 a_22576_75126.n11 0.536
R10401 a_22576_75126.n18 a_22576_75126.n17 0.415
R10402 a_22576_75126.n14 a_22576_75126.n13 0.151
R10403 a_22576_75126.n7 a_22576_75126.n5 0.028
R10404 a_22576_75126.n3 a_22576_75126.n2 0.025
R10405 a_22576_75126.n17 a_22576_75126.n16 0.021
R10406 a_22576_75126.n9 a_22576_75126.n7 0.012
R10407 a_22576_75126.n16 a_22576_75126.n15 0.006
R10408 bit0.n7 bit0.t0 552.693
R10409 bit0.n4 bit0.t1 300.446
R10410 bit0.n2 bit0.t3 300.446
R10411 bit0.n7 bit0.t2 279.56
R10412 bit0.n8 bit0.n7 120.317
R10413 bit0.n3 bit0.n2 27.537
R10414 bit0.n5 bit0.n4 24.127
R10415 bit0.n1 bit0.n0 8.764
R10416 bit0 bit0.n8 4.876
R10417 bit0.n6 bit0.n5 4.661
R10418 bit0.n3 bit0.n1 3.401
R10419 bit0.n6 bit0.n3 0.626
R10420 bit0.n8 bit0.n6 0.298
R10421 VDD.n5 VDD.t8 1362.76
R10422 VDD.n24 VDD.t10 1362.76
R10423 VDD.n43 VDD.t6 1362.76
R10424 VDD.n62 VDD.t0 1362.76
R10425 VDD.n81 VDD.t4 1362.76
R10426 VDD.n100 VDD.t2 1362.76
R10427 VDD.n2 VDD.t9 145.803
R10428 VDD.n21 VDD.t11 145.803
R10429 VDD.n40 VDD.t7 145.803
R10430 VDD.n59 VDD.t1 145.803
R10431 VDD.n78 VDD.t5 145.803
R10432 VDD.n97 VDD.t3 145.803
R10433 VDD.n12 VDD.n11 35.555
R10434 VDD.n31 VDD.n30 35.555
R10435 VDD.n50 VDD.n49 35.555
R10436 VDD.n69 VDD.n68 35.555
R10437 VDD.n88 VDD.n87 35.555
R10438 VDD.n107 VDD.n106 35.555
R10439 VDD.n15 VDD.n14 9.3
R10440 VDD.n1 VDD.n0 9.3
R10441 VDD.n20 VDD.n19 9.3
R10442 VDD.n34 VDD.n33 9.3
R10443 VDD.n39 VDD.n38 9.3
R10444 VDD.n53 VDD.n52 9.3
R10445 VDD.n58 VDD.n57 9.3
R10446 VDD.n72 VDD.n71 9.3
R10447 VDD.n77 VDD.n76 9.3
R10448 VDD.n91 VDD.n90 9.3
R10449 VDD.n96 VDD.n95 9.3
R10450 VDD.n110 VDD.n109 9.3
R10451 VDD.n114 VDD.n113 7.97
R10452 VDD.n118 VDD.n18 5.513
R10453 VDD.n117 VDD.n37 5.513
R10454 VDD.n116 VDD.n56 5.513
R10455 VDD.n115 VDD.n75 5.513
R10456 VDD.n114 VDD.n94 5.513
R10457 VDD.n5 VDD.n4 4.68
R10458 VDD.n24 VDD.n23 4.68
R10459 VDD.n43 VDD.n42 4.68
R10460 VDD.n62 VDD.n61 4.68
R10461 VDD.n81 VDD.n80 4.68
R10462 VDD.n100 VDD.n99 4.68
R10463 VDD.n13 VDD.n3 2.007
R10464 VDD.n32 VDD.n22 2.007
R10465 VDD.n51 VDD.n41 2.007
R10466 VDD.n70 VDD.n60 2.007
R10467 VDD.n89 VDD.n79 2.007
R10468 VDD.n108 VDD.n98 2.007
R10469 VDD.n36 VDD.n20 1.651
R10470 VDD.n55 VDD.n39 1.651
R10471 VDD.n74 VDD.n58 1.651
R10472 VDD.n93 VDD.n77 1.651
R10473 VDD.n112 VDD.n96 1.651
R10474 VDD.n17 VDD.n1 1.65
R10475 VDD.n115 VDD.n114 1.228
R10476 VDD.n15 VDD.n13 1.003
R10477 VDD.n34 VDD.n32 1.003
R10478 VDD.n53 VDD.n51 1.003
R10479 VDD.n72 VDD.n70 1.003
R10480 VDD.n91 VDD.n89 1.003
R10481 VDD.n110 VDD.n108 1.003
R10482 VDD VDD.n118 0.953
R10483 VDD.n118 VDD.n117 0.614
R10484 VDD.n117 VDD.n116 0.614
R10485 VDD.n116 VDD.n115 0.614
R10486 VDD.n16 VDD.n15 0.535
R10487 VDD.n35 VDD.n34 0.533
R10488 VDD.n54 VDD.n53 0.533
R10489 VDD.n73 VDD.n72 0.533
R10490 VDD.n92 VDD.n91 0.533
R10491 VDD.n111 VDD.n110 0.533
R10492 VDD.n8 VDD.n7 0.501
R10493 VDD.n27 VDD.n26 0.501
R10494 VDD.n46 VDD.n45 0.501
R10495 VDD.n65 VDD.n64 0.501
R10496 VDD.n84 VDD.n83 0.501
R10497 VDD.n103 VDD.n102 0.501
R10498 VDD.n3 VDD.n2 0.125
R10499 VDD.n22 VDD.n21 0.125
R10500 VDD.n41 VDD.n40 0.125
R10501 VDD.n60 VDD.n59 0.125
R10502 VDD.n79 VDD.n78 0.125
R10503 VDD.n98 VDD.n97 0.125
R10504 VDD.n18 VDD.n17 0.05
R10505 VDD.n37 VDD.n36 0.049
R10506 VDD.n56 VDD.n55 0.049
R10507 VDD.n75 VDD.n74 0.049
R10508 VDD.n94 VDD.n93 0.049
R10509 VDD.n113 VDD.n112 0.049
R10510 VDD.n7 VDD.n6 0.032
R10511 VDD.n6 VDD.n5 0.032
R10512 VDD.n26 VDD.n25 0.032
R10513 VDD.n25 VDD.n24 0.032
R10514 VDD.n45 VDD.n44 0.032
R10515 VDD.n44 VDD.n43 0.032
R10516 VDD.n64 VDD.n63 0.032
R10517 VDD.n63 VDD.n62 0.032
R10518 VDD.n83 VDD.n82 0.032
R10519 VDD.n82 VDD.n81 0.032
R10520 VDD.n102 VDD.n101 0.032
R10521 VDD.n101 VDD.n100 0.032
R10522 VDD.n12 VDD.n10 0.008
R10523 VDD.n29 VDD.n28 0.008
R10524 VDD.n48 VDD.n47 0.008
R10525 VDD.n67 VDD.n66 0.008
R10526 VDD.n86 VDD.n85 0.008
R10527 VDD.n105 VDD.n104 0.008
R10528 VDD.n10 VDD.n9 0.007
R10529 VDD.n31 VDD.n29 0.007
R10530 VDD.n50 VDD.n48 0.007
R10531 VDD.n69 VDD.n67 0.007
R10532 VDD.n88 VDD.n86 0.007
R10533 VDD.n107 VDD.n105 0.007
R10534 VDD.n9 VDD.n8 0.007
R10535 VDD.n13 VDD.n12 0.007
R10536 VDD.n28 VDD.n27 0.007
R10537 VDD.n32 VDD.n31 0.007
R10538 VDD.n47 VDD.n46 0.007
R10539 VDD.n51 VDD.n50 0.007
R10540 VDD.n66 VDD.n65 0.007
R10541 VDD.n70 VDD.n69 0.007
R10542 VDD.n85 VDD.n84 0.007
R10543 VDD.n89 VDD.n88 0.007
R10544 VDD.n104 VDD.n103 0.007
R10545 VDD.n108 VDD.n107 0.007
R10546 VDD.n36 VDD.n35 0.003
R10547 VDD.n55 VDD.n54 0.003
R10548 VDD.n74 VDD.n73 0.003
R10549 VDD.n93 VDD.n92 0.003
R10550 VDD.n112 VDD.n111 0.003
R10551 VDD.n17 VDD.n16 0.003
R10552 a_32066_35682.n26 a_32066_35682.t1 10.181
R10553 a_32066_35682.n18 a_32066_35682.t0 10.181
R10554 a_32066_35682.t3 a_32066_35682.n39 9.68
R10555 a_32066_35682.n3 a_32066_35682.n2 9.302
R10556 a_32066_35682.n13 a_32066_35682.n12 9.302
R10557 a_32066_35682.n32 a_32066_35682.n31 9.3
R10558 a_32066_35682.n34 a_32066_35682.n33 9.3
R10559 a_32066_35682.n7 a_32066_35682.n6 9.3
R10560 a_32066_35682.n5 a_32066_35682.n4 9.3
R10561 a_32066_35682.n36 a_32066_35682.n35 9
R10562 a_32066_35682.n9 a_32066_35682.n8 9
R10563 a_32066_35682.n27 a_32066_35682.n25 7.729
R10564 a_32066_35682.n19 a_32066_35682.n17 7.729
R10565 a_32066_35682.n27 a_32066_35682.n26 6.296
R10566 a_32066_35682.n19 a_32066_35682.n18 6.296
R10567 a_32066_35682.n30 a_32066_35682.n3 4.508
R10568 a_32066_35682.n14 a_32066_35682.n13 4.508
R10569 a_32066_35682.n37 a_32066_35682.n36 4.496
R10570 a_32066_35682.n21 a_32066_35682.n20 4.496
R10571 a_32066_35682.n29 a_32066_35682.n28 4.495
R10572 a_32066_35682.n10 a_32066_35682.n9 4.495
R10573 a_32066_35682.n14 a_32066_35682.n11 4.494
R10574 a_32066_35682.n30 a_32066_35682.n1 4.494
R10575 a_32066_35682.n39 a_32066_35682.t2 1.087
R10576 a_32066_35682.n25 a_32066_35682.n24 0.536
R10577 a_32066_35682.n17 a_32066_35682.n16 0.536
R10578 a_32066_35682.n39 a_32066_35682.n38 0.255
R10579 a_32066_35682.n28 a_32066_35682.n27 0.151
R10580 a_32066_35682.n20 a_32066_35682.n19 0.151
R10581 a_32066_35682.n23 a_32066_35682.n22 0.125
R10582 a_32066_35682.n34 a_32066_35682.n32 0.028
R10583 a_32066_35682.n7 a_32066_35682.n5 0.028
R10584 a_32066_35682.n1 a_32066_35682.n0 0.025
R10585 a_32066_35682.n20 a_32066_35682.n15 0.024
R10586 a_32066_35682.n36 a_32066_35682.n34 0.012
R10587 a_32066_35682.n9 a_32066_35682.n7 0.012
R10588 a_32066_35682.n29 a_32066_35682.n23 0.011
R10589 a_32066_35682.n30 a_32066_35682.n29 0.011
R10590 a_32066_35682.n14 a_32066_35682.n10 0.011
R10591 a_32066_35682.n38 a_32066_35682.n37 0.01
R10592 a_32066_35682.n22 a_32066_35682.n21 0.01
R10593 a_32066_35682.n21 a_32066_35682.n14 0.01
R10594 a_32066_35682.n37 a_32066_35682.n30 0.01
R10595 a_4176_65246.n10 a_4176_65246.t1 10.181
R10596 a_4176_65246.n10 a_4176_65246.t2 10.181
R10597 a_4176_65246.t0 a_4176_65246.n18 9.68
R10598 a_4176_65246.n1 a_4176_65246.n0 9.302
R10599 a_4176_65246.n7 a_4176_65246.n6 9.3
R10600 a_4176_65246.n5 a_4176_65246.n4 9.3
R10601 a_4176_65246.n9 a_4176_65246.n8 9
R10602 a_4176_65246.n13 a_4176_65246.n12 7.729
R10603 a_4176_65246.n13 a_4176_65246.n10 6.296
R10604 a_4176_65246.n16 a_4176_65246.n1 4.508
R10605 a_4176_65246.n15 a_4176_65246.n14 4.501
R10606 a_4176_65246.n15 a_4176_65246.n9 4.501
R10607 a_4176_65246.n16 a_4176_65246.n3 4.494
R10608 a_4176_65246.n18 a_4176_65246.t3 1.259
R10609 a_4176_65246.n12 a_4176_65246.n11 0.536
R10610 a_4176_65246.n18 a_4176_65246.n17 0.415
R10611 a_4176_65246.n14 a_4176_65246.n13 0.151
R10612 a_4176_65246.n7 a_4176_65246.n5 0.028
R10613 a_4176_65246.n3 a_4176_65246.n2 0.025
R10614 a_4176_65246.n17 a_4176_65246.n16 0.021
R10615 a_4176_65246.n9 a_4176_65246.n7 0.012
R10616 a_4176_65246.n16 a_4176_65246.n15 0.006
R10617 a_31776_5966.n10 a_31776_5966.t2 10.181
R10618 a_31776_5966.n10 a_31776_5966.t1 10.181
R10619 a_31776_5966.t0 a_31776_5966.n18 9.68
R10620 a_31776_5966.n1 a_31776_5966.n0 9.302
R10621 a_31776_5966.n7 a_31776_5966.n6 9.3
R10622 a_31776_5966.n5 a_31776_5966.n4 9.3
R10623 a_31776_5966.n9 a_31776_5966.n8 9
R10624 a_31776_5966.n13 a_31776_5966.n12 7.729
R10625 a_31776_5966.n13 a_31776_5966.n10 6.296
R10626 a_31776_5966.n16 a_31776_5966.n1 4.508
R10627 a_31776_5966.n15 a_31776_5966.n14 4.501
R10628 a_31776_5966.n15 a_31776_5966.n9 4.501
R10629 a_31776_5966.n16 a_31776_5966.n3 4.494
R10630 a_31776_5966.n18 a_31776_5966.t3 1.259
R10631 a_31776_5966.n12 a_31776_5966.n11 0.536
R10632 a_31776_5966.n18 a_31776_5966.n17 0.415
R10633 a_31776_5966.n14 a_31776_5966.n13 0.151
R10634 a_31776_5966.n7 a_31776_5966.n5 0.028
R10635 a_31776_5966.n3 a_31776_5966.n2 0.025
R10636 a_31776_5966.n17 a_31776_5966.n16 0.021
R10637 a_31776_5966.n9 a_31776_5966.n7 0.012
R10638 a_31776_5966.n16 a_31776_5966.n15 0.006
R10639 a_41266_35682.n26 a_41266_35682.t2 10.181
R10640 a_41266_35682.n18 a_41266_35682.t1 10.181
R10641 a_41266_35682.t0 a_41266_35682.n39 9.68
R10642 a_41266_35682.n3 a_41266_35682.n2 9.302
R10643 a_41266_35682.n13 a_41266_35682.n12 9.302
R10644 a_41266_35682.n32 a_41266_35682.n31 9.3
R10645 a_41266_35682.n34 a_41266_35682.n33 9.3
R10646 a_41266_35682.n7 a_41266_35682.n6 9.3
R10647 a_41266_35682.n5 a_41266_35682.n4 9.3
R10648 a_41266_35682.n36 a_41266_35682.n35 9
R10649 a_41266_35682.n9 a_41266_35682.n8 9
R10650 a_41266_35682.n27 a_41266_35682.n25 7.729
R10651 a_41266_35682.n19 a_41266_35682.n17 7.729
R10652 a_41266_35682.n27 a_41266_35682.n26 6.296
R10653 a_41266_35682.n19 a_41266_35682.n18 6.296
R10654 a_41266_35682.n30 a_41266_35682.n3 4.508
R10655 a_41266_35682.n14 a_41266_35682.n13 4.508
R10656 a_41266_35682.n37 a_41266_35682.n36 4.496
R10657 a_41266_35682.n21 a_41266_35682.n20 4.496
R10658 a_41266_35682.n29 a_41266_35682.n28 4.495
R10659 a_41266_35682.n10 a_41266_35682.n9 4.495
R10660 a_41266_35682.n14 a_41266_35682.n11 4.494
R10661 a_41266_35682.n30 a_41266_35682.n1 4.494
R10662 a_41266_35682.n39 a_41266_35682.t3 1.087
R10663 a_41266_35682.n25 a_41266_35682.n24 0.536
R10664 a_41266_35682.n17 a_41266_35682.n16 0.536
R10665 a_41266_35682.n39 a_41266_35682.n38 0.255
R10666 a_41266_35682.n28 a_41266_35682.n27 0.151
R10667 a_41266_35682.n20 a_41266_35682.n19 0.151
R10668 a_41266_35682.n23 a_41266_35682.n22 0.125
R10669 a_41266_35682.n34 a_41266_35682.n32 0.028
R10670 a_41266_35682.n7 a_41266_35682.n5 0.028
R10671 a_41266_35682.n1 a_41266_35682.n0 0.025
R10672 a_41266_35682.n20 a_41266_35682.n15 0.024
R10673 a_41266_35682.n36 a_41266_35682.n34 0.012
R10674 a_41266_35682.n9 a_41266_35682.n7 0.012
R10675 a_41266_35682.n29 a_41266_35682.n23 0.011
R10676 a_41266_35682.n30 a_41266_35682.n29 0.011
R10677 a_41266_35682.n14 a_41266_35682.n10 0.011
R10678 a_41266_35682.n38 a_41266_35682.n37 0.01
R10679 a_41266_35682.n22 a_41266_35682.n21 0.01
R10680 a_41266_35682.n21 a_41266_35682.n14 0.01
R10681 a_41266_35682.n37 a_41266_35682.n30 0.01
R10682 a_31776_15846.n10 a_31776_15846.t0 10.181
R10683 a_31776_15846.n10 a_31776_15846.t1 10.181
R10684 a_31776_15846.t3 a_31776_15846.n18 9.68
R10685 a_31776_15846.n1 a_31776_15846.n0 9.302
R10686 a_31776_15846.n7 a_31776_15846.n6 9.3
R10687 a_31776_15846.n5 a_31776_15846.n4 9.3
R10688 a_31776_15846.n9 a_31776_15846.n8 9
R10689 a_31776_15846.n13 a_31776_15846.n12 7.729
R10690 a_31776_15846.n13 a_31776_15846.n10 6.296
R10691 a_31776_15846.n16 a_31776_15846.n1 4.508
R10692 a_31776_15846.n15 a_31776_15846.n14 4.501
R10693 a_31776_15846.n15 a_31776_15846.n9 4.501
R10694 a_31776_15846.n16 a_31776_15846.n3 4.494
R10695 a_31776_15846.n18 a_31776_15846.t2 1.259
R10696 a_31776_15846.n12 a_31776_15846.n11 0.536
R10697 a_31776_15846.n18 a_31776_15846.n17 0.415
R10698 a_31776_15846.n14 a_31776_15846.n13 0.151
R10699 a_31776_15846.n7 a_31776_15846.n5 0.028
R10700 a_31776_15846.n3 a_31776_15846.n2 0.025
R10701 a_31776_15846.n17 a_31776_15846.n16 0.021
R10702 a_31776_15846.n9 a_31776_15846.n7 0.012
R10703 a_31776_15846.n16 a_31776_15846.n15 0.006
R10704 a_50466_35682.n26 a_50466_35682.t1 10.181
R10705 a_50466_35682.n18 a_50466_35682.t0 10.181
R10706 a_50466_35682.t2 a_50466_35682.n39 9.68
R10707 a_50466_35682.n3 a_50466_35682.n2 9.302
R10708 a_50466_35682.n13 a_50466_35682.n12 9.302
R10709 a_50466_35682.n32 a_50466_35682.n31 9.3
R10710 a_50466_35682.n34 a_50466_35682.n33 9.3
R10711 a_50466_35682.n7 a_50466_35682.n6 9.3
R10712 a_50466_35682.n5 a_50466_35682.n4 9.3
R10713 a_50466_35682.n36 a_50466_35682.n35 9
R10714 a_50466_35682.n9 a_50466_35682.n8 9
R10715 a_50466_35682.n27 a_50466_35682.n25 7.729
R10716 a_50466_35682.n19 a_50466_35682.n17 7.729
R10717 a_50466_35682.n27 a_50466_35682.n26 6.296
R10718 a_50466_35682.n19 a_50466_35682.n18 6.296
R10719 a_50466_35682.n30 a_50466_35682.n3 4.508
R10720 a_50466_35682.n14 a_50466_35682.n13 4.508
R10721 a_50466_35682.n37 a_50466_35682.n36 4.496
R10722 a_50466_35682.n21 a_50466_35682.n20 4.496
R10723 a_50466_35682.n29 a_50466_35682.n28 4.495
R10724 a_50466_35682.n10 a_50466_35682.n9 4.495
R10725 a_50466_35682.n14 a_50466_35682.n11 4.494
R10726 a_50466_35682.n30 a_50466_35682.n1 4.494
R10727 a_50466_35682.n39 a_50466_35682.t3 1.087
R10728 a_50466_35682.n25 a_50466_35682.n24 0.536
R10729 a_50466_35682.n17 a_50466_35682.n16 0.536
R10730 a_50466_35682.n39 a_50466_35682.n38 0.255
R10731 a_50466_35682.n28 a_50466_35682.n27 0.151
R10732 a_50466_35682.n20 a_50466_35682.n19 0.151
R10733 a_50466_35682.n23 a_50466_35682.n22 0.125
R10734 a_50466_35682.n34 a_50466_35682.n32 0.028
R10735 a_50466_35682.n7 a_50466_35682.n5 0.028
R10736 a_50466_35682.n1 a_50466_35682.n0 0.025
R10737 a_50466_35682.n20 a_50466_35682.n15 0.024
R10738 a_50466_35682.n36 a_50466_35682.n34 0.012
R10739 a_50466_35682.n9 a_50466_35682.n7 0.012
R10740 a_50466_35682.n29 a_50466_35682.n23 0.011
R10741 a_50466_35682.n30 a_50466_35682.n29 0.011
R10742 a_50466_35682.n14 a_50466_35682.n10 0.011
R10743 a_50466_35682.n38 a_50466_35682.n37 0.01
R10744 a_50466_35682.n22 a_50466_35682.n21 0.01
R10745 a_50466_35682.n21 a_50466_35682.n14 0.01
R10746 a_50466_35682.n37 a_50466_35682.n30 0.01
R10747 a_59666_65322.n26 a_59666_65322.t2 10.181
R10748 a_59666_65322.n18 a_59666_65322.t1 10.181
R10749 a_59666_65322.t0 a_59666_65322.n39 9.68
R10750 a_59666_65322.n3 a_59666_65322.n2 9.302
R10751 a_59666_65322.n13 a_59666_65322.n12 9.302
R10752 a_59666_65322.n32 a_59666_65322.n31 9.3
R10753 a_59666_65322.n34 a_59666_65322.n33 9.3
R10754 a_59666_65322.n7 a_59666_65322.n6 9.3
R10755 a_59666_65322.n5 a_59666_65322.n4 9.3
R10756 a_59666_65322.n36 a_59666_65322.n35 9
R10757 a_59666_65322.n9 a_59666_65322.n8 9
R10758 a_59666_65322.n27 a_59666_65322.n25 7.729
R10759 a_59666_65322.n19 a_59666_65322.n17 7.729
R10760 a_59666_65322.n27 a_59666_65322.n26 6.296
R10761 a_59666_65322.n19 a_59666_65322.n18 6.296
R10762 a_59666_65322.n30 a_59666_65322.n3 4.508
R10763 a_59666_65322.n14 a_59666_65322.n13 4.508
R10764 a_59666_65322.n37 a_59666_65322.n36 4.496
R10765 a_59666_65322.n21 a_59666_65322.n20 4.496
R10766 a_59666_65322.n29 a_59666_65322.n28 4.495
R10767 a_59666_65322.n10 a_59666_65322.n9 4.495
R10768 a_59666_65322.n14 a_59666_65322.n11 4.494
R10769 a_59666_65322.n30 a_59666_65322.n1 4.494
R10770 a_59666_65322.n39 a_59666_65322.t3 1.087
R10771 a_59666_65322.n25 a_59666_65322.n24 0.536
R10772 a_59666_65322.n17 a_59666_65322.n16 0.536
R10773 a_59666_65322.n39 a_59666_65322.n38 0.255
R10774 a_59666_65322.n28 a_59666_65322.n27 0.151
R10775 a_59666_65322.n20 a_59666_65322.n19 0.151
R10776 a_59666_65322.n23 a_59666_65322.n22 0.125
R10777 a_59666_65322.n34 a_59666_65322.n32 0.028
R10778 a_59666_65322.n7 a_59666_65322.n5 0.028
R10779 a_59666_65322.n1 a_59666_65322.n0 0.025
R10780 a_59666_65322.n20 a_59666_65322.n15 0.024
R10781 a_59666_65322.n36 a_59666_65322.n34 0.012
R10782 a_59666_65322.n9 a_59666_65322.n7 0.012
R10783 a_59666_65322.n29 a_59666_65322.n23 0.011
R10784 a_59666_65322.n30 a_59666_65322.n29 0.011
R10785 a_59666_65322.n14 a_59666_65322.n10 0.011
R10786 a_59666_65322.n38 a_59666_65322.n37 0.01
R10787 a_59666_65322.n22 a_59666_65322.n21 0.01
R10788 a_59666_65322.n21 a_59666_65322.n14 0.01
R10789 a_59666_65322.n37 a_59666_65322.n30 0.01
R10790 a_41266_45562.n26 a_41266_45562.t1 10.181
R10791 a_41266_45562.n18 a_41266_45562.t0 10.181
R10792 a_41266_45562.t2 a_41266_45562.n39 9.68
R10793 a_41266_45562.n3 a_41266_45562.n2 9.302
R10794 a_41266_45562.n13 a_41266_45562.n12 9.302
R10795 a_41266_45562.n32 a_41266_45562.n31 9.3
R10796 a_41266_45562.n34 a_41266_45562.n33 9.3
R10797 a_41266_45562.n7 a_41266_45562.n6 9.3
R10798 a_41266_45562.n5 a_41266_45562.n4 9.3
R10799 a_41266_45562.n36 a_41266_45562.n35 9
R10800 a_41266_45562.n9 a_41266_45562.n8 9
R10801 a_41266_45562.n27 a_41266_45562.n25 7.729
R10802 a_41266_45562.n19 a_41266_45562.n17 7.729
R10803 a_41266_45562.n27 a_41266_45562.n26 6.296
R10804 a_41266_45562.n19 a_41266_45562.n18 6.296
R10805 a_41266_45562.n30 a_41266_45562.n3 4.508
R10806 a_41266_45562.n14 a_41266_45562.n13 4.508
R10807 a_41266_45562.n37 a_41266_45562.n36 4.496
R10808 a_41266_45562.n21 a_41266_45562.n20 4.496
R10809 a_41266_45562.n29 a_41266_45562.n28 4.495
R10810 a_41266_45562.n10 a_41266_45562.n9 4.495
R10811 a_41266_45562.n14 a_41266_45562.n11 4.494
R10812 a_41266_45562.n30 a_41266_45562.n1 4.494
R10813 a_41266_45562.n39 a_41266_45562.t3 1.087
R10814 a_41266_45562.n25 a_41266_45562.n24 0.536
R10815 a_41266_45562.n17 a_41266_45562.n16 0.536
R10816 a_41266_45562.n39 a_41266_45562.n38 0.255
R10817 a_41266_45562.n28 a_41266_45562.n27 0.151
R10818 a_41266_45562.n20 a_41266_45562.n19 0.151
R10819 a_41266_45562.n23 a_41266_45562.n22 0.125
R10820 a_41266_45562.n34 a_41266_45562.n32 0.028
R10821 a_41266_45562.n7 a_41266_45562.n5 0.028
R10822 a_41266_45562.n1 a_41266_45562.n0 0.025
R10823 a_41266_45562.n20 a_41266_45562.n15 0.024
R10824 a_41266_45562.n36 a_41266_45562.n34 0.012
R10825 a_41266_45562.n9 a_41266_45562.n7 0.012
R10826 a_41266_45562.n29 a_41266_45562.n23 0.011
R10827 a_41266_45562.n30 a_41266_45562.n29 0.011
R10828 a_41266_45562.n14 a_41266_45562.n10 0.011
R10829 a_41266_45562.n38 a_41266_45562.n37 0.01
R10830 a_41266_45562.n22 a_41266_45562.n21 0.01
R10831 a_41266_45562.n21 a_41266_45562.n14 0.01
R10832 a_41266_45562.n37 a_41266_45562.n30 0.01
R10833 a_22576_15846.n10 a_22576_15846.t1 10.181
R10834 a_22576_15846.n10 a_22576_15846.t2 10.181
R10835 a_22576_15846.t0 a_22576_15846.n18 9.68
R10836 a_22576_15846.n1 a_22576_15846.n0 9.302
R10837 a_22576_15846.n7 a_22576_15846.n6 9.3
R10838 a_22576_15846.n5 a_22576_15846.n4 9.3
R10839 a_22576_15846.n9 a_22576_15846.n8 9
R10840 a_22576_15846.n13 a_22576_15846.n12 7.729
R10841 a_22576_15846.n13 a_22576_15846.n10 6.296
R10842 a_22576_15846.n16 a_22576_15846.n1 4.508
R10843 a_22576_15846.n15 a_22576_15846.n14 4.501
R10844 a_22576_15846.n15 a_22576_15846.n9 4.501
R10845 a_22576_15846.n16 a_22576_15846.n3 4.494
R10846 a_22576_15846.n18 a_22576_15846.t3 1.259
R10847 a_22576_15846.n12 a_22576_15846.n11 0.536
R10848 a_22576_15846.n18 a_22576_15846.n17 0.415
R10849 a_22576_15846.n14 a_22576_15846.n13 0.151
R10850 a_22576_15846.n7 a_22576_15846.n5 0.028
R10851 a_22576_15846.n3 a_22576_15846.n2 0.025
R10852 a_22576_15846.n17 a_22576_15846.n16 0.021
R10853 a_22576_15846.n9 a_22576_15846.n7 0.012
R10854 a_22576_15846.n16 a_22576_15846.n15 0.006
R10855 a_4176_5966.n10 a_4176_5966.t2 10.181
R10856 a_4176_5966.n10 a_4176_5966.t1 10.181
R10857 a_4176_5966.t0 a_4176_5966.n18 9.68
R10858 a_4176_5966.n1 a_4176_5966.n0 9.302
R10859 a_4176_5966.n7 a_4176_5966.n6 9.3
R10860 a_4176_5966.n5 a_4176_5966.n4 9.3
R10861 a_4176_5966.n9 a_4176_5966.n8 9
R10862 a_4176_5966.n13 a_4176_5966.n12 7.729
R10863 a_4176_5966.n13 a_4176_5966.n10 6.296
R10864 a_4176_5966.n16 a_4176_5966.n1 4.508
R10865 a_4176_5966.n15 a_4176_5966.n14 4.501
R10866 a_4176_5966.n15 a_4176_5966.n9 4.501
R10867 a_4176_5966.n16 a_4176_5966.n3 4.494
R10868 a_4176_5966.n18 a_4176_5966.t3 1.259
R10869 a_4176_5966.n12 a_4176_5966.n11 0.536
R10870 a_4176_5966.n18 a_4176_5966.n17 0.415
R10871 a_4176_5966.n14 a_4176_5966.n13 0.151
R10872 a_4176_5966.n7 a_4176_5966.n5 0.028
R10873 a_4176_5966.n3 a_4176_5966.n2 0.025
R10874 a_4176_5966.n17 a_4176_5966.n16 0.021
R10875 a_4176_5966.n9 a_4176_5966.n7 0.012
R10876 a_4176_5966.n16 a_4176_5966.n15 0.006
C21 OUT_P GND 575.40fF
C22 OUT_N GND 576.12fF
C23 bit5 GND 460.90fF
C24 bit4 GND 229.48fF
C25 bit3 GND 125.29fF
C26 bit2 GND 148.13fF
C27 bit1 GND 157.90fF
C28 bit0 GND 162.36fF
C29 VDD GND 146.97fF
C30 a_4176_5966.n0 GND 0.01fF
C31 a_4176_5966.n1 GND 0.01fF
C32 a_4176_5966.n2 GND 0.00fF
C33 a_4176_5966.n3 GND 0.00fF
C34 a_4176_5966.n4 GND 0.00fF
C35 a_4176_5966.n5 GND 0.00fF
C36 a_4176_5966.n6 GND 0.00fF
C37 a_4176_5966.n7 GND 0.00fF
C38 a_4176_5966.n8 GND 0.00fF
C39 a_4176_5966.n9 GND 0.00fF
C40 a_4176_5966.t2 GND 0.02fF $ **FLOATING
C41 a_4176_5966.t1 GND 0.02fF $ **FLOATING
C42 a_4176_5966.n10 GND 0.05fF
C43 a_4176_5966.n11 GND 0.00fF
C44 a_4176_5966.n12 GND 0.00fF
C45 a_4176_5966.n13 GND 0.02fF
C46 a_4176_5966.n14 GND 0.04fF
C47 a_4176_5966.n15 GND 0.12fF
C48 a_4176_5966.n16 GND 0.01fF
C49 a_4176_5966.n17 GND 0.12fF
C50 a_4176_5966.t3 GND 3.87fF $ **FLOATING
C51 a_4176_5966.n18 GND 0.52fF
C52 a_4176_5966.t0 GND 0.24fF $ **FLOATING
C53 a_22576_15846.n0 GND 0.01fF
C54 a_22576_15846.n1 GND 0.01fF
C55 a_22576_15846.n2 GND 0.00fF
C56 a_22576_15846.n3 GND 0.00fF
C57 a_22576_15846.n4 GND 0.00fF
C58 a_22576_15846.n5 GND 0.00fF
C59 a_22576_15846.n6 GND 0.00fF
C60 a_22576_15846.n7 GND 0.00fF
C61 a_22576_15846.n8 GND 0.00fF
C62 a_22576_15846.n9 GND 0.00fF
C63 a_22576_15846.t1 GND 0.02fF $ **FLOATING
C64 a_22576_15846.t2 GND 0.02fF $ **FLOATING
C65 a_22576_15846.n10 GND 0.05fF
C66 a_22576_15846.n11 GND 0.00fF
C67 a_22576_15846.n12 GND 0.00fF
C68 a_22576_15846.n13 GND 0.02fF
C69 a_22576_15846.n14 GND 0.04fF
C70 a_22576_15846.n15 GND 0.12fF
C71 a_22576_15846.n16 GND 0.01fF
C72 a_22576_15846.n17 GND 0.12fF
C73 a_22576_15846.t3 GND 3.87fF $ **FLOATING
C74 a_22576_15846.n18 GND 0.52fF
C75 a_22576_15846.t0 GND 0.24fF $ **FLOATING
C76 a_41266_45562.n0 GND 0.00fF
C77 a_41266_45562.n1 GND 0.00fF
C78 a_41266_45562.n2 GND 0.01fF
C79 a_41266_45562.n3 GND 0.01fF
C80 a_41266_45562.n4 GND 0.00fF
C81 a_41266_45562.n5 GND 0.00fF
C82 a_41266_45562.n6 GND 0.00fF
C83 a_41266_45562.n7 GND 0.00fF
C84 a_41266_45562.n8 GND 0.00fF
C85 a_41266_45562.n9 GND 0.00fF
C86 a_41266_45562.n10 GND 0.09fF
C87 a_41266_45562.n11 GND 0.00fF
C88 a_41266_45562.n12 GND 0.01fF
C89 a_41266_45562.n13 GND 0.01fF
C90 a_41266_45562.n14 GND 0.01fF
C91 a_41266_45562.n15 GND 0.00fF
C92 a_41266_45562.n16 GND 0.00fF
C93 a_41266_45562.n17 GND 0.00fF
C94 a_41266_45562.t0 GND 0.02fF $ **FLOATING
C95 a_41266_45562.n18 GND 0.07fF
C96 a_41266_45562.n19 GND 0.02fF
C97 a_41266_45562.n20 GND 0.05fF
C98 a_41266_45562.n22 GND 0.04fF
C99 a_41266_45562.n23 GND 0.04fF
C100 a_41266_45562.n24 GND 0.00fF
C101 a_41266_45562.n25 GND 0.00fF
C102 a_41266_45562.t1 GND 0.02fF $ **FLOATING
C103 a_41266_45562.n26 GND 0.07fF
C104 a_41266_45562.n27 GND 0.02fF
C105 a_41266_45562.n28 GND 0.05fF
C106 a_41266_45562.n30 GND 0.01fF
C107 a_41266_45562.n31 GND 0.00fF
C108 a_41266_45562.n32 GND 0.00fF
C109 a_41266_45562.n33 GND 0.00fF
C110 a_41266_45562.n34 GND 0.00fF
C111 a_41266_45562.n35 GND 0.00fF
C112 a_41266_45562.n36 GND 0.00fF
C113 a_41266_45562.n38 GND 0.08fF
C114 a_41266_45562.t3 GND 4.19fF $ **FLOATING
C115 a_41266_45562.n39 GND 0.61fF
C116 a_41266_45562.t2 GND 0.26fF $ **FLOATING
C117 a_59666_65322.n0 GND 0.00fF
C118 a_59666_65322.n1 GND 0.00fF
C119 a_59666_65322.n2 GND 0.01fF
C120 a_59666_65322.n3 GND 0.01fF
C121 a_59666_65322.n4 GND 0.00fF
C122 a_59666_65322.n5 GND 0.00fF
C123 a_59666_65322.n6 GND 0.00fF
C124 a_59666_65322.n7 GND 0.00fF
C125 a_59666_65322.n8 GND 0.00fF
C126 a_59666_65322.n9 GND 0.00fF
C127 a_59666_65322.n10 GND 0.09fF
C128 a_59666_65322.n11 GND 0.00fF
C129 a_59666_65322.n12 GND 0.01fF
C130 a_59666_65322.n13 GND 0.01fF
C131 a_59666_65322.n14 GND 0.01fF
C132 a_59666_65322.n15 GND 0.00fF
C133 a_59666_65322.n16 GND 0.00fF
C134 a_59666_65322.n17 GND 0.00fF
C135 a_59666_65322.t1 GND 0.02fF $ **FLOATING
C136 a_59666_65322.n18 GND 0.07fF
C137 a_59666_65322.n19 GND 0.02fF
C138 a_59666_65322.n20 GND 0.05fF
C139 a_59666_65322.n22 GND 0.04fF
C140 a_59666_65322.n23 GND 0.04fF
C141 a_59666_65322.n24 GND 0.00fF
C142 a_59666_65322.n25 GND 0.00fF
C143 a_59666_65322.t2 GND 0.02fF $ **FLOATING
C144 a_59666_65322.n26 GND 0.07fF
C145 a_59666_65322.n27 GND 0.02fF
C146 a_59666_65322.n28 GND 0.05fF
C147 a_59666_65322.n30 GND 0.01fF
C148 a_59666_65322.n31 GND 0.00fF
C149 a_59666_65322.n32 GND 0.00fF
C150 a_59666_65322.n33 GND 0.00fF
C151 a_59666_65322.n34 GND 0.00fF
C152 a_59666_65322.n35 GND 0.00fF
C153 a_59666_65322.n36 GND 0.00fF
C154 a_59666_65322.n38 GND 0.08fF
C155 a_59666_65322.t3 GND 4.19fF $ **FLOATING
C156 a_59666_65322.n39 GND 0.61fF
C157 a_59666_65322.t0 GND 0.26fF $ **FLOATING
C158 a_50466_35682.n0 GND 0.00fF
C159 a_50466_35682.n1 GND 0.00fF
C160 a_50466_35682.n2 GND 0.01fF
C161 a_50466_35682.n3 GND 0.01fF
C162 a_50466_35682.n4 GND 0.00fF
C163 a_50466_35682.n5 GND 0.00fF
C164 a_50466_35682.n6 GND 0.00fF
C165 a_50466_35682.n7 GND 0.00fF
C166 a_50466_35682.n8 GND 0.00fF
C167 a_50466_35682.n9 GND 0.00fF
C168 a_50466_35682.n10 GND 0.09fF
C169 a_50466_35682.n11 GND 0.00fF
C170 a_50466_35682.n12 GND 0.01fF
C171 a_50466_35682.n13 GND 0.01fF
C172 a_50466_35682.n14 GND 0.01fF
C173 a_50466_35682.n15 GND 0.00fF
C174 a_50466_35682.n16 GND 0.00fF
C175 a_50466_35682.n17 GND 0.00fF
C176 a_50466_35682.t0 GND 0.02fF $ **FLOATING
C177 a_50466_35682.n18 GND 0.07fF
C178 a_50466_35682.n19 GND 0.02fF
C179 a_50466_35682.n20 GND 0.05fF
C180 a_50466_35682.n22 GND 0.04fF
C181 a_50466_35682.n23 GND 0.04fF
C182 a_50466_35682.n24 GND 0.00fF
C183 a_50466_35682.n25 GND 0.00fF
C184 a_50466_35682.t1 GND 0.02fF $ **FLOATING
C185 a_50466_35682.n26 GND 0.07fF
C186 a_50466_35682.n27 GND 0.02fF
C187 a_50466_35682.n28 GND 0.05fF
C188 a_50466_35682.n30 GND 0.01fF
C189 a_50466_35682.n31 GND 0.00fF
C190 a_50466_35682.n32 GND 0.00fF
C191 a_50466_35682.n33 GND 0.00fF
C192 a_50466_35682.n34 GND 0.00fF
C193 a_50466_35682.n35 GND 0.00fF
C194 a_50466_35682.n36 GND 0.00fF
C195 a_50466_35682.n38 GND 0.08fF
C196 a_50466_35682.t3 GND 4.19fF $ **FLOATING
C197 a_50466_35682.n39 GND 0.61fF
C198 a_50466_35682.t2 GND 0.26fF $ **FLOATING
C199 a_31776_15846.n0 GND 0.01fF
C200 a_31776_15846.n1 GND 0.01fF
C201 a_31776_15846.n2 GND 0.00fF
C202 a_31776_15846.n3 GND 0.00fF
C203 a_31776_15846.n4 GND 0.00fF
C204 a_31776_15846.n5 GND 0.00fF
C205 a_31776_15846.n6 GND 0.00fF
C206 a_31776_15846.n7 GND 0.00fF
C207 a_31776_15846.n8 GND 0.00fF
C208 a_31776_15846.n9 GND 0.00fF
C209 a_31776_15846.t0 GND 0.02fF $ **FLOATING
C210 a_31776_15846.t1 GND 0.02fF $ **FLOATING
C211 a_31776_15846.n10 GND 0.05fF
C212 a_31776_15846.n11 GND 0.00fF
C213 a_31776_15846.n12 GND 0.00fF
C214 a_31776_15846.n13 GND 0.02fF
C215 a_31776_15846.n14 GND 0.04fF
C216 a_31776_15846.n15 GND 0.12fF
C217 a_31776_15846.n16 GND 0.01fF
C218 a_31776_15846.n17 GND 0.12fF
C219 a_31776_15846.t2 GND 3.87fF $ **FLOATING
C220 a_31776_15846.n18 GND 0.52fF
C221 a_31776_15846.t3 GND 0.24fF $ **FLOATING
C222 a_41266_35682.n0 GND 0.00fF
C223 a_41266_35682.n1 GND 0.00fF
C224 a_41266_35682.n2 GND 0.01fF
C225 a_41266_35682.n3 GND 0.01fF
C226 a_41266_35682.n4 GND 0.00fF
C227 a_41266_35682.n5 GND 0.00fF
C228 a_41266_35682.n6 GND 0.00fF
C229 a_41266_35682.n7 GND 0.00fF
C230 a_41266_35682.n8 GND 0.00fF
C231 a_41266_35682.n9 GND 0.00fF
C232 a_41266_35682.n10 GND 0.09fF
C233 a_41266_35682.n11 GND 0.00fF
C234 a_41266_35682.n12 GND 0.01fF
C235 a_41266_35682.n13 GND 0.01fF
C236 a_41266_35682.n14 GND 0.01fF
C237 a_41266_35682.n15 GND 0.00fF
C238 a_41266_35682.n16 GND 0.00fF
C239 a_41266_35682.n17 GND 0.00fF
C240 a_41266_35682.t1 GND 0.02fF $ **FLOATING
C241 a_41266_35682.n18 GND 0.07fF
C242 a_41266_35682.n19 GND 0.02fF
C243 a_41266_35682.n20 GND 0.05fF
C244 a_41266_35682.n22 GND 0.04fF
C245 a_41266_35682.n23 GND 0.04fF
C246 a_41266_35682.n24 GND 0.00fF
C247 a_41266_35682.n25 GND 0.00fF
C248 a_41266_35682.t2 GND 0.02fF $ **FLOATING
C249 a_41266_35682.n26 GND 0.07fF
C250 a_41266_35682.n27 GND 0.02fF
C251 a_41266_35682.n28 GND 0.05fF
C252 a_41266_35682.n30 GND 0.01fF
C253 a_41266_35682.n31 GND 0.00fF
C254 a_41266_35682.n32 GND 0.00fF
C255 a_41266_35682.n33 GND 0.00fF
C256 a_41266_35682.n34 GND 0.00fF
C257 a_41266_35682.n35 GND 0.00fF
C258 a_41266_35682.n36 GND 0.00fF
C259 a_41266_35682.n38 GND 0.08fF
C260 a_41266_35682.t3 GND 4.19fF $ **FLOATING
C261 a_41266_35682.n39 GND 0.61fF
C262 a_41266_35682.t0 GND 0.26fF $ **FLOATING
C263 a_31776_5966.n0 GND 0.01fF
C264 a_31776_5966.n1 GND 0.01fF
C265 a_31776_5966.n2 GND 0.00fF
C266 a_31776_5966.n3 GND 0.00fF
C267 a_31776_5966.n4 GND 0.00fF
C268 a_31776_5966.n5 GND 0.00fF
C269 a_31776_5966.n6 GND 0.00fF
C270 a_31776_5966.n7 GND 0.00fF
C271 a_31776_5966.n8 GND 0.00fF
C272 a_31776_5966.n9 GND 0.00fF
C273 a_31776_5966.t2 GND 0.02fF $ **FLOATING
C274 a_31776_5966.t1 GND 0.02fF $ **FLOATING
C275 a_31776_5966.n10 GND 0.05fF
C276 a_31776_5966.n11 GND 0.00fF
C277 a_31776_5966.n12 GND 0.00fF
C278 a_31776_5966.n13 GND 0.02fF
C279 a_31776_5966.n14 GND 0.04fF
C280 a_31776_5966.n15 GND 0.12fF
C281 a_31776_5966.n16 GND 0.01fF
C282 a_31776_5966.n17 GND 0.12fF
C283 a_31776_5966.t3 GND 3.87fF $ **FLOATING
C284 a_31776_5966.n18 GND 0.52fF
C285 a_31776_5966.t0 GND 0.24fF $ **FLOATING
C286 a_4176_65246.n0 GND 0.01fF
C287 a_4176_65246.n1 GND 0.01fF
C288 a_4176_65246.n2 GND 0.00fF
C289 a_4176_65246.n3 GND 0.00fF
C290 a_4176_65246.n4 GND 0.00fF
C291 a_4176_65246.n5 GND 0.00fF
C292 a_4176_65246.n6 GND 0.00fF
C293 a_4176_65246.n7 GND 0.00fF
C294 a_4176_65246.n8 GND 0.00fF
C295 a_4176_65246.n9 GND 0.00fF
C296 a_4176_65246.t1 GND 0.02fF $ **FLOATING
C297 a_4176_65246.t2 GND 0.02fF $ **FLOATING
C298 a_4176_65246.n10 GND 0.05fF
C299 a_4176_65246.n11 GND 0.00fF
C300 a_4176_65246.n12 GND 0.00fF
C301 a_4176_65246.n13 GND 0.02fF
C302 a_4176_65246.n14 GND 0.04fF
C303 a_4176_65246.n15 GND 0.12fF
C304 a_4176_65246.n16 GND 0.01fF
C305 a_4176_65246.n17 GND 0.12fF
C306 a_4176_65246.t3 GND 3.87fF $ **FLOATING
C307 a_4176_65246.n18 GND 0.52fF
C308 a_4176_65246.t0 GND 0.24fF $ **FLOATING
C309 a_32066_35682.n0 GND 0.00fF
C310 a_32066_35682.n1 GND 0.00fF
C311 a_32066_35682.n2 GND 0.01fF
C312 a_32066_35682.n3 GND 0.01fF
C313 a_32066_35682.n4 GND 0.00fF
C314 a_32066_35682.n5 GND 0.00fF
C315 a_32066_35682.n6 GND 0.00fF
C316 a_32066_35682.n7 GND 0.00fF
C317 a_32066_35682.n8 GND 0.00fF
C318 a_32066_35682.n9 GND 0.00fF
C319 a_32066_35682.n10 GND 0.09fF
C320 a_32066_35682.n11 GND 0.00fF
C321 a_32066_35682.n12 GND 0.01fF
C322 a_32066_35682.n13 GND 0.01fF
C323 a_32066_35682.n14 GND 0.01fF
C324 a_32066_35682.n15 GND 0.00fF
C325 a_32066_35682.n16 GND 0.00fF
C326 a_32066_35682.n17 GND 0.00fF
C327 a_32066_35682.t0 GND 0.02fF $ **FLOATING
C328 a_32066_35682.n18 GND 0.07fF
C329 a_32066_35682.n19 GND 0.02fF
C330 a_32066_35682.n20 GND 0.05fF
C331 a_32066_35682.n22 GND 0.04fF
C332 a_32066_35682.n23 GND 0.04fF
C333 a_32066_35682.n24 GND 0.00fF
C334 a_32066_35682.n25 GND 0.00fF
C335 a_32066_35682.t1 GND 0.02fF $ **FLOATING
C336 a_32066_35682.n26 GND 0.07fF
C337 a_32066_35682.n27 GND 0.02fF
C338 a_32066_35682.n28 GND 0.05fF
C339 a_32066_35682.n30 GND 0.01fF
C340 a_32066_35682.n31 GND 0.00fF
C341 a_32066_35682.n32 GND 0.00fF
C342 a_32066_35682.n33 GND 0.00fF
C343 a_32066_35682.n34 GND 0.00fF
C344 a_32066_35682.n35 GND 0.00fF
C345 a_32066_35682.n36 GND 0.00fF
C346 a_32066_35682.n38 GND 0.08fF
C347 a_32066_35682.t2 GND 4.19fF $ **FLOATING
C348 a_32066_35682.n39 GND 0.61fF
C349 a_32066_35682.t3 GND 0.26fF $ **FLOATING
C350 VDD.n0 GND 0.00fF
C351 VDD.n1 GND 0.00fF
C352 VDD.t9 GND 0.05fF $ **FLOATING
C353 VDD.n2 GND 0.01fF
C354 VDD.n3 GND 0.00fF
C355 VDD.t8 GND 0.11fF $ **FLOATING
C356 VDD.n5 GND 0.04fF
C357 VDD.n6 GND 0.00fF
C358 VDD.n7 GND 0.00fF
C359 VDD.n8 GND 0.00fF
C360 VDD.n9 GND 0.00fF
C361 VDD.n10 GND 0.01fF
C362 VDD.n11 GND 0.00fF
C363 VDD.n12 GND 0.00fF
C364 VDD.n13 GND 0.00fF
C365 VDD.n14 GND 0.00fF
C366 VDD.n15 GND 0.00fF
C367 VDD.n16 GND 0.03fF
C368 VDD.n17 GND 0.00fF
C369 VDD.n18 GND 0.17fF
C370 VDD.n19 GND 0.00fF
C371 VDD.n20 GND 0.00fF
C372 VDD.t11 GND 0.05fF $ **FLOATING
C373 VDD.n21 GND 0.01fF
C374 VDD.n22 GND 0.00fF
C375 VDD.t10 GND 0.11fF $ **FLOATING
C376 VDD.n24 GND 0.04fF
C377 VDD.n25 GND 0.00fF
C378 VDD.n26 GND 0.00fF
C379 VDD.n27 GND 0.00fF
C380 VDD.n28 GND 0.00fF
C381 VDD.n29 GND 0.01fF
C382 VDD.n30 GND 0.00fF
C383 VDD.n31 GND 0.00fF
C384 VDD.n32 GND 0.00fF
C385 VDD.n33 GND 0.00fF
C386 VDD.n34 GND 0.00fF
C387 VDD.n35 GND 0.03fF
C388 VDD.n36 GND 0.00fF
C389 VDD.n37 GND 0.17fF
C390 VDD.n38 GND 0.00fF
C391 VDD.n39 GND 0.00fF
C392 VDD.t7 GND 0.05fF $ **FLOATING
C393 VDD.n40 GND 0.01fF
C394 VDD.n41 GND 0.00fF
C395 VDD.t6 GND 0.11fF $ **FLOATING
C396 VDD.n43 GND 0.04fF
C397 VDD.n44 GND 0.00fF
C398 VDD.n45 GND 0.00fF
C399 VDD.n46 GND 0.00fF
C400 VDD.n47 GND 0.00fF
C401 VDD.n48 GND 0.01fF
C402 VDD.n49 GND 0.00fF
C403 VDD.n50 GND 0.00fF
C404 VDD.n51 GND 0.00fF
C405 VDD.n52 GND 0.00fF
C406 VDD.n53 GND 0.00fF
C407 VDD.n54 GND 0.03fF
C408 VDD.n55 GND 0.00fF
C409 VDD.n56 GND 0.17fF
C410 VDD.n57 GND 0.00fF
C411 VDD.n58 GND 0.00fF
C412 VDD.t1 GND 0.05fF $ **FLOATING
C413 VDD.n59 GND 0.01fF
C414 VDD.n60 GND 0.00fF
C415 VDD.t0 GND 0.11fF $ **FLOATING
C416 VDD.n62 GND 0.04fF
C417 VDD.n63 GND 0.00fF
C418 VDD.n64 GND 0.00fF
C419 VDD.n65 GND 0.00fF
C420 VDD.n66 GND 0.00fF
C421 VDD.n67 GND 0.01fF
C422 VDD.n68 GND 0.00fF
C423 VDD.n69 GND 0.00fF
C424 VDD.n70 GND 0.00fF
C425 VDD.n71 GND 0.00fF
C426 VDD.n72 GND 0.00fF
C427 VDD.n73 GND 0.03fF
C428 VDD.n74 GND 0.00fF
C429 VDD.n75 GND 0.17fF
C430 VDD.n76 GND 0.00fF
C431 VDD.n77 GND 0.00fF
C432 VDD.t5 GND 0.05fF $ **FLOATING
C433 VDD.n78 GND 0.01fF
C434 VDD.n79 GND 0.00fF
C435 VDD.t4 GND 0.11fF $ **FLOATING
C436 VDD.n81 GND 0.04fF
C437 VDD.n82 GND 0.00fF
C438 VDD.n83 GND 0.00fF
C439 VDD.n84 GND 0.00fF
C440 VDD.n85 GND 0.00fF
C441 VDD.n86 GND 0.01fF
C442 VDD.n87 GND 0.00fF
C443 VDD.n88 GND 0.00fF
C444 VDD.n89 GND 0.00fF
C445 VDD.n90 GND 0.00fF
C446 VDD.n91 GND 0.00fF
C447 VDD.n92 GND 0.03fF
C448 VDD.n93 GND 0.00fF
C449 VDD.n94 GND 0.17fF
C450 VDD.n95 GND 0.00fF
C451 VDD.n96 GND 0.00fF
C452 VDD.t3 GND 0.05fF $ **FLOATING
C453 VDD.n97 GND 0.01fF
C454 VDD.n98 GND 0.00fF
C455 VDD.t2 GND 0.11fF $ **FLOATING
C456 VDD.n100 GND 0.04fF
C457 VDD.n101 GND 0.00fF
C458 VDD.n102 GND 0.00fF
C459 VDD.n103 GND 0.00fF
C460 VDD.n104 GND 0.00fF
C461 VDD.n105 GND 0.01fF
C462 VDD.n106 GND 0.00fF
C463 VDD.n107 GND 0.00fF
C464 VDD.n108 GND 0.00fF
C465 VDD.n109 GND 0.00fF
C466 VDD.n110 GND 0.00fF
C467 VDD.n111 GND 0.03fF
C468 VDD.n112 GND 0.00fF
C469 VDD.n113 GND 11.56fF
C470 VDD.n114 GND 67.08fF
C471 VDD.n115 GND 20.84fF
C472 VDD.n116 GND 13.94fF
C473 VDD.n117 GND 13.94fF
C474 VDD.n118 GND 17.70fF
C475 bit0.n0 GND 0.00fF
C476 bit0.n1 GND 0.00fF
C477 bit0.t3 GND 0.02fF $ **FLOATING
C478 bit0.n2 GND 0.01fF
C479 bit0.n3 GND 0.00fF
C480 bit0.t1 GND 0.02fF $ **FLOATING
C481 bit0.n4 GND 0.01fF
C482 bit0.n5 GND 0.00fF
C483 bit0.n6 GND 0.06fF
C484 bit0.t0 GND 0.01fF $ **FLOATING
C485 bit0.t2 GND 0.01fF $ **FLOATING
C486 bit0.n7 GND 0.02fF
C487 bit0.n8 GND 77.65fF
C488 a_22576_75126.n0 GND 0.01fF
C489 a_22576_75126.n1 GND 0.01fF
C490 a_22576_75126.n2 GND 0.00fF
C491 a_22576_75126.n3 GND 0.00fF
C492 a_22576_75126.n4 GND 0.00fF
C493 a_22576_75126.n5 GND 0.00fF
C494 a_22576_75126.n6 GND 0.00fF
C495 a_22576_75126.n7 GND 0.00fF
C496 a_22576_75126.n8 GND 0.00fF
C497 a_22576_75126.n9 GND 0.00fF
C498 a_22576_75126.t1 GND 0.02fF $ **FLOATING
C499 a_22576_75126.t2 GND 0.02fF $ **FLOATING
C500 a_22576_75126.n10 GND 0.05fF
C501 a_22576_75126.n11 GND 0.00fF
C502 a_22576_75126.n12 GND 0.00fF
C503 a_22576_75126.n13 GND 0.02fF
C504 a_22576_75126.n14 GND 0.04fF
C505 a_22576_75126.n15 GND 0.12fF
C506 a_22576_75126.n16 GND 0.01fF
C507 a_22576_75126.n17 GND 0.12fF
C508 a_22576_75126.t3 GND 3.87fF $ **FLOATING
C509 a_22576_75126.n18 GND 0.52fF
C510 a_22576_75126.t0 GND 0.24fF $ **FLOATING
C511 a_22866_75202.n0 GND 0.00fF
C512 a_22866_75202.n1 GND 0.00fF
C513 a_22866_75202.n2 GND 0.01fF
C514 a_22866_75202.n3 GND 0.01fF
C515 a_22866_75202.n4 GND 0.00fF
C516 a_22866_75202.n5 GND 0.00fF
C517 a_22866_75202.n6 GND 0.00fF
C518 a_22866_75202.n7 GND 0.00fF
C519 a_22866_75202.n8 GND 0.00fF
C520 a_22866_75202.n9 GND 0.00fF
C521 a_22866_75202.n10 GND 0.09fF
C522 a_22866_75202.n11 GND 0.00fF
C523 a_22866_75202.n12 GND 0.01fF
C524 a_22866_75202.n13 GND 0.01fF
C525 a_22866_75202.n14 GND 0.01fF
C526 a_22866_75202.n15 GND 0.00fF
C527 a_22866_75202.n16 GND 0.00fF
C528 a_22866_75202.n17 GND 0.00fF
C529 a_22866_75202.t1 GND 0.02fF $ **FLOATING
C530 a_22866_75202.n18 GND 0.07fF
C531 a_22866_75202.n19 GND 0.02fF
C532 a_22866_75202.n20 GND 0.05fF
C533 a_22866_75202.n22 GND 0.04fF
C534 a_22866_75202.n23 GND 0.04fF
C535 a_22866_75202.n24 GND 0.00fF
C536 a_22866_75202.n25 GND 0.00fF
C537 a_22866_75202.t0 GND 0.02fF $ **FLOATING
C538 a_22866_75202.n26 GND 0.07fF
C539 a_22866_75202.n27 GND 0.02fF
C540 a_22866_75202.n28 GND 0.05fF
C541 a_22866_75202.n30 GND 0.01fF
C542 a_22866_75202.n31 GND 0.00fF
C543 a_22866_75202.n32 GND 0.00fF
C544 a_22866_75202.n33 GND 0.00fF
C545 a_22866_75202.n34 GND 0.00fF
C546 a_22866_75202.n35 GND 0.00fF
C547 a_22866_75202.n36 GND 0.00fF
C548 a_22866_75202.n38 GND 0.08fF
C549 a_22866_75202.t2 GND 4.19fF $ **FLOATING
C550 a_22866_75202.n39 GND 0.61fF
C551 a_22866_75202.t3 GND 0.26fF $ **FLOATING
C552 a_4466_25802.n0 GND 0.00fF
C553 a_4466_25802.n1 GND 0.00fF
C554 a_4466_25802.n2 GND 0.01fF
C555 a_4466_25802.n3 GND 0.01fF
C556 a_4466_25802.n4 GND 0.00fF
C557 a_4466_25802.n5 GND 0.00fF
C558 a_4466_25802.n6 GND 0.00fF
C559 a_4466_25802.n7 GND 0.00fF
C560 a_4466_25802.n8 GND 0.00fF
C561 a_4466_25802.n9 GND 0.00fF
C562 a_4466_25802.n10 GND 0.09fF
C563 a_4466_25802.n11 GND 0.00fF
C564 a_4466_25802.n12 GND 0.01fF
C565 a_4466_25802.n13 GND 0.01fF
C566 a_4466_25802.n14 GND 0.01fF
C567 a_4466_25802.n15 GND 0.00fF
C568 a_4466_25802.n16 GND 0.00fF
C569 a_4466_25802.n17 GND 0.00fF
C570 a_4466_25802.t0 GND 0.02fF $ **FLOATING
C571 a_4466_25802.n18 GND 0.07fF
C572 a_4466_25802.n19 GND 0.02fF
C573 a_4466_25802.n20 GND 0.05fF
C574 a_4466_25802.n22 GND 0.04fF
C575 a_4466_25802.n23 GND 0.04fF
C576 a_4466_25802.n24 GND 0.00fF
C577 a_4466_25802.n25 GND 0.00fF
C578 a_4466_25802.t1 GND 0.02fF $ **FLOATING
C579 a_4466_25802.n26 GND 0.07fF
C580 a_4466_25802.n27 GND 0.02fF
C581 a_4466_25802.n28 GND 0.05fF
C582 a_4466_25802.n30 GND 0.01fF
C583 a_4466_25802.n31 GND 0.00fF
C584 a_4466_25802.n32 GND 0.00fF
C585 a_4466_25802.n33 GND 0.00fF
C586 a_4466_25802.n34 GND 0.00fF
C587 a_4466_25802.n35 GND 0.00fF
C588 a_4466_25802.n36 GND 0.00fF
C589 a_4466_25802.n38 GND 0.08fF
C590 a_4466_25802.t3 GND 4.19fF $ **FLOATING
C591 a_4466_25802.n39 GND 0.61fF
C592 a_4466_25802.t2 GND 0.26fF $ **FLOATING
C593 a_13666_45562.n0 GND 0.00fF
C594 a_13666_45562.n1 GND 0.00fF
C595 a_13666_45562.n2 GND 0.01fF
C596 a_13666_45562.n3 GND 0.01fF
C597 a_13666_45562.n4 GND 0.00fF
C598 a_13666_45562.n5 GND 0.00fF
C599 a_13666_45562.n6 GND 0.00fF
C600 a_13666_45562.n7 GND 0.00fF
C601 a_13666_45562.n8 GND 0.00fF
C602 a_13666_45562.n9 GND 0.00fF
C603 a_13666_45562.n10 GND 0.09fF
C604 a_13666_45562.n11 GND 0.00fF
C605 a_13666_45562.n12 GND 0.01fF
C606 a_13666_45562.n13 GND 0.01fF
C607 a_13666_45562.n14 GND 0.01fF
C608 a_13666_45562.n15 GND 0.00fF
C609 a_13666_45562.n16 GND 0.00fF
C610 a_13666_45562.n17 GND 0.00fF
C611 a_13666_45562.t0 GND 0.02fF $ **FLOATING
C612 a_13666_45562.n18 GND 0.07fF
C613 a_13666_45562.n19 GND 0.02fF
C614 a_13666_45562.n20 GND 0.05fF
C615 a_13666_45562.n22 GND 0.04fF
C616 a_13666_45562.n23 GND 0.04fF
C617 a_13666_45562.n24 GND 0.00fF
C618 a_13666_45562.n25 GND 0.00fF
C619 a_13666_45562.t1 GND 0.02fF $ **FLOATING
C620 a_13666_45562.n26 GND 0.07fF
C621 a_13666_45562.n27 GND 0.02fF
C622 a_13666_45562.n28 GND 0.05fF
C623 a_13666_45562.n30 GND 0.01fF
C624 a_13666_45562.n31 GND 0.00fF
C625 a_13666_45562.n32 GND 0.00fF
C626 a_13666_45562.n33 GND 0.00fF
C627 a_13666_45562.n34 GND 0.00fF
C628 a_13666_45562.n35 GND 0.00fF
C629 a_13666_45562.n36 GND 0.00fF
C630 a_13666_45562.n38 GND 0.08fF
C631 a_13666_45562.t2 GND 4.19fF $ **FLOATING
C632 a_13666_45562.n39 GND 0.61fF
C633 a_13666_45562.t3 GND 0.26fF $ **FLOATING
C634 a_22866_35682.n0 GND 0.00fF
C635 a_22866_35682.n1 GND 0.00fF
C636 a_22866_35682.n2 GND 0.01fF
C637 a_22866_35682.n3 GND 0.01fF
C638 a_22866_35682.n4 GND 0.00fF
C639 a_22866_35682.n5 GND 0.00fF
C640 a_22866_35682.n6 GND 0.00fF
C641 a_22866_35682.n7 GND 0.00fF
C642 a_22866_35682.n8 GND 0.00fF
C643 a_22866_35682.n9 GND 0.00fF
C644 a_22866_35682.n10 GND 0.09fF
C645 a_22866_35682.n11 GND 0.00fF
C646 a_22866_35682.n12 GND 0.01fF
C647 a_22866_35682.n13 GND 0.01fF
C648 a_22866_35682.n14 GND 0.01fF
C649 a_22866_35682.n15 GND 0.00fF
C650 a_22866_35682.n16 GND 0.00fF
C651 a_22866_35682.n17 GND 0.00fF
C652 a_22866_35682.t0 GND 0.02fF $ **FLOATING
C653 a_22866_35682.n18 GND 0.07fF
C654 a_22866_35682.n19 GND 0.02fF
C655 a_22866_35682.n20 GND 0.05fF
C656 a_22866_35682.n22 GND 0.04fF
C657 a_22866_35682.n23 GND 0.04fF
C658 a_22866_35682.n24 GND 0.00fF
C659 a_22866_35682.n25 GND 0.00fF
C660 a_22866_35682.t1 GND 0.02fF $ **FLOATING
C661 a_22866_35682.n26 GND 0.07fF
C662 a_22866_35682.n27 GND 0.02fF
C663 a_22866_35682.n28 GND 0.05fF
C664 a_22866_35682.n30 GND 0.01fF
C665 a_22866_35682.n31 GND 0.00fF
C666 a_22866_35682.n32 GND 0.00fF
C667 a_22866_35682.n33 GND 0.00fF
C668 a_22866_35682.n34 GND 0.00fF
C669 a_22866_35682.n35 GND 0.00fF
C670 a_22866_35682.n36 GND 0.00fF
C671 a_22866_35682.n38 GND 0.08fF
C672 a_22866_35682.t2 GND 4.19fF $ **FLOATING
C673 a_22866_35682.n39 GND 0.61fF
C674 a_22866_35682.t3 GND 0.26fF $ **FLOATING
C675 a_68866_55442.n0 GND 0.00fF
C676 a_68866_55442.n1 GND 0.00fF
C677 a_68866_55442.n2 GND 0.01fF
C678 a_68866_55442.n3 GND 0.01fF
C679 a_68866_55442.n4 GND 0.00fF
C680 a_68866_55442.n5 GND 0.00fF
C681 a_68866_55442.n6 GND 0.00fF
C682 a_68866_55442.n7 GND 0.00fF
C683 a_68866_55442.n8 GND 0.00fF
C684 a_68866_55442.n9 GND 0.00fF
C685 a_68866_55442.n10 GND 0.09fF
C686 a_68866_55442.n11 GND 0.00fF
C687 a_68866_55442.n12 GND 0.01fF
C688 a_68866_55442.n13 GND 0.01fF
C689 a_68866_55442.n14 GND 0.01fF
C690 a_68866_55442.n15 GND 0.00fF
C691 a_68866_55442.n16 GND 0.00fF
C692 a_68866_55442.n17 GND 0.00fF
C693 a_68866_55442.t1 GND 0.02fF $ **FLOATING
C694 a_68866_55442.n18 GND 0.07fF
C695 a_68866_55442.n19 GND 0.02fF
C696 a_68866_55442.n20 GND 0.05fF
C697 a_68866_55442.n22 GND 0.04fF
C698 a_68866_55442.n23 GND 0.04fF
C699 a_68866_55442.n24 GND 0.00fF
C700 a_68866_55442.n25 GND 0.00fF
C701 a_68866_55442.t2 GND 0.02fF $ **FLOATING
C702 a_68866_55442.n26 GND 0.07fF
C703 a_68866_55442.n27 GND 0.02fF
C704 a_68866_55442.n28 GND 0.05fF
C705 a_68866_55442.n30 GND 0.01fF
C706 a_68866_55442.n31 GND 0.00fF
C707 a_68866_55442.n32 GND 0.00fF
C708 a_68866_55442.n33 GND 0.00fF
C709 a_68866_55442.n34 GND 0.00fF
C710 a_68866_55442.n35 GND 0.00fF
C711 a_68866_55442.n36 GND 0.00fF
C712 a_68866_55442.n38 GND 0.08fF
C713 a_68866_55442.t3 GND 4.19fF $ **FLOATING
C714 a_68866_55442.n39 GND 0.61fF
C715 a_68866_55442.t0 GND 0.26fF $ **FLOATING
C716 a_13376_75126.n0 GND 0.01fF
C717 a_13376_75126.n1 GND 0.01fF
C718 a_13376_75126.n2 GND 0.00fF
C719 a_13376_75126.n3 GND 0.00fF
C720 a_13376_75126.n4 GND 0.00fF
C721 a_13376_75126.n5 GND 0.00fF
C722 a_13376_75126.n6 GND 0.00fF
C723 a_13376_75126.n7 GND 0.00fF
C724 a_13376_75126.n8 GND 0.00fF
C725 a_13376_75126.n9 GND 0.00fF
C726 a_13376_75126.t0 GND 0.02fF $ **FLOATING
C727 a_13376_75126.t1 GND 0.02fF $ **FLOATING
C728 a_13376_75126.n10 GND 0.05fF
C729 a_13376_75126.n11 GND 0.00fF
C730 a_13376_75126.n12 GND 0.00fF
C731 a_13376_75126.n13 GND 0.02fF
C732 a_13376_75126.n14 GND 0.04fF
C733 a_13376_75126.n15 GND 0.12fF
C734 a_13376_75126.n16 GND 0.01fF
C735 a_13376_75126.n17 GND 0.12fF
C736 a_13376_75126.t2 GND 3.87fF $ **FLOATING
C737 a_13376_75126.n18 GND 0.52fF
C738 a_13376_75126.t3 GND 0.24fF $ **FLOATING
C739 a_13666_75202.n0 GND 0.00fF
C740 a_13666_75202.n1 GND 0.00fF
C741 a_13666_75202.n2 GND 0.01fF
C742 a_13666_75202.n3 GND 0.01fF
C743 a_13666_75202.n4 GND 0.00fF
C744 a_13666_75202.n5 GND 0.00fF
C745 a_13666_75202.n6 GND 0.00fF
C746 a_13666_75202.n7 GND 0.00fF
C747 a_13666_75202.n8 GND 0.00fF
C748 a_13666_75202.n9 GND 0.00fF
C749 a_13666_75202.n10 GND 0.09fF
C750 a_13666_75202.n11 GND 0.00fF
C751 a_13666_75202.n12 GND 0.01fF
C752 a_13666_75202.n13 GND 0.01fF
C753 a_13666_75202.n14 GND 0.01fF
C754 a_13666_75202.n15 GND 0.00fF
C755 a_13666_75202.n16 GND 0.00fF
C756 a_13666_75202.n17 GND 0.00fF
C757 a_13666_75202.t2 GND 0.02fF $ **FLOATING
C758 a_13666_75202.n18 GND 0.07fF
C759 a_13666_75202.n19 GND 0.02fF
C760 a_13666_75202.n20 GND 0.05fF
C761 a_13666_75202.n22 GND 0.04fF
C762 a_13666_75202.n23 GND 0.04fF
C763 a_13666_75202.n24 GND 0.00fF
C764 a_13666_75202.n25 GND 0.00fF
C765 a_13666_75202.t1 GND 0.02fF $ **FLOATING
C766 a_13666_75202.n26 GND 0.07fF
C767 a_13666_75202.n27 GND 0.02fF
C768 a_13666_75202.n28 GND 0.05fF
C769 a_13666_75202.n30 GND 0.01fF
C770 a_13666_75202.n31 GND 0.00fF
C771 a_13666_75202.n32 GND 0.00fF
C772 a_13666_75202.n33 GND 0.00fF
C773 a_13666_75202.n34 GND 0.00fF
C774 a_13666_75202.n35 GND 0.00fF
C775 a_13666_75202.n36 GND 0.00fF
C776 a_13666_75202.n38 GND 0.08fF
C777 a_13666_75202.t3 GND 4.19fF $ **FLOATING
C778 a_13666_75202.n39 GND 0.61fF
C779 a_13666_75202.t0 GND 0.26fF $ **FLOATING
C780 a_41266_6042.n0 GND 0.00fF
C781 a_41266_6042.n1 GND 0.00fF
C782 a_41266_6042.n2 GND 0.01fF
C783 a_41266_6042.n3 GND 0.01fF
C784 a_41266_6042.n4 GND 0.00fF
C785 a_41266_6042.n5 GND 0.00fF
C786 a_41266_6042.n6 GND 0.00fF
C787 a_41266_6042.n7 GND 0.00fF
C788 a_41266_6042.n8 GND 0.00fF
C789 a_41266_6042.n9 GND 0.00fF
C790 a_41266_6042.n10 GND 0.09fF
C791 a_41266_6042.n11 GND 0.00fF
C792 a_41266_6042.n12 GND 0.01fF
C793 a_41266_6042.n13 GND 0.01fF
C794 a_41266_6042.n14 GND 0.01fF
C795 a_41266_6042.n15 GND 0.00fF
C796 a_41266_6042.n16 GND 0.00fF
C797 a_41266_6042.n17 GND 0.00fF
C798 a_41266_6042.t1 GND 0.02fF $ **FLOATING
C799 a_41266_6042.n18 GND 0.07fF
C800 a_41266_6042.n19 GND 0.02fF
C801 a_41266_6042.n20 GND 0.05fF
C802 a_41266_6042.n22 GND 0.04fF
C803 a_41266_6042.n23 GND 0.04fF
C804 a_41266_6042.n24 GND 0.00fF
C805 a_41266_6042.n25 GND 0.00fF
C806 a_41266_6042.t2 GND 0.02fF $ **FLOATING
C807 a_41266_6042.n26 GND 0.07fF
C808 a_41266_6042.n27 GND 0.02fF
C809 a_41266_6042.n28 GND 0.05fF
C810 a_41266_6042.n30 GND 0.01fF
C811 a_41266_6042.n31 GND 0.00fF
C812 a_41266_6042.n32 GND 0.00fF
C813 a_41266_6042.n33 GND 0.00fF
C814 a_41266_6042.n34 GND 0.00fF
C815 a_41266_6042.n35 GND 0.00fF
C816 a_41266_6042.n36 GND 0.00fF
C817 a_41266_6042.n38 GND 0.08fF
C818 a_41266_6042.t3 GND 4.19fF $ **FLOATING
C819 a_41266_6042.n39 GND 0.61fF
C820 a_41266_6042.t0 GND 0.26fF $ **FLOATING
C821 a_13666_35682.n0 GND 0.00fF
C822 a_13666_35682.n1 GND 0.00fF
C823 a_13666_35682.n2 GND 0.01fF
C824 a_13666_35682.n3 GND 0.01fF
C825 a_13666_35682.n4 GND 0.00fF
C826 a_13666_35682.n5 GND 0.00fF
C827 a_13666_35682.n6 GND 0.00fF
C828 a_13666_35682.n7 GND 0.00fF
C829 a_13666_35682.n8 GND 0.00fF
C830 a_13666_35682.n9 GND 0.00fF
C831 a_13666_35682.n10 GND 0.09fF
C832 a_13666_35682.n11 GND 0.00fF
C833 a_13666_35682.n12 GND 0.01fF
C834 a_13666_35682.n13 GND 0.01fF
C835 a_13666_35682.n14 GND 0.01fF
C836 a_13666_35682.n15 GND 0.00fF
C837 a_13666_35682.n16 GND 0.00fF
C838 a_13666_35682.n17 GND 0.00fF
C839 a_13666_35682.t0 GND 0.02fF $ **FLOATING
C840 a_13666_35682.n18 GND 0.07fF
C841 a_13666_35682.n19 GND 0.02fF
C842 a_13666_35682.n20 GND 0.05fF
C843 a_13666_35682.n22 GND 0.04fF
C844 a_13666_35682.n23 GND 0.04fF
C845 a_13666_35682.n24 GND 0.00fF
C846 a_13666_35682.n25 GND 0.00fF
C847 a_13666_35682.t1 GND 0.02fF $ **FLOATING
C848 a_13666_35682.n26 GND 0.07fF
C849 a_13666_35682.n27 GND 0.02fF
C850 a_13666_35682.n28 GND 0.05fF
C851 a_13666_35682.n30 GND 0.01fF
C852 a_13666_35682.n31 GND 0.00fF
C853 a_13666_35682.n32 GND 0.00fF
C854 a_13666_35682.n33 GND 0.00fF
C855 a_13666_35682.n34 GND 0.00fF
C856 a_13666_35682.n35 GND 0.00fF
C857 a_13666_35682.n36 GND 0.00fF
C858 a_13666_35682.n38 GND 0.08fF
C859 a_13666_35682.t2 GND 4.19fF $ **FLOATING
C860 a_13666_35682.n39 GND 0.61fF
C861 a_13666_35682.t3 GND 0.26fF $ **FLOATING
C862 a_40976_5966.n0 GND 0.01fF
C863 a_40976_5966.n1 GND 0.01fF
C864 a_40976_5966.n2 GND 0.00fF
C865 a_40976_5966.n3 GND 0.00fF
C866 a_40976_5966.n4 GND 0.00fF
C867 a_40976_5966.n5 GND 0.00fF
C868 a_40976_5966.n6 GND 0.00fF
C869 a_40976_5966.n7 GND 0.00fF
C870 a_40976_5966.n8 GND 0.00fF
C871 a_40976_5966.n9 GND 0.00fF
C872 a_40976_5966.t1 GND 0.02fF $ **FLOATING
C873 a_40976_5966.t0 GND 0.02fF $ **FLOATING
C874 a_40976_5966.n10 GND 0.05fF
C875 a_40976_5966.n11 GND 0.00fF
C876 a_40976_5966.n12 GND 0.00fF
C877 a_40976_5966.n13 GND 0.02fF
C878 a_40976_5966.n14 GND 0.04fF
C879 a_40976_5966.n15 GND 0.12fF
C880 a_40976_5966.n16 GND 0.01fF
C881 a_40976_5966.n17 GND 0.12fF
C882 a_40976_5966.t2 GND 3.87fF $ **FLOATING
C883 a_40976_5966.n18 GND 0.52fF
C884 a_40976_5966.t3 GND 0.24fF $ **FLOATING
C885 a_n436_84486.t2 GND 0.04fF $ **FLOATING
C886 a_n436_84486.t1 GND 0.07fF $ **FLOATING
C887 a_n436_84486.t4 GND 0.07fF $ **FLOATING
C888 a_n436_84486.t0 GND 0.07fF $ **FLOATING
C889 a_n436_84486.t5 GND 0.12fF $ **FLOATING
C890 a_n436_84486.n0 GND 21.77fF
C891 a_n436_84486.n1 GND 10.89fF
C892 a_n436_84486.n2 GND 12.33fF
C893 a_n436_84486.n3 GND 0.06fF
C894 a_n436_84486.t3 GND 0.09fF $ **FLOATING
C895 a_68576_25726.n0 GND 0.01fF
C896 a_68576_25726.n1 GND 0.01fF
C897 a_68576_25726.n2 GND 0.00fF
C898 a_68576_25726.n3 GND 0.00fF
C899 a_68576_25726.n4 GND 0.00fF
C900 a_68576_25726.n5 GND 0.00fF
C901 a_68576_25726.n6 GND 0.00fF
C902 a_68576_25726.n7 GND 0.00fF
C903 a_68576_25726.n8 GND 0.00fF
C904 a_68576_25726.n9 GND 0.00fF
C905 a_68576_25726.t1 GND 0.02fF $ **FLOATING
C906 a_68576_25726.t2 GND 0.02fF $ **FLOATING
C907 a_68576_25726.n10 GND 0.05fF
C908 a_68576_25726.n11 GND 0.00fF
C909 a_68576_25726.n12 GND 0.00fF
C910 a_68576_25726.n13 GND 0.02fF
C911 a_68576_25726.n14 GND 0.04fF
C912 a_68576_25726.n15 GND 0.12fF
C913 a_68576_25726.n16 GND 0.01fF
C914 a_68576_25726.n17 GND 0.12fF
C915 a_68576_25726.t3 GND 3.87fF $ **FLOATING
C916 a_68576_25726.n18 GND 0.52fF
C917 a_68576_25726.t0 GND 0.24fF $ **FLOATING
C918 a_68866_25802.n0 GND 0.00fF
C919 a_68866_25802.n1 GND 0.00fF
C920 a_68866_25802.n2 GND 0.01fF
C921 a_68866_25802.n3 GND 0.01fF
C922 a_68866_25802.n4 GND 0.00fF
C923 a_68866_25802.n5 GND 0.00fF
C924 a_68866_25802.n6 GND 0.00fF
C925 a_68866_25802.n7 GND 0.00fF
C926 a_68866_25802.n8 GND 0.00fF
C927 a_68866_25802.n9 GND 0.00fF
C928 a_68866_25802.n10 GND 0.09fF
C929 a_68866_25802.n11 GND 0.00fF
C930 a_68866_25802.n12 GND 0.01fF
C931 a_68866_25802.n13 GND 0.01fF
C932 a_68866_25802.n14 GND 0.01fF
C933 a_68866_25802.n15 GND 0.00fF
C934 a_68866_25802.n16 GND 0.00fF
C935 a_68866_25802.n17 GND 0.00fF
C936 a_68866_25802.t2 GND 0.02fF $ **FLOATING
C937 a_68866_25802.n18 GND 0.07fF
C938 a_68866_25802.n19 GND 0.02fF
C939 a_68866_25802.n20 GND 0.05fF
C940 a_68866_25802.n22 GND 0.04fF
C941 a_68866_25802.n23 GND 0.04fF
C942 a_68866_25802.n24 GND 0.00fF
C943 a_68866_25802.n25 GND 0.00fF
C944 a_68866_25802.t1 GND 0.02fF $ **FLOATING
C945 a_68866_25802.n26 GND 0.07fF
C946 a_68866_25802.n27 GND 0.02fF
C947 a_68866_25802.n28 GND 0.05fF
C948 a_68866_25802.n30 GND 0.01fF
C949 a_68866_25802.n31 GND 0.00fF
C950 a_68866_25802.n32 GND 0.00fF
C951 a_68866_25802.n33 GND 0.00fF
C952 a_68866_25802.n34 GND 0.00fF
C953 a_68866_25802.n35 GND 0.00fF
C954 a_68866_25802.n36 GND 0.00fF
C955 a_68866_25802.n38 GND 0.08fF
C956 a_68866_25802.t3 GND 4.19fF $ **FLOATING
C957 a_68866_25802.n39 GND 0.61fF
C958 a_68866_25802.t0 GND 0.26fF $ **FLOATING
C959 a_59666_45562.n0 GND 0.00fF
C960 a_59666_45562.n1 GND 0.00fF
C961 a_59666_45562.n2 GND 0.01fF
C962 a_59666_45562.n3 GND 0.01fF
C963 a_59666_45562.n4 GND 0.00fF
C964 a_59666_45562.n5 GND 0.00fF
C965 a_59666_45562.n6 GND 0.00fF
C966 a_59666_45562.n7 GND 0.00fF
C967 a_59666_45562.n8 GND 0.00fF
C968 a_59666_45562.n9 GND 0.00fF
C969 a_59666_45562.n10 GND 0.09fF
C970 a_59666_45562.n11 GND 0.00fF
C971 a_59666_45562.n12 GND 0.01fF
C972 a_59666_45562.n13 GND 0.01fF
C973 a_59666_45562.n14 GND 0.01fF
C974 a_59666_45562.n15 GND 0.00fF
C975 a_59666_45562.n16 GND 0.00fF
C976 a_59666_45562.n17 GND 0.00fF
C977 a_59666_45562.t0 GND 0.02fF $ **FLOATING
C978 a_59666_45562.n18 GND 0.07fF
C979 a_59666_45562.n19 GND 0.02fF
C980 a_59666_45562.n20 GND 0.05fF
C981 a_59666_45562.n22 GND 0.04fF
C982 a_59666_45562.n23 GND 0.04fF
C983 a_59666_45562.n24 GND 0.00fF
C984 a_59666_45562.n25 GND 0.00fF
C985 a_59666_45562.t1 GND 0.02fF $ **FLOATING
C986 a_59666_45562.n26 GND 0.07fF
C987 a_59666_45562.n27 GND 0.02fF
C988 a_59666_45562.n28 GND 0.05fF
C989 a_59666_45562.n30 GND 0.01fF
C990 a_59666_45562.n31 GND 0.00fF
C991 a_59666_45562.n32 GND 0.00fF
C992 a_59666_45562.n33 GND 0.00fF
C993 a_59666_45562.n34 GND 0.00fF
C994 a_59666_45562.n35 GND 0.00fF
C995 a_59666_45562.n36 GND 0.00fF
C996 a_59666_45562.n38 GND 0.08fF
C997 a_59666_45562.t3 GND 4.19fF $ **FLOATING
C998 a_59666_45562.n39 GND 0.61fF
C999 a_59666_45562.t2 GND 0.26fF $ **FLOATING
C1000 a_32066_75202.n0 GND 0.00fF
C1001 a_32066_75202.n1 GND 0.00fF
C1002 a_32066_75202.n2 GND 0.01fF
C1003 a_32066_75202.n3 GND 0.01fF
C1004 a_32066_75202.n4 GND 0.00fF
C1005 a_32066_75202.n5 GND 0.00fF
C1006 a_32066_75202.n6 GND 0.00fF
C1007 a_32066_75202.n7 GND 0.00fF
C1008 a_32066_75202.n8 GND 0.00fF
C1009 a_32066_75202.n9 GND 0.00fF
C1010 a_32066_75202.n10 GND 0.09fF
C1011 a_32066_75202.n11 GND 0.00fF
C1012 a_32066_75202.n12 GND 0.01fF
C1013 a_32066_75202.n13 GND 0.01fF
C1014 a_32066_75202.n14 GND 0.01fF
C1015 a_32066_75202.n15 GND 0.00fF
C1016 a_32066_75202.n16 GND 0.00fF
C1017 a_32066_75202.n17 GND 0.00fF
C1018 a_32066_75202.t1 GND 0.02fF $ **FLOATING
C1019 a_32066_75202.n18 GND 0.07fF
C1020 a_32066_75202.n19 GND 0.02fF
C1021 a_32066_75202.n20 GND 0.05fF
C1022 a_32066_75202.n22 GND 0.04fF
C1023 a_32066_75202.n23 GND 0.04fF
C1024 a_32066_75202.n24 GND 0.00fF
C1025 a_32066_75202.n25 GND 0.00fF
C1026 a_32066_75202.t0 GND 0.02fF $ **FLOATING
C1027 a_32066_75202.n26 GND 0.07fF
C1028 a_32066_75202.n27 GND 0.02fF
C1029 a_32066_75202.n28 GND 0.05fF
C1030 a_32066_75202.n30 GND 0.01fF
C1031 a_32066_75202.n31 GND 0.00fF
C1032 a_32066_75202.n32 GND 0.00fF
C1033 a_32066_75202.n33 GND 0.00fF
C1034 a_32066_75202.n34 GND 0.00fF
C1035 a_32066_75202.n35 GND 0.00fF
C1036 a_32066_75202.n36 GND 0.00fF
C1037 a_32066_75202.n38 GND 0.08fF
C1038 a_32066_75202.t2 GND 4.19fF $ **FLOATING
C1039 a_32066_75202.n39 GND 0.61fF
C1040 a_32066_75202.t3 GND 0.26fF $ **FLOATING
C1041 a_50176_65246.n0 GND 0.01fF
C1042 a_50176_65246.n1 GND 0.01fF
C1043 a_50176_65246.n2 GND 0.00fF
C1044 a_50176_65246.n3 GND 0.00fF
C1045 a_50176_65246.n4 GND 0.00fF
C1046 a_50176_65246.n5 GND 0.00fF
C1047 a_50176_65246.n6 GND 0.00fF
C1048 a_50176_65246.n7 GND 0.00fF
C1049 a_50176_65246.n8 GND 0.00fF
C1050 a_50176_65246.n9 GND 0.00fF
C1051 a_50176_65246.t0 GND 0.02fF $ **FLOATING
C1052 a_50176_65246.t1 GND 0.02fF $ **FLOATING
C1053 a_50176_65246.n10 GND 0.05fF
C1054 a_50176_65246.n11 GND 0.00fF
C1055 a_50176_65246.n12 GND 0.00fF
C1056 a_50176_65246.n13 GND 0.02fF
C1057 a_50176_65246.n14 GND 0.04fF
C1058 a_50176_65246.n15 GND 0.12fF
C1059 a_50176_65246.n16 GND 0.01fF
C1060 a_50176_65246.n17 GND 0.12fF
C1061 a_50176_65246.t2 GND 3.87fF $ **FLOATING
C1062 a_50176_65246.n18 GND 0.52fF
C1063 a_50176_65246.t3 GND 0.24fF $ **FLOATING
C1064 a_31776_75126.n0 GND 0.01fF
C1065 a_31776_75126.n1 GND 0.01fF
C1066 a_31776_75126.n2 GND 0.00fF
C1067 a_31776_75126.n3 GND 0.00fF
C1068 a_31776_75126.n4 GND 0.00fF
C1069 a_31776_75126.n5 GND 0.00fF
C1070 a_31776_75126.n6 GND 0.00fF
C1071 a_31776_75126.n7 GND 0.00fF
C1072 a_31776_75126.n8 GND 0.00fF
C1073 a_31776_75126.n9 GND 0.00fF
C1074 a_31776_75126.t1 GND 0.02fF $ **FLOATING
C1075 a_31776_75126.t2 GND 0.02fF $ **FLOATING
C1076 a_31776_75126.n10 GND 0.05fF
C1077 a_31776_75126.n11 GND 0.00fF
C1078 a_31776_75126.n12 GND 0.00fF
C1079 a_31776_75126.n13 GND 0.02fF
C1080 a_31776_75126.n14 GND 0.04fF
C1081 a_31776_75126.n15 GND 0.12fF
C1082 a_31776_75126.n16 GND 0.01fF
C1083 a_31776_75126.n17 GND 0.12fF
C1084 a_31776_75126.t3 GND 3.87fF $ **FLOATING
C1085 a_31776_75126.n18 GND 0.52fF
C1086 a_31776_75126.t0 GND 0.24fF $ **FLOATING
C1087 a_59376_5966.n0 GND 0.01fF
C1088 a_59376_5966.n1 GND 0.01fF
C1089 a_59376_5966.n2 GND 0.00fF
C1090 a_59376_5966.n3 GND 0.00fF
C1091 a_59376_5966.n4 GND 0.00fF
C1092 a_59376_5966.n5 GND 0.00fF
C1093 a_59376_5966.n6 GND 0.00fF
C1094 a_59376_5966.n7 GND 0.00fF
C1095 a_59376_5966.n8 GND 0.00fF
C1096 a_59376_5966.n9 GND 0.00fF
C1097 a_59376_5966.t1 GND 0.02fF $ **FLOATING
C1098 a_59376_5966.t0 GND 0.02fF $ **FLOATING
C1099 a_59376_5966.n10 GND 0.05fF
C1100 a_59376_5966.n11 GND 0.00fF
C1101 a_59376_5966.n12 GND 0.00fF
C1102 a_59376_5966.n13 GND 0.02fF
C1103 a_59376_5966.n14 GND 0.04fF
C1104 a_59376_5966.n15 GND 0.12fF
C1105 a_59376_5966.n16 GND 0.01fF
C1106 a_59376_5966.n17 GND 0.12fF
C1107 a_59376_5966.t2 GND 3.87fF $ **FLOATING
C1108 a_59376_5966.n18 GND 0.52fF
C1109 a_59376_5966.t3 GND 0.24fF $ **FLOATING
C1110 a_40976_45486.n0 GND 0.01fF
C1111 a_40976_45486.n1 GND 0.01fF
C1112 a_40976_45486.n2 GND 0.00fF
C1113 a_40976_45486.n3 GND 0.00fF
C1114 a_40976_45486.n4 GND 0.00fF
C1115 a_40976_45486.n5 GND 0.00fF
C1116 a_40976_45486.n6 GND 0.00fF
C1117 a_40976_45486.n7 GND 0.00fF
C1118 a_40976_45486.n8 GND 0.00fF
C1119 a_40976_45486.n9 GND 0.00fF
C1120 a_40976_45486.t1 GND 0.02fF $ **FLOATING
C1121 a_40976_45486.t0 GND 0.02fF $ **FLOATING
C1122 a_40976_45486.n10 GND 0.05fF
C1123 a_40976_45486.n11 GND 0.00fF
C1124 a_40976_45486.n12 GND 0.00fF
C1125 a_40976_45486.n13 GND 0.02fF
C1126 a_40976_45486.n14 GND 0.04fF
C1127 a_40976_45486.n15 GND 0.12fF
C1128 a_40976_45486.n16 GND 0.01fF
C1129 a_40976_45486.n17 GND 0.12fF
C1130 a_40976_45486.t2 GND 3.87fF $ **FLOATING
C1131 a_40976_45486.n18 GND 0.52fF
C1132 a_40976_45486.t3 GND 0.24fF $ **FLOATING
C1133 a_68866_65322.n0 GND 0.00fF
C1134 a_68866_65322.n1 GND 0.00fF
C1135 a_68866_65322.n2 GND 0.01fF
C1136 a_68866_65322.n3 GND 0.01fF
C1137 a_68866_65322.n4 GND 0.00fF
C1138 a_68866_65322.n5 GND 0.00fF
C1139 a_68866_65322.n6 GND 0.00fF
C1140 a_68866_65322.n7 GND 0.00fF
C1141 a_68866_65322.n8 GND 0.00fF
C1142 a_68866_65322.n9 GND 0.00fF
C1143 a_68866_65322.n10 GND 0.09fF
C1144 a_68866_65322.n11 GND 0.00fF
C1145 a_68866_65322.n12 GND 0.01fF
C1146 a_68866_65322.n13 GND 0.01fF
C1147 a_68866_65322.n14 GND 0.01fF
C1148 a_68866_65322.n15 GND 0.00fF
C1149 a_68866_65322.n16 GND 0.00fF
C1150 a_68866_65322.n17 GND 0.00fF
C1151 a_68866_65322.t0 GND 0.02fF $ **FLOATING
C1152 a_68866_65322.n18 GND 0.07fF
C1153 a_68866_65322.n19 GND 0.02fF
C1154 a_68866_65322.n20 GND 0.05fF
C1155 a_68866_65322.n22 GND 0.04fF
C1156 a_68866_65322.n23 GND 0.04fF
C1157 a_68866_65322.n24 GND 0.00fF
C1158 a_68866_65322.n25 GND 0.00fF
C1159 a_68866_65322.t1 GND 0.02fF $ **FLOATING
C1160 a_68866_65322.n26 GND 0.07fF
C1161 a_68866_65322.n27 GND 0.02fF
C1162 a_68866_65322.n28 GND 0.05fF
C1163 a_68866_65322.n30 GND 0.01fF
C1164 a_68866_65322.n31 GND 0.00fF
C1165 a_68866_65322.n32 GND 0.00fF
C1166 a_68866_65322.n33 GND 0.00fF
C1167 a_68866_65322.n34 GND 0.00fF
C1168 a_68866_65322.n35 GND 0.00fF
C1169 a_68866_65322.n36 GND 0.00fF
C1170 a_68866_65322.n38 GND 0.08fF
C1171 a_68866_65322.t3 GND 4.19fF $ **FLOATING
C1172 a_68866_65322.n39 GND 0.61fF
C1173 a_68866_65322.t2 GND 0.26fF $ **FLOATING
C1174 a_22576_65246.n0 GND 0.01fF
C1175 a_22576_65246.n1 GND 0.01fF
C1176 a_22576_65246.n2 GND 0.00fF
C1177 a_22576_65246.n3 GND 0.00fF
C1178 a_22576_65246.n4 GND 0.00fF
C1179 a_22576_65246.n5 GND 0.00fF
C1180 a_22576_65246.n6 GND 0.00fF
C1181 a_22576_65246.n7 GND 0.00fF
C1182 a_22576_65246.n8 GND 0.00fF
C1183 a_22576_65246.n9 GND 0.00fF
C1184 a_22576_65246.t0 GND 0.02fF $ **FLOATING
C1185 a_22576_65246.t1 GND 0.02fF $ **FLOATING
C1186 a_22576_65246.n10 GND 0.05fF
C1187 a_22576_65246.n11 GND 0.00fF
C1188 a_22576_65246.n12 GND 0.00fF
C1189 a_22576_65246.n13 GND 0.02fF
C1190 a_22576_65246.n14 GND 0.04fF
C1191 a_22576_65246.n15 GND 0.12fF
C1192 a_22576_65246.n16 GND 0.01fF
C1193 a_22576_65246.n17 GND 0.12fF
C1194 a_22576_65246.t2 GND 3.87fF $ **FLOATING
C1195 a_22576_65246.n18 GND 0.52fF
C1196 a_22576_65246.t3 GND 0.24fF $ **FLOATING
C1197 a_22866_65322.n0 GND 0.00fF
C1198 a_22866_65322.n1 GND 0.00fF
C1199 a_22866_65322.n2 GND 0.01fF
C1200 a_22866_65322.n3 GND 0.01fF
C1201 a_22866_65322.n4 GND 0.00fF
C1202 a_22866_65322.n5 GND 0.00fF
C1203 a_22866_65322.n6 GND 0.00fF
C1204 a_22866_65322.n7 GND 0.00fF
C1205 a_22866_65322.n8 GND 0.00fF
C1206 a_22866_65322.n9 GND 0.00fF
C1207 a_22866_65322.n10 GND 0.09fF
C1208 a_22866_65322.n11 GND 0.00fF
C1209 a_22866_65322.n12 GND 0.01fF
C1210 a_22866_65322.n13 GND 0.01fF
C1211 a_22866_65322.n14 GND 0.01fF
C1212 a_22866_65322.n15 GND 0.00fF
C1213 a_22866_65322.n16 GND 0.00fF
C1214 a_22866_65322.n17 GND 0.00fF
C1215 a_22866_65322.t1 GND 0.02fF $ **FLOATING
C1216 a_22866_65322.n18 GND 0.07fF
C1217 a_22866_65322.n19 GND 0.02fF
C1218 a_22866_65322.n20 GND 0.05fF
C1219 a_22866_65322.n22 GND 0.04fF
C1220 a_22866_65322.n23 GND 0.04fF
C1221 a_22866_65322.n24 GND 0.00fF
C1222 a_22866_65322.n25 GND 0.00fF
C1223 a_22866_65322.t0 GND 0.02fF $ **FLOATING
C1224 a_22866_65322.n26 GND 0.07fF
C1225 a_22866_65322.n27 GND 0.02fF
C1226 a_22866_65322.n28 GND 0.05fF
C1227 a_22866_65322.n30 GND 0.01fF
C1228 a_22866_65322.n31 GND 0.00fF
C1229 a_22866_65322.n32 GND 0.00fF
C1230 a_22866_65322.n33 GND 0.00fF
C1231 a_22866_65322.n34 GND 0.00fF
C1232 a_22866_65322.n35 GND 0.00fF
C1233 a_22866_65322.n36 GND 0.00fF
C1234 a_22866_65322.n38 GND 0.08fF
C1235 a_22866_65322.t2 GND 4.19fF $ **FLOATING
C1236 a_22866_65322.n39 GND 0.61fF
C1237 a_22866_65322.t3 GND 0.26fF $ **FLOATING
C1238 a_4466_15922.n0 GND 0.00fF
C1239 a_4466_15922.n1 GND 0.00fF
C1240 a_4466_15922.n2 GND 0.01fF
C1241 a_4466_15922.n3 GND 0.01fF
C1242 a_4466_15922.n4 GND 0.00fF
C1243 a_4466_15922.n5 GND 0.00fF
C1244 a_4466_15922.n6 GND 0.00fF
C1245 a_4466_15922.n7 GND 0.00fF
C1246 a_4466_15922.n8 GND 0.00fF
C1247 a_4466_15922.n9 GND 0.00fF
C1248 a_4466_15922.n10 GND 0.09fF
C1249 a_4466_15922.n11 GND 0.00fF
C1250 a_4466_15922.n12 GND 0.01fF
C1251 a_4466_15922.n13 GND 0.01fF
C1252 a_4466_15922.n14 GND 0.01fF
C1253 a_4466_15922.n15 GND 0.00fF
C1254 a_4466_15922.n16 GND 0.00fF
C1255 a_4466_15922.n17 GND 0.00fF
C1256 a_4466_15922.t1 GND 0.02fF $ **FLOATING
C1257 a_4466_15922.n18 GND 0.07fF
C1258 a_4466_15922.n19 GND 0.02fF
C1259 a_4466_15922.n20 GND 0.05fF
C1260 a_4466_15922.n22 GND 0.04fF
C1261 a_4466_15922.n23 GND 0.04fF
C1262 a_4466_15922.n24 GND 0.00fF
C1263 a_4466_15922.n25 GND 0.00fF
C1264 a_4466_15922.t2 GND 0.02fF $ **FLOATING
C1265 a_4466_15922.n26 GND 0.07fF
C1266 a_4466_15922.n27 GND 0.02fF
C1267 a_4466_15922.n28 GND 0.05fF
C1268 a_4466_15922.n30 GND 0.01fF
C1269 a_4466_15922.n31 GND 0.00fF
C1270 a_4466_15922.n32 GND 0.00fF
C1271 a_4466_15922.n33 GND 0.00fF
C1272 a_4466_15922.n34 GND 0.00fF
C1273 a_4466_15922.n35 GND 0.00fF
C1274 a_4466_15922.n36 GND 0.00fF
C1275 a_4466_15922.n38 GND 0.08fF
C1276 a_4466_15922.t3 GND 4.19fF $ **FLOATING
C1277 a_4466_15922.n39 GND 0.61fF
C1278 a_4466_15922.t0 GND 0.26fF $ **FLOATING
C1279 a_59376_65246.n0 GND 0.01fF
C1280 a_59376_65246.n1 GND 0.01fF
C1281 a_59376_65246.n2 GND 0.00fF
C1282 a_59376_65246.n3 GND 0.00fF
C1283 a_59376_65246.n4 GND 0.00fF
C1284 a_59376_65246.n5 GND 0.00fF
C1285 a_59376_65246.n6 GND 0.00fF
C1286 a_59376_65246.n7 GND 0.00fF
C1287 a_59376_65246.n8 GND 0.00fF
C1288 a_59376_65246.n9 GND 0.00fF
C1289 a_59376_65246.t1 GND 0.02fF $ **FLOATING
C1290 a_59376_65246.t0 GND 0.02fF $ **FLOATING
C1291 a_59376_65246.n10 GND 0.05fF
C1292 a_59376_65246.n11 GND 0.00fF
C1293 a_59376_65246.n12 GND 0.00fF
C1294 a_59376_65246.n13 GND 0.02fF
C1295 a_59376_65246.n14 GND 0.04fF
C1296 a_59376_65246.n15 GND 0.12fF
C1297 a_59376_65246.n16 GND 0.01fF
C1298 a_59376_65246.n17 GND 0.12fF
C1299 a_59376_65246.t2 GND 3.87fF $ **FLOATING
C1300 a_59376_65246.n18 GND 0.52fF
C1301 a_59376_65246.t3 GND 0.24fF $ **FLOATING
C1302 a_13666_85082.n0 GND 0.00fF
C1303 a_13666_85082.n1 GND 0.00fF
C1304 a_13666_85082.n2 GND 0.01fF
C1305 a_13666_85082.n3 GND 0.01fF
C1306 a_13666_85082.n4 GND 0.00fF
C1307 a_13666_85082.n5 GND 0.00fF
C1308 a_13666_85082.n6 GND 0.00fF
C1309 a_13666_85082.n7 GND 0.00fF
C1310 a_13666_85082.n8 GND 0.00fF
C1311 a_13666_85082.n9 GND 0.00fF
C1312 a_13666_85082.n10 GND 0.09fF
C1313 a_13666_85082.n11 GND 0.00fF
C1314 a_13666_85082.n12 GND 0.01fF
C1315 a_13666_85082.n13 GND 0.01fF
C1316 a_13666_85082.n14 GND 0.01fF
C1317 a_13666_85082.n15 GND 0.00fF
C1318 a_13666_85082.n16 GND 0.00fF
C1319 a_13666_85082.n17 GND 0.00fF
C1320 a_13666_85082.t1 GND 0.02fF $ **FLOATING
C1321 a_13666_85082.n18 GND 0.07fF
C1322 a_13666_85082.n19 GND 0.02fF
C1323 a_13666_85082.n20 GND 0.05fF
C1324 a_13666_85082.n22 GND 0.04fF
C1325 a_13666_85082.n23 GND 0.04fF
C1326 a_13666_85082.n24 GND 0.00fF
C1327 a_13666_85082.n25 GND 0.00fF
C1328 a_13666_85082.t2 GND 0.02fF $ **FLOATING
C1329 a_13666_85082.n26 GND 0.07fF
C1330 a_13666_85082.n27 GND 0.02fF
C1331 a_13666_85082.n28 GND 0.05fF
C1332 a_13666_85082.n30 GND 0.01fF
C1333 a_13666_85082.n31 GND 0.00fF
C1334 a_13666_85082.n32 GND 0.00fF
C1335 a_13666_85082.n33 GND 0.00fF
C1336 a_13666_85082.n34 GND 0.00fF
C1337 a_13666_85082.n35 GND 0.00fF
C1338 a_13666_85082.n36 GND 0.00fF
C1339 a_13666_85082.n38 GND 0.08fF
C1340 a_13666_85082.t0 GND 4.19fF $ **FLOATING
C1341 a_13666_85082.n39 GND 0.61fF
C1342 a_13666_85082.t3 GND 0.26fF $ **FLOATING
C1343 a_13376_85006.n0 GND 0.01fF
C1344 a_13376_85006.n1 GND 0.01fF
C1345 a_13376_85006.n2 GND 0.00fF
C1346 a_13376_85006.n3 GND 0.00fF
C1347 a_13376_85006.n4 GND 0.00fF
C1348 a_13376_85006.n5 GND 0.00fF
C1349 a_13376_85006.n6 GND 0.00fF
C1350 a_13376_85006.n7 GND 0.00fF
C1351 a_13376_85006.n8 GND 0.00fF
C1352 a_13376_85006.n9 GND 0.00fF
C1353 a_13376_85006.t3 GND 0.02fF $ **FLOATING
C1354 a_13376_85006.t2 GND 0.02fF $ **FLOATING
C1355 a_13376_85006.n10 GND 0.05fF
C1356 a_13376_85006.n11 GND 0.00fF
C1357 a_13376_85006.n12 GND 0.00fF
C1358 a_13376_85006.n13 GND 0.02fF
C1359 a_13376_85006.n14 GND 0.04fF
C1360 a_13376_85006.n15 GND 0.12fF
C1361 a_13376_85006.n16 GND 0.01fF
C1362 a_13376_85006.n17 GND 0.12fF
C1363 a_13376_85006.t1 GND 3.87fF $ **FLOATING
C1364 a_13376_85006.n18 GND 0.52fF
C1365 a_13376_85006.t0 GND 0.24fF $ **FLOATING
C1366 bit1.t3 GND 0.02fF $ **FLOATING
C1367 bit1.n0 GND 0.01fF
C1368 bit1.n1 GND 0.00fF
C1369 bit1.t0 GND 0.02fF $ **FLOATING
C1370 bit1.n2 GND 0.01fF
C1371 bit1.n3 GND 0.00fF
C1372 bit1.n4 GND 0.00fF
C1373 bit1.n5 GND 0.00fF
C1374 bit1.n6 GND 0.07fF
C1375 bit1.n7 GND 0.00fF
C1376 bit1.n8 GND 0.00fF
C1377 bit1.t4 GND 0.02fF $ **FLOATING
C1378 bit1.n9 GND 0.01fF
C1379 bit1.n10 GND 0.00fF
C1380 bit1.t1 GND 0.02fF $ **FLOATING
C1381 bit1.n11 GND 0.01fF
C1382 bit1.n12 GND 0.00fF
C1383 bit1.n13 GND 0.07fF
C1384 bit1.t5 GND 0.01fF $ **FLOATING
C1385 bit1.t2 GND 0.01fF $ **FLOATING
C1386 bit1.n14 GND 0.02fF
C1387 bit1.n15 GND 16.94fF
C1388 bit1.n16 GND 70.36fF
C1389 a_59376_25726.n0 GND 0.01fF
C1390 a_59376_25726.n1 GND 0.01fF
C1391 a_59376_25726.n2 GND 0.00fF
C1392 a_59376_25726.n3 GND 0.00fF
C1393 a_59376_25726.n4 GND 0.00fF
C1394 a_59376_25726.n5 GND 0.00fF
C1395 a_59376_25726.n6 GND 0.00fF
C1396 a_59376_25726.n7 GND 0.00fF
C1397 a_59376_25726.n8 GND 0.00fF
C1398 a_59376_25726.n9 GND 0.00fF
C1399 a_59376_25726.t0 GND 0.02fF $ **FLOATING
C1400 a_59376_25726.t1 GND 0.02fF $ **FLOATING
C1401 a_59376_25726.n10 GND 0.05fF
C1402 a_59376_25726.n11 GND 0.00fF
C1403 a_59376_25726.n12 GND 0.00fF
C1404 a_59376_25726.n13 GND 0.02fF
C1405 a_59376_25726.n14 GND 0.04fF
C1406 a_59376_25726.n15 GND 0.12fF
C1407 a_59376_25726.n16 GND 0.01fF
C1408 a_59376_25726.n17 GND 0.12fF
C1409 a_59376_25726.t2 GND 3.87fF $ **FLOATING
C1410 a_59376_25726.n18 GND 0.52fF
C1411 a_59376_25726.t3 GND 0.24fF $ **FLOATING
C1412 a_59666_25802.n0 GND 0.00fF
C1413 a_59666_25802.n1 GND 0.00fF
C1414 a_59666_25802.n2 GND 0.01fF
C1415 a_59666_25802.n3 GND 0.01fF
C1416 a_59666_25802.n4 GND 0.00fF
C1417 a_59666_25802.n5 GND 0.00fF
C1418 a_59666_25802.n6 GND 0.00fF
C1419 a_59666_25802.n7 GND 0.00fF
C1420 a_59666_25802.n8 GND 0.00fF
C1421 a_59666_25802.n9 GND 0.00fF
C1422 a_59666_25802.n10 GND 0.09fF
C1423 a_59666_25802.n11 GND 0.00fF
C1424 a_59666_25802.n12 GND 0.01fF
C1425 a_59666_25802.n13 GND 0.01fF
C1426 a_59666_25802.n14 GND 0.01fF
C1427 a_59666_25802.n15 GND 0.00fF
C1428 a_59666_25802.n16 GND 0.00fF
C1429 a_59666_25802.n17 GND 0.00fF
C1430 a_59666_25802.t0 GND 0.02fF $ **FLOATING
C1431 a_59666_25802.n18 GND 0.07fF
C1432 a_59666_25802.n19 GND 0.02fF
C1433 a_59666_25802.n20 GND 0.05fF
C1434 a_59666_25802.n22 GND 0.04fF
C1435 a_59666_25802.n23 GND 0.04fF
C1436 a_59666_25802.n24 GND 0.00fF
C1437 a_59666_25802.n25 GND 0.00fF
C1438 a_59666_25802.t1 GND 0.02fF $ **FLOATING
C1439 a_59666_25802.n26 GND 0.07fF
C1440 a_59666_25802.n27 GND 0.02fF
C1441 a_59666_25802.n28 GND 0.05fF
C1442 a_59666_25802.n30 GND 0.01fF
C1443 a_59666_25802.n31 GND 0.00fF
C1444 a_59666_25802.n32 GND 0.00fF
C1445 a_59666_25802.n33 GND 0.00fF
C1446 a_59666_25802.n34 GND 0.00fF
C1447 a_59666_25802.n35 GND 0.00fF
C1448 a_59666_25802.n36 GND 0.00fF
C1449 a_59666_25802.n38 GND 0.08fF
C1450 a_59666_25802.t3 GND 4.19fF $ **FLOATING
C1451 a_59666_25802.n39 GND 0.61fF
C1452 a_59666_25802.t2 GND 0.26fF $ **FLOATING
C1453 a_4466_85082.n0 GND 0.00fF
C1454 a_4466_85082.n1 GND 0.00fF
C1455 a_4466_85082.n2 GND 0.01fF
C1456 a_4466_85082.n3 GND 0.01fF
C1457 a_4466_85082.n4 GND 0.00fF
C1458 a_4466_85082.n5 GND 0.00fF
C1459 a_4466_85082.n6 GND 0.00fF
C1460 a_4466_85082.n7 GND 0.00fF
C1461 a_4466_85082.n8 GND 0.00fF
C1462 a_4466_85082.n9 GND 0.00fF
C1463 a_4466_85082.n10 GND 0.09fF
C1464 a_4466_85082.n11 GND 0.00fF
C1465 a_4466_85082.n12 GND 0.01fF
C1466 a_4466_85082.n13 GND 0.01fF
C1467 a_4466_85082.n14 GND 0.01fF
C1468 a_4466_85082.n15 GND 0.00fF
C1469 a_4466_85082.n16 GND 0.00fF
C1470 a_4466_85082.n17 GND 0.00fF
C1471 a_4466_85082.t3 GND 0.02fF $ **FLOATING
C1472 a_4466_85082.n18 GND 0.07fF
C1473 a_4466_85082.n19 GND 0.02fF
C1474 a_4466_85082.n20 GND 0.05fF
C1475 a_4466_85082.n22 GND 0.04fF
C1476 a_4466_85082.n23 GND 0.04fF
C1477 a_4466_85082.n24 GND 0.00fF
C1478 a_4466_85082.n25 GND 0.00fF
C1479 a_4466_85082.t2 GND 0.02fF $ **FLOATING
C1480 a_4466_85082.n26 GND 0.07fF
C1481 a_4466_85082.n27 GND 0.02fF
C1482 a_4466_85082.n28 GND 0.05fF
C1483 a_4466_85082.n30 GND 0.01fF
C1484 a_4466_85082.n31 GND 0.00fF
C1485 a_4466_85082.n32 GND 0.00fF
C1486 a_4466_85082.n33 GND 0.00fF
C1487 a_4466_85082.n34 GND 0.00fF
C1488 a_4466_85082.n35 GND 0.00fF
C1489 a_4466_85082.n36 GND 0.00fF
C1490 a_4466_85082.n38 GND 0.08fF
C1491 a_4466_85082.t0 GND 4.19fF $ **FLOATING
C1492 a_4466_85082.n39 GND 0.61fF
C1493 a_4466_85082.t1 GND 0.26fF $ **FLOATING
C1494 a_68576_65246.n0 GND 0.01fF
C1495 a_68576_65246.n1 GND 0.01fF
C1496 a_68576_65246.n2 GND 0.00fF
C1497 a_68576_65246.n3 GND 0.00fF
C1498 a_68576_65246.n4 GND 0.00fF
C1499 a_68576_65246.n5 GND 0.00fF
C1500 a_68576_65246.n6 GND 0.00fF
C1501 a_68576_65246.n7 GND 0.00fF
C1502 a_68576_65246.n8 GND 0.00fF
C1503 a_68576_65246.n9 GND 0.00fF
C1504 a_68576_65246.t1 GND 0.02fF $ **FLOATING
C1505 a_68576_65246.t0 GND 0.02fF $ **FLOATING
C1506 a_68576_65246.n10 GND 0.05fF
C1507 a_68576_65246.n11 GND 0.00fF
C1508 a_68576_65246.n12 GND 0.00fF
C1509 a_68576_65246.n13 GND 0.02fF
C1510 a_68576_65246.n14 GND 0.04fF
C1511 a_68576_65246.n15 GND 0.12fF
C1512 a_68576_65246.n16 GND 0.01fF
C1513 a_68576_65246.n17 GND 0.12fF
C1514 a_68576_65246.t2 GND 3.87fF $ **FLOATING
C1515 a_68576_65246.n18 GND 0.52fF
C1516 a_68576_65246.t3 GND 0.24fF $ **FLOATING
C1517 a_40976_65246.n0 GND 0.01fF
C1518 a_40976_65246.n1 GND 0.01fF
C1519 a_40976_65246.n2 GND 0.00fF
C1520 a_40976_65246.n3 GND 0.00fF
C1521 a_40976_65246.n4 GND 0.00fF
C1522 a_40976_65246.n5 GND 0.00fF
C1523 a_40976_65246.n6 GND 0.00fF
C1524 a_40976_65246.n7 GND 0.00fF
C1525 a_40976_65246.n8 GND 0.00fF
C1526 a_40976_65246.n9 GND 0.00fF
C1527 a_40976_65246.t0 GND 0.02fF $ **FLOATING
C1528 a_40976_65246.t1 GND 0.02fF $ **FLOATING
C1529 a_40976_65246.n10 GND 0.05fF
C1530 a_40976_65246.n11 GND 0.00fF
C1531 a_40976_65246.n12 GND 0.00fF
C1532 a_40976_65246.n13 GND 0.02fF
C1533 a_40976_65246.n14 GND 0.04fF
C1534 a_40976_65246.n15 GND 0.12fF
C1535 a_40976_65246.n16 GND 0.01fF
C1536 a_40976_65246.n17 GND 0.12fF
C1537 a_40976_65246.t3 GND 3.87fF $ **FLOATING
C1538 a_40976_65246.n18 GND 0.52fF
C1539 a_40976_65246.t2 GND 0.24fF $ **FLOATING
C1540 a_41266_65322.n0 GND 0.00fF
C1541 a_41266_65322.n1 GND 0.00fF
C1542 a_41266_65322.n2 GND 0.01fF
C1543 a_41266_65322.n3 GND 0.01fF
C1544 a_41266_65322.n4 GND 0.00fF
C1545 a_41266_65322.n5 GND 0.00fF
C1546 a_41266_65322.n6 GND 0.00fF
C1547 a_41266_65322.n7 GND 0.00fF
C1548 a_41266_65322.n8 GND 0.00fF
C1549 a_41266_65322.n9 GND 0.00fF
C1550 a_41266_65322.n10 GND 0.09fF
C1551 a_41266_65322.n11 GND 0.00fF
C1552 a_41266_65322.n12 GND 0.01fF
C1553 a_41266_65322.n13 GND 0.01fF
C1554 a_41266_65322.n14 GND 0.01fF
C1555 a_41266_65322.n15 GND 0.00fF
C1556 a_41266_65322.n16 GND 0.00fF
C1557 a_41266_65322.n17 GND 0.00fF
C1558 a_41266_65322.t2 GND 0.02fF $ **FLOATING
C1559 a_41266_65322.n18 GND 0.07fF
C1560 a_41266_65322.n19 GND 0.02fF
C1561 a_41266_65322.n20 GND 0.05fF
C1562 a_41266_65322.n22 GND 0.04fF
C1563 a_41266_65322.n23 GND 0.04fF
C1564 a_41266_65322.n24 GND 0.00fF
C1565 a_41266_65322.n25 GND 0.00fF
C1566 a_41266_65322.t1 GND 0.02fF $ **FLOATING
C1567 a_41266_65322.n26 GND 0.07fF
C1568 a_41266_65322.n27 GND 0.02fF
C1569 a_41266_65322.n28 GND 0.05fF
C1570 a_41266_65322.n30 GND 0.01fF
C1571 a_41266_65322.n31 GND 0.00fF
C1572 a_41266_65322.n32 GND 0.00fF
C1573 a_41266_65322.n33 GND 0.00fF
C1574 a_41266_65322.n34 GND 0.00fF
C1575 a_41266_65322.n35 GND 0.00fF
C1576 a_41266_65322.n36 GND 0.00fF
C1577 a_41266_65322.n38 GND 0.08fF
C1578 a_41266_65322.t3 GND 4.19fF $ **FLOATING
C1579 a_41266_65322.n39 GND 0.61fF
C1580 a_41266_65322.t0 GND 0.26fF $ **FLOATING
C1581 a_50466_25802.n0 GND 0.00fF
C1582 a_50466_25802.n1 GND 0.00fF
C1583 a_50466_25802.n2 GND 0.01fF
C1584 a_50466_25802.n3 GND 0.01fF
C1585 a_50466_25802.n4 GND 0.00fF
C1586 a_50466_25802.n5 GND 0.00fF
C1587 a_50466_25802.n6 GND 0.00fF
C1588 a_50466_25802.n7 GND 0.00fF
C1589 a_50466_25802.n8 GND 0.00fF
C1590 a_50466_25802.n9 GND 0.00fF
C1591 a_50466_25802.n10 GND 0.09fF
C1592 a_50466_25802.n11 GND 0.00fF
C1593 a_50466_25802.n12 GND 0.01fF
C1594 a_50466_25802.n13 GND 0.01fF
C1595 a_50466_25802.n14 GND 0.01fF
C1596 a_50466_25802.n15 GND 0.00fF
C1597 a_50466_25802.n16 GND 0.00fF
C1598 a_50466_25802.n17 GND 0.00fF
C1599 a_50466_25802.t0 GND 0.02fF $ **FLOATING
C1600 a_50466_25802.n18 GND 0.07fF
C1601 a_50466_25802.n19 GND 0.02fF
C1602 a_50466_25802.n20 GND 0.05fF
C1603 a_50466_25802.n22 GND 0.04fF
C1604 a_50466_25802.n23 GND 0.04fF
C1605 a_50466_25802.n24 GND 0.00fF
C1606 a_50466_25802.n25 GND 0.00fF
C1607 a_50466_25802.t1 GND 0.02fF $ **FLOATING
C1608 a_50466_25802.n26 GND 0.07fF
C1609 a_50466_25802.n27 GND 0.02fF
C1610 a_50466_25802.n28 GND 0.05fF
C1611 a_50466_25802.n30 GND 0.01fF
C1612 a_50466_25802.n31 GND 0.00fF
C1613 a_50466_25802.n32 GND 0.00fF
C1614 a_50466_25802.n33 GND 0.00fF
C1615 a_50466_25802.n34 GND 0.00fF
C1616 a_50466_25802.n35 GND 0.00fF
C1617 a_50466_25802.n36 GND 0.00fF
C1618 a_50466_25802.n38 GND 0.08fF
C1619 a_50466_25802.t2 GND 4.19fF $ **FLOATING
C1620 a_50466_25802.n39 GND 0.61fF
C1621 a_50466_25802.t3 GND 0.26fF $ **FLOATING
C1622 a_50176_25726.n0 GND 0.01fF
C1623 a_50176_25726.n1 GND 0.01fF
C1624 a_50176_25726.n2 GND 0.00fF
C1625 a_50176_25726.n3 GND 0.00fF
C1626 a_50176_25726.n4 GND 0.00fF
C1627 a_50176_25726.n5 GND 0.00fF
C1628 a_50176_25726.n6 GND 0.00fF
C1629 a_50176_25726.n7 GND 0.00fF
C1630 a_50176_25726.n8 GND 0.00fF
C1631 a_50176_25726.n9 GND 0.00fF
C1632 a_50176_25726.t1 GND 0.02fF $ **FLOATING
C1633 a_50176_25726.t0 GND 0.02fF $ **FLOATING
C1634 a_50176_25726.n10 GND 0.05fF
C1635 a_50176_25726.n11 GND 0.00fF
C1636 a_50176_25726.n12 GND 0.00fF
C1637 a_50176_25726.n13 GND 0.02fF
C1638 a_50176_25726.n14 GND 0.04fF
C1639 a_50176_25726.n15 GND 0.12fF
C1640 a_50176_25726.n16 GND 0.01fF
C1641 a_50176_25726.n17 GND 0.12fF
C1642 a_50176_25726.t2 GND 3.87fF $ **FLOATING
C1643 a_50176_25726.n18 GND 0.52fF
C1644 a_50176_25726.t3 GND 0.24fF $ **FLOATING
C1645 a_68576_45486.n0 GND 0.01fF
C1646 a_68576_45486.n1 GND 0.01fF
C1647 a_68576_45486.n2 GND 0.00fF
C1648 a_68576_45486.n3 GND 0.00fF
C1649 a_68576_45486.n4 GND 0.00fF
C1650 a_68576_45486.n5 GND 0.00fF
C1651 a_68576_45486.n6 GND 0.00fF
C1652 a_68576_45486.n7 GND 0.00fF
C1653 a_68576_45486.n8 GND 0.00fF
C1654 a_68576_45486.n9 GND 0.00fF
C1655 a_68576_45486.t1 GND 0.02fF $ **FLOATING
C1656 a_68576_45486.t0 GND 0.02fF $ **FLOATING
C1657 a_68576_45486.n10 GND 0.05fF
C1658 a_68576_45486.n11 GND 0.00fF
C1659 a_68576_45486.n12 GND 0.00fF
C1660 a_68576_45486.n13 GND 0.02fF
C1661 a_68576_45486.n14 GND 0.04fF
C1662 a_68576_45486.n15 GND 0.12fF
C1663 a_68576_45486.n16 GND 0.01fF
C1664 a_68576_45486.n17 GND 0.12fF
C1665 a_68576_45486.t2 GND 3.87fF $ **FLOATING
C1666 a_68576_45486.n18 GND 0.52fF
C1667 a_68576_45486.t3 GND 0.24fF $ **FLOATING
C1668 a_40976_35606.n0 GND 0.01fF
C1669 a_40976_35606.n1 GND 0.01fF
C1670 a_40976_35606.n2 GND 0.00fF
C1671 a_40976_35606.n3 GND 0.00fF
C1672 a_40976_35606.n4 GND 0.00fF
C1673 a_40976_35606.n5 GND 0.00fF
C1674 a_40976_35606.n6 GND 0.00fF
C1675 a_40976_35606.n7 GND 0.00fF
C1676 a_40976_35606.n8 GND 0.00fF
C1677 a_40976_35606.n9 GND 0.00fF
C1678 a_40976_35606.t2 GND 0.02fF $ **FLOATING
C1679 a_40976_35606.t1 GND 0.02fF $ **FLOATING
C1680 a_40976_35606.n10 GND 0.05fF
C1681 a_40976_35606.n11 GND 0.00fF
C1682 a_40976_35606.n12 GND 0.00fF
C1683 a_40976_35606.n13 GND 0.02fF
C1684 a_40976_35606.n14 GND 0.04fF
C1685 a_40976_35606.n15 GND 0.12fF
C1686 a_40976_35606.n16 GND 0.01fF
C1687 a_40976_35606.n17 GND 0.12fF
C1688 a_40976_35606.t3 GND 3.87fF $ **FLOATING
C1689 a_40976_35606.n18 GND 0.52fF
C1690 a_40976_35606.t0 GND 0.24fF $ **FLOATING
C1691 a_13666_6042.n0 GND 0.00fF
C1692 a_13666_6042.n1 GND 0.00fF
C1693 a_13666_6042.n2 GND 0.01fF
C1694 a_13666_6042.n3 GND 0.01fF
C1695 a_13666_6042.n4 GND 0.00fF
C1696 a_13666_6042.n5 GND 0.00fF
C1697 a_13666_6042.n6 GND 0.00fF
C1698 a_13666_6042.n7 GND 0.00fF
C1699 a_13666_6042.n8 GND 0.00fF
C1700 a_13666_6042.n9 GND 0.00fF
C1701 a_13666_6042.n10 GND 0.09fF
C1702 a_13666_6042.n11 GND 0.00fF
C1703 a_13666_6042.n12 GND 0.01fF
C1704 a_13666_6042.n13 GND 0.01fF
C1705 a_13666_6042.n14 GND 0.01fF
C1706 a_13666_6042.n15 GND 0.00fF
C1707 a_13666_6042.n16 GND 0.00fF
C1708 a_13666_6042.n17 GND 0.00fF
C1709 a_13666_6042.t0 GND 0.02fF $ **FLOATING
C1710 a_13666_6042.n18 GND 0.07fF
C1711 a_13666_6042.n19 GND 0.02fF
C1712 a_13666_6042.n20 GND 0.05fF
C1713 a_13666_6042.n22 GND 0.04fF
C1714 a_13666_6042.n23 GND 0.04fF
C1715 a_13666_6042.n24 GND 0.00fF
C1716 a_13666_6042.n25 GND 0.00fF
C1717 a_13666_6042.t1 GND 0.02fF $ **FLOATING
C1718 a_13666_6042.n26 GND 0.07fF
C1719 a_13666_6042.n27 GND 0.02fF
C1720 a_13666_6042.n28 GND 0.05fF
C1721 a_13666_6042.n30 GND 0.01fF
C1722 a_13666_6042.n31 GND 0.00fF
C1723 a_13666_6042.n32 GND 0.00fF
C1724 a_13666_6042.n33 GND 0.00fF
C1725 a_13666_6042.n34 GND 0.00fF
C1726 a_13666_6042.n35 GND 0.00fF
C1727 a_13666_6042.n36 GND 0.00fF
C1728 a_13666_6042.n38 GND 0.08fF
C1729 a_13666_6042.t2 GND 4.19fF $ **FLOATING
C1730 a_13666_6042.n39 GND 0.61fF
C1731 a_13666_6042.t3 GND 0.26fF $ **FLOATING
C1732 a_13376_5966.n0 GND 0.01fF
C1733 a_13376_5966.n1 GND 0.01fF
C1734 a_13376_5966.n2 GND 0.00fF
C1735 a_13376_5966.n3 GND 0.00fF
C1736 a_13376_5966.n4 GND 0.00fF
C1737 a_13376_5966.n5 GND 0.00fF
C1738 a_13376_5966.n6 GND 0.00fF
C1739 a_13376_5966.n7 GND 0.00fF
C1740 a_13376_5966.n8 GND 0.00fF
C1741 a_13376_5966.n9 GND 0.00fF
C1742 a_13376_5966.t1 GND 0.02fF $ **FLOATING
C1743 a_13376_5966.t0 GND 0.02fF $ **FLOATING
C1744 a_13376_5966.n10 GND 0.05fF
C1745 a_13376_5966.n11 GND 0.00fF
C1746 a_13376_5966.n12 GND 0.00fF
C1747 a_13376_5966.n13 GND 0.02fF
C1748 a_13376_5966.n14 GND 0.04fF
C1749 a_13376_5966.n15 GND 0.12fF
C1750 a_13376_5966.n16 GND 0.01fF
C1751 a_13376_5966.n17 GND 0.12fF
C1752 a_13376_5966.t2 GND 3.87fF $ **FLOATING
C1753 a_13376_5966.n18 GND 0.52fF
C1754 a_13376_5966.t3 GND 0.24fF $ **FLOATING
C1755 a_59666_6042.n0 GND 0.00fF
C1756 a_59666_6042.n1 GND 0.00fF
C1757 a_59666_6042.n2 GND 0.01fF
C1758 a_59666_6042.n3 GND 0.01fF
C1759 a_59666_6042.n4 GND 0.00fF
C1760 a_59666_6042.n5 GND 0.00fF
C1761 a_59666_6042.n6 GND 0.00fF
C1762 a_59666_6042.n7 GND 0.00fF
C1763 a_59666_6042.n8 GND 0.00fF
C1764 a_59666_6042.n9 GND 0.00fF
C1765 a_59666_6042.n10 GND 0.09fF
C1766 a_59666_6042.n11 GND 0.00fF
C1767 a_59666_6042.n12 GND 0.01fF
C1768 a_59666_6042.n13 GND 0.01fF
C1769 a_59666_6042.n14 GND 0.01fF
C1770 a_59666_6042.n15 GND 0.00fF
C1771 a_59666_6042.n16 GND 0.00fF
C1772 a_59666_6042.n17 GND 0.00fF
C1773 a_59666_6042.t1 GND 0.02fF $ **FLOATING
C1774 a_59666_6042.n18 GND 0.07fF
C1775 a_59666_6042.n19 GND 0.02fF
C1776 a_59666_6042.n20 GND 0.05fF
C1777 a_59666_6042.n22 GND 0.04fF
C1778 a_59666_6042.n23 GND 0.04fF
C1779 a_59666_6042.n24 GND 0.00fF
C1780 a_59666_6042.n25 GND 0.00fF
C1781 a_59666_6042.t2 GND 0.02fF $ **FLOATING
C1782 a_59666_6042.n26 GND 0.07fF
C1783 a_59666_6042.n27 GND 0.02fF
C1784 a_59666_6042.n28 GND 0.05fF
C1785 a_59666_6042.n30 GND 0.01fF
C1786 a_59666_6042.n31 GND 0.00fF
C1787 a_59666_6042.n32 GND 0.00fF
C1788 a_59666_6042.n33 GND 0.00fF
C1789 a_59666_6042.n34 GND 0.00fF
C1790 a_59666_6042.n35 GND 0.00fF
C1791 a_59666_6042.n36 GND 0.00fF
C1792 a_59666_6042.n38 GND 0.08fF
C1793 a_59666_6042.t3 GND 4.19fF $ **FLOATING
C1794 a_59666_6042.n39 GND 0.61fF
C1795 a_59666_6042.t0 GND 0.26fF $ **FLOATING
C1796 a_4176_85006.n0 GND 0.01fF
C1797 a_4176_85006.n1 GND 0.01fF
C1798 a_4176_85006.n2 GND 0.00fF
C1799 a_4176_85006.n3 GND 0.00fF
C1800 a_4176_85006.n4 GND 0.00fF
C1801 a_4176_85006.n5 GND 0.00fF
C1802 a_4176_85006.n6 GND 0.00fF
C1803 a_4176_85006.n7 GND 0.00fF
C1804 a_4176_85006.n8 GND 0.00fF
C1805 a_4176_85006.n9 GND 0.00fF
C1806 a_4176_85006.t2 GND 0.02fF $ **FLOATING
C1807 a_4176_85006.t3 GND 0.02fF $ **FLOATING
C1808 a_4176_85006.n10 GND 0.05fF
C1809 a_4176_85006.n11 GND 0.00fF
C1810 a_4176_85006.n12 GND 0.00fF
C1811 a_4176_85006.n13 GND 0.02fF
C1812 a_4176_85006.n14 GND 0.04fF
C1813 a_4176_85006.n15 GND 0.12fF
C1814 a_4176_85006.n16 GND 0.01fF
C1815 a_4176_85006.n17 GND 0.12fF
C1816 a_4176_85006.t0 GND 3.87fF $ **FLOATING
C1817 a_4176_85006.n18 GND 0.52fF
C1818 a_4176_85006.t1 GND 0.24fF $ **FLOATING
C1819 a_68576_5966.n0 GND 0.01fF
C1820 a_68576_5966.n1 GND 0.01fF
C1821 a_68576_5966.n2 GND 0.00fF
C1822 a_68576_5966.n3 GND 0.00fF
C1823 a_68576_5966.n4 GND 0.00fF
C1824 a_68576_5966.n5 GND 0.00fF
C1825 a_68576_5966.n6 GND 0.00fF
C1826 a_68576_5966.n7 GND 0.00fF
C1827 a_68576_5966.n8 GND 0.00fF
C1828 a_68576_5966.n9 GND 0.00fF
C1829 a_68576_5966.t1 GND 0.02fF $ **FLOATING
C1830 a_68576_5966.t2 GND 0.02fF $ **FLOATING
C1831 a_68576_5966.n10 GND 0.05fF
C1832 a_68576_5966.n11 GND 0.00fF
C1833 a_68576_5966.n12 GND 0.00fF
C1834 a_68576_5966.n13 GND 0.02fF
C1835 a_68576_5966.n14 GND 0.04fF
C1836 a_68576_5966.n15 GND 0.12fF
C1837 a_68576_5966.n16 GND 0.01fF
C1838 a_68576_5966.n17 GND 0.12fF
C1839 a_68576_5966.t3 GND 3.87fF $ **FLOATING
C1840 a_68576_5966.n18 GND 0.52fF
C1841 a_68576_5966.t0 GND 0.24fF $ **FLOATING
C1842 a_68576_55366.n0 GND 0.01fF
C1843 a_68576_55366.n1 GND 0.01fF
C1844 a_68576_55366.n2 GND 0.00fF
C1845 a_68576_55366.n3 GND 0.00fF
C1846 a_68576_55366.n4 GND 0.00fF
C1847 a_68576_55366.n5 GND 0.00fF
C1848 a_68576_55366.n6 GND 0.00fF
C1849 a_68576_55366.n7 GND 0.00fF
C1850 a_68576_55366.n8 GND 0.00fF
C1851 a_68576_55366.n9 GND 0.00fF
C1852 a_68576_55366.t1 GND 0.02fF $ **FLOATING
C1853 a_68576_55366.t0 GND 0.02fF $ **FLOATING
C1854 a_68576_55366.n10 GND 0.05fF
C1855 a_68576_55366.n11 GND 0.00fF
C1856 a_68576_55366.n12 GND 0.00fF
C1857 a_68576_55366.n13 GND 0.02fF
C1858 a_68576_55366.n14 GND 0.04fF
C1859 a_68576_55366.n15 GND 0.12fF
C1860 a_68576_55366.n16 GND 0.01fF
C1861 a_68576_55366.n17 GND 0.12fF
C1862 a_68576_55366.t2 GND 3.87fF $ **FLOATING
C1863 a_68576_55366.n18 GND 0.52fF
C1864 a_68576_55366.t3 GND 0.24fF $ **FLOATING
C1865 a_4176_45486.n0 GND 0.01fF
C1866 a_4176_45486.n1 GND 0.01fF
C1867 a_4176_45486.n2 GND 0.00fF
C1868 a_4176_45486.n3 GND 0.00fF
C1869 a_4176_45486.n4 GND 0.00fF
C1870 a_4176_45486.n5 GND 0.00fF
C1871 a_4176_45486.n6 GND 0.00fF
C1872 a_4176_45486.n7 GND 0.00fF
C1873 a_4176_45486.n8 GND 0.00fF
C1874 a_4176_45486.n9 GND 0.00fF
C1875 a_4176_45486.t0 GND 0.02fF $ **FLOATING
C1876 a_4176_45486.t1 GND 0.02fF $ **FLOATING
C1877 a_4176_45486.n10 GND 0.05fF
C1878 a_4176_45486.n11 GND 0.00fF
C1879 a_4176_45486.n12 GND 0.00fF
C1880 a_4176_45486.n13 GND 0.02fF
C1881 a_4176_45486.n14 GND 0.04fF
C1882 a_4176_45486.n15 GND 0.12fF
C1883 a_4176_45486.n16 GND 0.01fF
C1884 a_4176_45486.n17 GND 0.12fF
C1885 a_4176_45486.t3 GND 3.87fF $ **FLOATING
C1886 a_4176_45486.n18 GND 0.52fF
C1887 a_4176_45486.t2 GND 0.24fF $ **FLOATING
C1888 a_4466_45562.n0 GND 0.00fF
C1889 a_4466_45562.n1 GND 0.00fF
C1890 a_4466_45562.n2 GND 0.01fF
C1891 a_4466_45562.n3 GND 0.01fF
C1892 a_4466_45562.n4 GND 0.00fF
C1893 a_4466_45562.n5 GND 0.00fF
C1894 a_4466_45562.n6 GND 0.00fF
C1895 a_4466_45562.n7 GND 0.00fF
C1896 a_4466_45562.n8 GND 0.00fF
C1897 a_4466_45562.n9 GND 0.00fF
C1898 a_4466_45562.n10 GND 0.09fF
C1899 a_4466_45562.n11 GND 0.00fF
C1900 a_4466_45562.n12 GND 0.01fF
C1901 a_4466_45562.n13 GND 0.01fF
C1902 a_4466_45562.n14 GND 0.01fF
C1903 a_4466_45562.n15 GND 0.00fF
C1904 a_4466_45562.n16 GND 0.00fF
C1905 a_4466_45562.n17 GND 0.00fF
C1906 a_4466_45562.t1 GND 0.02fF $ **FLOATING
C1907 a_4466_45562.n18 GND 0.07fF
C1908 a_4466_45562.n19 GND 0.02fF
C1909 a_4466_45562.n20 GND 0.05fF
C1910 a_4466_45562.n22 GND 0.04fF
C1911 a_4466_45562.n23 GND 0.04fF
C1912 a_4466_45562.n24 GND 0.00fF
C1913 a_4466_45562.n25 GND 0.00fF
C1914 a_4466_45562.t0 GND 0.02fF $ **FLOATING
C1915 a_4466_45562.n26 GND 0.07fF
C1916 a_4466_45562.n27 GND 0.02fF
C1917 a_4466_45562.n28 GND 0.05fF
C1918 a_4466_45562.n30 GND 0.01fF
C1919 a_4466_45562.n31 GND 0.00fF
C1920 a_4466_45562.n32 GND 0.00fF
C1921 a_4466_45562.n33 GND 0.00fF
C1922 a_4466_45562.n34 GND 0.00fF
C1923 a_4466_45562.n35 GND 0.00fF
C1924 a_4466_45562.n36 GND 0.00fF
C1925 a_4466_45562.n38 GND 0.08fF
C1926 a_4466_45562.t2 GND 4.19fF $ **FLOATING
C1927 a_4466_45562.n39 GND 0.61fF
C1928 a_4466_45562.t3 GND 0.26fF $ **FLOATING
C1929 a_n436_74606.t3 GND 0.04fF $ **FLOATING
C1930 a_n436_74606.t6 GND 0.07fF $ **FLOATING
C1931 a_n436_74606.t9 GND 0.07fF $ **FLOATING
C1932 a_n436_74606.t5 GND 0.07fF $ **FLOATING
C1933 a_n436_74606.t0 GND 0.07fF $ **FLOATING
C1934 a_n436_74606.t2 GND 0.07fF $ **FLOATING
C1935 a_n436_74606.t7 GND 0.07fF $ **FLOATING
C1936 a_n436_74606.t1 GND 0.07fF $ **FLOATING
C1937 a_n436_74606.t8 GND 0.12fF $ **FLOATING
C1938 a_n436_74606.n0 GND 21.43fF
C1939 a_n436_74606.n1 GND 10.72fF
C1940 a_n436_74606.n2 GND 10.72fF
C1941 a_n436_74606.n3 GND 10.72fF
C1942 a_n436_74606.n4 GND 10.72fF
C1943 a_n436_74606.n5 GND 10.72fF
C1944 a_n436_74606.n6 GND 12.14fF
C1945 a_n436_74606.n7 GND 0.06fF
C1946 a_n436_74606.t4 GND 0.09fF $ **FLOATING
C1947 a_68576_15846.n0 GND 0.01fF
C1948 a_68576_15846.n1 GND 0.01fF
C1949 a_68576_15846.n2 GND 0.00fF
C1950 a_68576_15846.n3 GND 0.00fF
C1951 a_68576_15846.n4 GND 0.00fF
C1952 a_68576_15846.n5 GND 0.00fF
C1953 a_68576_15846.n6 GND 0.00fF
C1954 a_68576_15846.n7 GND 0.00fF
C1955 a_68576_15846.n8 GND 0.00fF
C1956 a_68576_15846.n9 GND 0.00fF
C1957 a_68576_15846.t0 GND 0.02fF $ **FLOATING
C1958 a_68576_15846.t1 GND 0.02fF $ **FLOATING
C1959 a_68576_15846.n10 GND 0.05fF
C1960 a_68576_15846.n11 GND 0.00fF
C1961 a_68576_15846.n12 GND 0.00fF
C1962 a_68576_15846.n13 GND 0.02fF
C1963 a_68576_15846.n14 GND 0.04fF
C1964 a_68576_15846.n15 GND 0.12fF
C1965 a_68576_15846.n16 GND 0.01fF
C1966 a_68576_15846.n17 GND 0.12fF
C1967 a_68576_15846.t3 GND 3.87fF $ **FLOATING
C1968 a_68576_15846.n18 GND 0.52fF
C1969 a_68576_15846.t2 GND 0.24fF $ **FLOATING
C1970 a_68866_15922.n0 GND 0.00fF
C1971 a_68866_15922.n1 GND 0.00fF
C1972 a_68866_15922.n2 GND 0.01fF
C1973 a_68866_15922.n3 GND 0.01fF
C1974 a_68866_15922.n4 GND 0.00fF
C1975 a_68866_15922.n5 GND 0.00fF
C1976 a_68866_15922.n6 GND 0.00fF
C1977 a_68866_15922.n7 GND 0.00fF
C1978 a_68866_15922.n8 GND 0.00fF
C1979 a_68866_15922.n9 GND 0.00fF
C1980 a_68866_15922.n10 GND 0.09fF
C1981 a_68866_15922.n11 GND 0.00fF
C1982 a_68866_15922.n12 GND 0.01fF
C1983 a_68866_15922.n13 GND 0.01fF
C1984 a_68866_15922.n14 GND 0.01fF
C1985 a_68866_15922.n15 GND 0.00fF
C1986 a_68866_15922.n16 GND 0.00fF
C1987 a_68866_15922.n17 GND 0.00fF
C1988 a_68866_15922.t0 GND 0.02fF $ **FLOATING
C1989 a_68866_15922.n18 GND 0.07fF
C1990 a_68866_15922.n19 GND 0.02fF
C1991 a_68866_15922.n20 GND 0.05fF
C1992 a_68866_15922.n22 GND 0.04fF
C1993 a_68866_15922.n23 GND 0.04fF
C1994 a_68866_15922.n24 GND 0.00fF
C1995 a_68866_15922.n25 GND 0.00fF
C1996 a_68866_15922.t1 GND 0.02fF $ **FLOATING
C1997 a_68866_15922.n26 GND 0.07fF
C1998 a_68866_15922.n27 GND 0.02fF
C1999 a_68866_15922.n28 GND 0.05fF
C2000 a_68866_15922.n30 GND 0.01fF
C2001 a_68866_15922.n31 GND 0.00fF
C2002 a_68866_15922.n32 GND 0.00fF
C2003 a_68866_15922.n33 GND 0.00fF
C2004 a_68866_15922.n34 GND 0.00fF
C2005 a_68866_15922.n35 GND 0.00fF
C2006 a_68866_15922.n36 GND 0.00fF
C2007 a_68866_15922.n38 GND 0.08fF
C2008 a_68866_15922.t2 GND 4.19fF $ **FLOATING
C2009 a_68866_15922.n39 GND 0.61fF
C2010 a_68866_15922.t3 GND 0.26fF $ **FLOATING
C2011 a_59666_35682.n0 GND 0.00fF
C2012 a_59666_35682.n1 GND 0.00fF
C2013 a_59666_35682.n2 GND 0.01fF
C2014 a_59666_35682.n3 GND 0.01fF
C2015 a_59666_35682.n4 GND 0.00fF
C2016 a_59666_35682.n5 GND 0.00fF
C2017 a_59666_35682.n6 GND 0.00fF
C2018 a_59666_35682.n7 GND 0.00fF
C2019 a_59666_35682.n8 GND 0.00fF
C2020 a_59666_35682.n9 GND 0.00fF
C2021 a_59666_35682.n10 GND 0.09fF
C2022 a_59666_35682.n11 GND 0.00fF
C2023 a_59666_35682.n12 GND 0.01fF
C2024 a_59666_35682.n13 GND 0.01fF
C2025 a_59666_35682.n14 GND 0.01fF
C2026 a_59666_35682.n15 GND 0.00fF
C2027 a_59666_35682.n16 GND 0.00fF
C2028 a_59666_35682.n17 GND 0.00fF
C2029 a_59666_35682.t1 GND 0.02fF $ **FLOATING
C2030 a_59666_35682.n18 GND 0.07fF
C2031 a_59666_35682.n19 GND 0.02fF
C2032 a_59666_35682.n20 GND 0.05fF
C2033 a_59666_35682.n22 GND 0.04fF
C2034 a_59666_35682.n23 GND 0.04fF
C2035 a_59666_35682.n24 GND 0.00fF
C2036 a_59666_35682.n25 GND 0.00fF
C2037 a_59666_35682.t2 GND 0.02fF $ **FLOATING
C2038 a_59666_35682.n26 GND 0.07fF
C2039 a_59666_35682.n27 GND 0.02fF
C2040 a_59666_35682.n28 GND 0.05fF
C2041 a_59666_35682.n30 GND 0.01fF
C2042 a_59666_35682.n31 GND 0.00fF
C2043 a_59666_35682.n32 GND 0.00fF
C2044 a_59666_35682.n33 GND 0.00fF
C2045 a_59666_35682.n34 GND 0.00fF
C2046 a_59666_35682.n35 GND 0.00fF
C2047 a_59666_35682.n36 GND 0.00fF
C2048 a_59666_35682.n38 GND 0.08fF
C2049 a_59666_35682.t3 GND 4.19fF $ **FLOATING
C2050 a_59666_35682.n39 GND 0.61fF
C2051 a_59666_35682.t0 GND 0.26fF $ **FLOATING
C2052 a_59376_35606.n0 GND 0.01fF
C2053 a_59376_35606.n1 GND 0.01fF
C2054 a_59376_35606.n2 GND 0.00fF
C2055 a_59376_35606.n3 GND 0.00fF
C2056 a_59376_35606.n4 GND 0.00fF
C2057 a_59376_35606.n5 GND 0.00fF
C2058 a_59376_35606.n6 GND 0.00fF
C2059 a_59376_35606.n7 GND 0.00fF
C2060 a_59376_35606.n8 GND 0.00fF
C2061 a_59376_35606.n9 GND 0.00fF
C2062 a_59376_35606.t2 GND 0.02fF $ **FLOATING
C2063 a_59376_35606.t1 GND 0.02fF $ **FLOATING
C2064 a_59376_35606.n10 GND 0.05fF
C2065 a_59376_35606.n11 GND 0.00fF
C2066 a_59376_35606.n12 GND 0.00fF
C2067 a_59376_35606.n13 GND 0.02fF
C2068 a_59376_35606.n14 GND 0.04fF
C2069 a_59376_35606.n15 GND 0.12fF
C2070 a_59376_35606.n16 GND 0.01fF
C2071 a_59376_35606.n17 GND 0.12fF
C2072 a_59376_35606.t3 GND 3.87fF $ **FLOATING
C2073 a_59376_35606.n18 GND 0.52fF
C2074 a_59376_35606.t0 GND 0.24fF $ **FLOATING
C2075 a_31776_65246.n0 GND 0.01fF
C2076 a_31776_65246.n1 GND 0.01fF
C2077 a_31776_65246.n2 GND 0.00fF
C2078 a_31776_65246.n3 GND 0.00fF
C2079 a_31776_65246.n4 GND 0.00fF
C2080 a_31776_65246.n5 GND 0.00fF
C2081 a_31776_65246.n6 GND 0.00fF
C2082 a_31776_65246.n7 GND 0.00fF
C2083 a_31776_65246.n8 GND 0.00fF
C2084 a_31776_65246.n9 GND 0.00fF
C2085 a_31776_65246.t0 GND 0.02fF $ **FLOATING
C2086 a_31776_65246.t1 GND 0.02fF $ **FLOATING
C2087 a_31776_65246.n10 GND 0.05fF
C2088 a_31776_65246.n11 GND 0.00fF
C2089 a_31776_65246.n12 GND 0.00fF
C2090 a_31776_65246.n13 GND 0.02fF
C2091 a_31776_65246.n14 GND 0.04fF
C2092 a_31776_65246.n15 GND 0.12fF
C2093 a_31776_65246.n16 GND 0.01fF
C2094 a_31776_65246.n17 GND 0.12fF
C2095 a_31776_65246.t2 GND 3.87fF $ **FLOATING
C2096 a_31776_65246.n18 GND 0.52fF
C2097 a_31776_65246.t3 GND 0.24fF $ **FLOATING
C2098 a_32066_65322.n0 GND 0.00fF
C2099 a_32066_65322.n1 GND 0.00fF
C2100 a_32066_65322.n2 GND 0.01fF
C2101 a_32066_65322.n3 GND 0.01fF
C2102 a_32066_65322.n4 GND 0.00fF
C2103 a_32066_65322.n5 GND 0.00fF
C2104 a_32066_65322.n6 GND 0.00fF
C2105 a_32066_65322.n7 GND 0.00fF
C2106 a_32066_65322.n8 GND 0.00fF
C2107 a_32066_65322.n9 GND 0.00fF
C2108 a_32066_65322.n10 GND 0.09fF
C2109 a_32066_65322.n11 GND 0.00fF
C2110 a_32066_65322.n12 GND 0.01fF
C2111 a_32066_65322.n13 GND 0.01fF
C2112 a_32066_65322.n14 GND 0.01fF
C2113 a_32066_65322.n15 GND 0.00fF
C2114 a_32066_65322.n16 GND 0.00fF
C2115 a_32066_65322.n17 GND 0.00fF
C2116 a_32066_65322.t1 GND 0.02fF $ **FLOATING
C2117 a_32066_65322.n18 GND 0.07fF
C2118 a_32066_65322.n19 GND 0.02fF
C2119 a_32066_65322.n20 GND 0.05fF
C2120 a_32066_65322.n22 GND 0.04fF
C2121 a_32066_65322.n23 GND 0.04fF
C2122 a_32066_65322.n24 GND 0.00fF
C2123 a_32066_65322.n25 GND 0.00fF
C2124 a_32066_65322.t0 GND 0.02fF $ **FLOATING
C2125 a_32066_65322.n26 GND 0.07fF
C2126 a_32066_65322.n27 GND 0.02fF
C2127 a_32066_65322.n28 GND 0.05fF
C2128 a_32066_65322.n30 GND 0.01fF
C2129 a_32066_65322.n31 GND 0.00fF
C2130 a_32066_65322.n32 GND 0.00fF
C2131 a_32066_65322.n33 GND 0.00fF
C2132 a_32066_65322.n34 GND 0.00fF
C2133 a_32066_65322.n35 GND 0.00fF
C2134 a_32066_65322.n36 GND 0.00fF
C2135 a_32066_65322.n38 GND 0.08fF
C2136 a_32066_65322.t2 GND 4.19fF $ **FLOATING
C2137 a_32066_65322.n39 GND 0.61fF
C2138 a_32066_65322.t3 GND 0.26fF $ **FLOATING
C2139 bit3.t16 GND 0.03fF $ **FLOATING
C2140 bit3.n0 GND 0.01fF
C2141 bit3.n1 GND 0.00fF
C2142 bit3.t7 GND 0.03fF $ **FLOATING
C2143 bit3.n2 GND 0.01fF
C2144 bit3.n3 GND 0.00fF
C2145 bit3.n4 GND 0.00fF
C2146 bit3.n5 GND 0.00fF
C2147 bit3.n6 GND 0.07fF
C2148 bit3.t15 GND 0.03fF $ **FLOATING
C2149 bit3.n7 GND 0.01fF
C2150 bit3.n8 GND 0.00fF
C2151 bit3.t8 GND 0.03fF $ **FLOATING
C2152 bit3.n9 GND 0.01fF
C2153 bit3.n10 GND 0.00fF
C2154 bit3.n11 GND 0.00fF
C2155 bit3.n12 GND 0.00fF
C2156 bit3.n13 GND 0.07fF
C2157 bit3.t5 GND 0.03fF $ **FLOATING
C2158 bit3.n14 GND 0.01fF
C2159 bit3.n15 GND 0.00fF
C2160 bit3.t13 GND 0.03fF $ **FLOATING
C2161 bit3.n16 GND 0.01fF
C2162 bit3.n17 GND 0.00fF
C2163 bit3.n18 GND 0.00fF
C2164 bit3.n19 GND 0.00fF
C2165 bit3.n20 GND 0.07fF
C2166 bit3.t3 GND 0.03fF $ **FLOATING
C2167 bit3.n21 GND 0.01fF
C2168 bit3.n22 GND 0.00fF
C2169 bit3.t12 GND 0.03fF $ **FLOATING
C2170 bit3.n23 GND 0.01fF
C2171 bit3.n24 GND 0.00fF
C2172 bit3.n25 GND 0.00fF
C2173 bit3.n26 GND 0.00fF
C2174 bit3.n27 GND 0.07fF
C2175 bit3.t1 GND 0.03fF $ **FLOATING
C2176 bit3.n28 GND 0.01fF
C2177 bit3.n29 GND 0.00fF
C2178 bit3.t10 GND 0.03fF $ **FLOATING
C2179 bit3.n30 GND 0.01fF
C2180 bit3.n31 GND 0.00fF
C2181 bit3.n32 GND 0.00fF
C2182 bit3.n33 GND 0.00fF
C2183 bit3.n34 GND 0.07fF
C2184 bit3.t4 GND 0.03fF $ **FLOATING
C2185 bit3.n35 GND 0.01fF
C2186 bit3.n36 GND 0.00fF
C2187 bit3.t9 GND 0.03fF $ **FLOATING
C2188 bit3.n37 GND 0.01fF
C2189 bit3.n38 GND 0.00fF
C2190 bit3.n39 GND 0.00fF
C2191 bit3.n40 GND 0.00fF
C2192 bit3.n41 GND 0.07fF
C2193 bit3.t2 GND 0.03fF $ **FLOATING
C2194 bit3.n42 GND 0.01fF
C2195 bit3.n43 GND 0.00fF
C2196 bit3.t11 GND 0.03fF $ **FLOATING
C2197 bit3.n44 GND 0.01fF
C2198 bit3.n45 GND 0.00fF
C2199 bit3.n46 GND 0.00fF
C2200 bit3.n47 GND 0.00fF
C2201 bit3.n48 GND 0.07fF
C2202 bit3.n49 GND 0.00fF
C2203 bit3.n50 GND 0.00fF
C2204 bit3.t6 GND 0.03fF $ **FLOATING
C2205 bit3.n51 GND 0.01fF
C2206 bit3.n52 GND 0.00fF
C2207 bit3.t17 GND 0.03fF $ **FLOATING
C2208 bit3.n53 GND 0.01fF
C2209 bit3.n54 GND 0.00fF
C2210 bit3.n55 GND 0.07fF
C2211 bit3.t14 GND 0.01fF $ **FLOATING
C2212 bit3.t0 GND 0.01fF $ **FLOATING
C2213 bit3.n56 GND 0.03fF
C2214 bit3.n57 GND 18.62fF
C2215 bit3.n58 GND 18.27fF
C2216 bit3.n59 GND 18.27fF
C2217 bit3.n60 GND 18.27fF
C2218 bit3.n61 GND 18.27fF
C2219 bit3.n62 GND 18.27fF
C2220 bit3.n63 GND 18.27fF
C2221 bit3.n64 GND 22.65fF
C2222 a_32066_15922.n0 GND 0.00fF
C2223 a_32066_15922.n1 GND 0.00fF
C2224 a_32066_15922.n2 GND 0.01fF
C2225 a_32066_15922.n3 GND 0.01fF
C2226 a_32066_15922.n4 GND 0.00fF
C2227 a_32066_15922.n5 GND 0.00fF
C2228 a_32066_15922.n6 GND 0.00fF
C2229 a_32066_15922.n7 GND 0.00fF
C2230 a_32066_15922.n8 GND 0.00fF
C2231 a_32066_15922.n9 GND 0.00fF
C2232 a_32066_15922.n10 GND 0.09fF
C2233 a_32066_15922.n11 GND 0.00fF
C2234 a_32066_15922.n12 GND 0.01fF
C2235 a_32066_15922.n13 GND 0.01fF
C2236 a_32066_15922.n14 GND 0.01fF
C2237 a_32066_15922.n15 GND 0.00fF
C2238 a_32066_15922.n16 GND 0.00fF
C2239 a_32066_15922.n17 GND 0.00fF
C2240 a_32066_15922.t2 GND 0.02fF $ **FLOATING
C2241 a_32066_15922.n18 GND 0.07fF
C2242 a_32066_15922.n19 GND 0.02fF
C2243 a_32066_15922.n20 GND 0.05fF
C2244 a_32066_15922.n22 GND 0.04fF
C2245 a_32066_15922.n23 GND 0.04fF
C2246 a_32066_15922.n24 GND 0.00fF
C2247 a_32066_15922.n25 GND 0.00fF
C2248 a_32066_15922.t1 GND 0.02fF $ **FLOATING
C2249 a_32066_15922.n26 GND 0.07fF
C2250 a_32066_15922.n27 GND 0.02fF
C2251 a_32066_15922.n28 GND 0.05fF
C2252 a_32066_15922.n30 GND 0.01fF
C2253 a_32066_15922.n31 GND 0.00fF
C2254 a_32066_15922.n32 GND 0.00fF
C2255 a_32066_15922.n33 GND 0.00fF
C2256 a_32066_15922.n34 GND 0.00fF
C2257 a_32066_15922.n35 GND 0.00fF
C2258 a_32066_15922.n36 GND 0.00fF
C2259 a_32066_15922.n38 GND 0.08fF
C2260 a_32066_15922.t3 GND 4.19fF $ **FLOATING
C2261 a_32066_15922.n39 GND 0.61fF
C2262 a_32066_15922.t0 GND 0.26fF $ **FLOATING
C2263 a_41266_25802.n0 GND 0.00fF
C2264 a_41266_25802.n1 GND 0.00fF
C2265 a_41266_25802.n2 GND 0.01fF
C2266 a_41266_25802.n3 GND 0.01fF
C2267 a_41266_25802.n4 GND 0.00fF
C2268 a_41266_25802.n5 GND 0.00fF
C2269 a_41266_25802.n6 GND 0.00fF
C2270 a_41266_25802.n7 GND 0.00fF
C2271 a_41266_25802.n8 GND 0.00fF
C2272 a_41266_25802.n9 GND 0.00fF
C2273 a_41266_25802.n10 GND 0.09fF
C2274 a_41266_25802.n11 GND 0.00fF
C2275 a_41266_25802.n12 GND 0.01fF
C2276 a_41266_25802.n13 GND 0.01fF
C2277 a_41266_25802.n14 GND 0.01fF
C2278 a_41266_25802.n15 GND 0.00fF
C2279 a_41266_25802.n16 GND 0.00fF
C2280 a_41266_25802.n17 GND 0.00fF
C2281 a_41266_25802.t0 GND 0.02fF $ **FLOATING
C2282 a_41266_25802.n18 GND 0.07fF
C2283 a_41266_25802.n19 GND 0.02fF
C2284 a_41266_25802.n20 GND 0.05fF
C2285 a_41266_25802.n22 GND 0.04fF
C2286 a_41266_25802.n23 GND 0.04fF
C2287 a_41266_25802.n24 GND 0.00fF
C2288 a_41266_25802.n25 GND 0.00fF
C2289 a_41266_25802.t1 GND 0.02fF $ **FLOATING
C2290 a_41266_25802.n26 GND 0.07fF
C2291 a_41266_25802.n27 GND 0.02fF
C2292 a_41266_25802.n28 GND 0.05fF
C2293 a_41266_25802.n30 GND 0.01fF
C2294 a_41266_25802.n31 GND 0.00fF
C2295 a_41266_25802.n32 GND 0.00fF
C2296 a_41266_25802.n33 GND 0.00fF
C2297 a_41266_25802.n34 GND 0.00fF
C2298 a_41266_25802.n35 GND 0.00fF
C2299 a_41266_25802.n36 GND 0.00fF
C2300 a_41266_25802.n38 GND 0.08fF
C2301 a_41266_25802.t3 GND 4.19fF $ **FLOATING
C2302 a_41266_25802.n39 GND 0.61fF
C2303 a_41266_25802.t2 GND 0.26fF $ **FLOATING
C2304 a_50466_55442.n0 GND 0.00fF
C2305 a_50466_55442.n1 GND 0.00fF
C2306 a_50466_55442.n2 GND 0.01fF
C2307 a_50466_55442.n3 GND 0.01fF
C2308 a_50466_55442.n4 GND 0.00fF
C2309 a_50466_55442.n5 GND 0.00fF
C2310 a_50466_55442.n6 GND 0.00fF
C2311 a_50466_55442.n7 GND 0.00fF
C2312 a_50466_55442.n8 GND 0.00fF
C2313 a_50466_55442.n9 GND 0.00fF
C2314 a_50466_55442.n10 GND 0.09fF
C2315 a_50466_55442.n11 GND 0.00fF
C2316 a_50466_55442.n12 GND 0.01fF
C2317 a_50466_55442.n13 GND 0.01fF
C2318 a_50466_55442.n14 GND 0.01fF
C2319 a_50466_55442.n15 GND 0.00fF
C2320 a_50466_55442.n16 GND 0.00fF
C2321 a_50466_55442.n17 GND 0.00fF
C2322 a_50466_55442.t1 GND 0.02fF $ **FLOATING
C2323 a_50466_55442.n18 GND 0.07fF
C2324 a_50466_55442.n19 GND 0.02fF
C2325 a_50466_55442.n20 GND 0.05fF
C2326 a_50466_55442.n22 GND 0.04fF
C2327 a_50466_55442.n23 GND 0.04fF
C2328 a_50466_55442.n24 GND 0.00fF
C2329 a_50466_55442.n25 GND 0.00fF
C2330 a_50466_55442.t0 GND 0.02fF $ **FLOATING
C2331 a_50466_55442.n26 GND 0.07fF
C2332 a_50466_55442.n27 GND 0.02fF
C2333 a_50466_55442.n28 GND 0.05fF
C2334 a_50466_55442.n30 GND 0.01fF
C2335 a_50466_55442.n31 GND 0.00fF
C2336 a_50466_55442.n32 GND 0.00fF
C2337 a_50466_55442.n33 GND 0.00fF
C2338 a_50466_55442.n34 GND 0.00fF
C2339 a_50466_55442.n35 GND 0.00fF
C2340 a_50466_55442.n36 GND 0.00fF
C2341 a_50466_55442.n38 GND 0.08fF
C2342 a_50466_55442.t2 GND 4.19fF $ **FLOATING
C2343 a_50466_55442.n39 GND 0.61fF
C2344 a_50466_55442.t3 GND 0.26fF $ **FLOATING
C2345 a_68866_6042.n0 GND 0.00fF
C2346 a_68866_6042.n1 GND 0.00fF
C2347 a_68866_6042.n2 GND 0.01fF
C2348 a_68866_6042.n3 GND 0.01fF
C2349 a_68866_6042.n4 GND 0.00fF
C2350 a_68866_6042.n5 GND 0.00fF
C2351 a_68866_6042.n6 GND 0.00fF
C2352 a_68866_6042.n7 GND 0.00fF
C2353 a_68866_6042.n8 GND 0.00fF
C2354 a_68866_6042.n9 GND 0.00fF
C2355 a_68866_6042.n10 GND 0.09fF
C2356 a_68866_6042.n11 GND 0.00fF
C2357 a_68866_6042.n12 GND 0.01fF
C2358 a_68866_6042.n13 GND 0.01fF
C2359 a_68866_6042.n14 GND 0.01fF
C2360 a_68866_6042.n15 GND 0.00fF
C2361 a_68866_6042.n16 GND 0.00fF
C2362 a_68866_6042.n17 GND 0.00fF
C2363 a_68866_6042.t2 GND 0.02fF $ **FLOATING
C2364 a_68866_6042.n18 GND 0.07fF
C2365 a_68866_6042.n19 GND 0.02fF
C2366 a_68866_6042.n20 GND 0.05fF
C2367 a_68866_6042.n22 GND 0.04fF
C2368 a_68866_6042.n23 GND 0.04fF
C2369 a_68866_6042.n24 GND 0.00fF
C2370 a_68866_6042.n25 GND 0.00fF
C2371 a_68866_6042.t1 GND 0.02fF $ **FLOATING
C2372 a_68866_6042.n26 GND 0.07fF
C2373 a_68866_6042.n27 GND 0.02fF
C2374 a_68866_6042.n28 GND 0.05fF
C2375 a_68866_6042.n30 GND 0.01fF
C2376 a_68866_6042.n31 GND 0.00fF
C2377 a_68866_6042.n32 GND 0.00fF
C2378 a_68866_6042.n33 GND 0.00fF
C2379 a_68866_6042.n34 GND 0.00fF
C2380 a_68866_6042.n35 GND 0.00fF
C2381 a_68866_6042.n36 GND 0.00fF
C2382 a_68866_6042.n38 GND 0.08fF
C2383 a_68866_6042.t3 GND 4.19fF $ **FLOATING
C2384 a_68866_6042.n39 GND 0.61fF
C2385 a_68866_6042.t0 GND 0.26fF $ **FLOATING
C2386 a_31776_35606.n0 GND 0.01fF
C2387 a_31776_35606.n1 GND 0.01fF
C2388 a_31776_35606.n2 GND 0.00fF
C2389 a_31776_35606.n3 GND 0.00fF
C2390 a_31776_35606.n4 GND 0.00fF
C2391 a_31776_35606.n5 GND 0.00fF
C2392 a_31776_35606.n6 GND 0.00fF
C2393 a_31776_35606.n7 GND 0.00fF
C2394 a_31776_35606.n8 GND 0.00fF
C2395 a_31776_35606.n9 GND 0.00fF
C2396 a_31776_35606.t1 GND 0.02fF $ **FLOATING
C2397 a_31776_35606.t0 GND 0.02fF $ **FLOATING
C2398 a_31776_35606.n10 GND 0.05fF
C2399 a_31776_35606.n11 GND 0.00fF
C2400 a_31776_35606.n12 GND 0.00fF
C2401 a_31776_35606.n13 GND 0.02fF
C2402 a_31776_35606.n14 GND 0.04fF
C2403 a_31776_35606.n15 GND 0.12fF
C2404 a_31776_35606.n16 GND 0.01fF
C2405 a_31776_35606.n17 GND 0.12fF
C2406 a_31776_35606.t2 GND 3.87fF $ **FLOATING
C2407 a_31776_35606.n18 GND 0.52fF
C2408 a_31776_35606.t3 GND 0.24fF $ **FLOATING
C2409 a_4176_25726.n0 GND 0.01fF
C2410 a_4176_25726.n1 GND 0.01fF
C2411 a_4176_25726.n2 GND 0.00fF
C2412 a_4176_25726.n3 GND 0.00fF
C2413 a_4176_25726.n4 GND 0.00fF
C2414 a_4176_25726.n5 GND 0.00fF
C2415 a_4176_25726.n6 GND 0.00fF
C2416 a_4176_25726.n7 GND 0.00fF
C2417 a_4176_25726.n8 GND 0.00fF
C2418 a_4176_25726.n9 GND 0.00fF
C2419 a_4176_25726.t0 GND 0.02fF $ **FLOATING
C2420 a_4176_25726.t1 GND 0.02fF $ **FLOATING
C2421 a_4176_25726.n10 GND 0.05fF
C2422 a_4176_25726.n11 GND 0.00fF
C2423 a_4176_25726.n12 GND 0.00fF
C2424 a_4176_25726.n13 GND 0.02fF
C2425 a_4176_25726.n14 GND 0.04fF
C2426 a_4176_25726.n15 GND 0.12fF
C2427 a_4176_25726.n16 GND 0.01fF
C2428 a_4176_25726.n17 GND 0.12fF
C2429 a_4176_25726.t2 GND 3.87fF $ **FLOATING
C2430 a_4176_25726.n18 GND 0.52fF
C2431 a_4176_25726.t3 GND 0.24fF $ **FLOATING
C2432 a_13666_25802.n0 GND 0.00fF
C2433 a_13666_25802.n1 GND 0.00fF
C2434 a_13666_25802.n2 GND 0.01fF
C2435 a_13666_25802.n3 GND 0.01fF
C2436 a_13666_25802.n4 GND 0.00fF
C2437 a_13666_25802.n5 GND 0.00fF
C2438 a_13666_25802.n6 GND 0.00fF
C2439 a_13666_25802.n7 GND 0.00fF
C2440 a_13666_25802.n8 GND 0.00fF
C2441 a_13666_25802.n9 GND 0.00fF
C2442 a_13666_25802.n10 GND 0.09fF
C2443 a_13666_25802.n11 GND 0.00fF
C2444 a_13666_25802.n12 GND 0.01fF
C2445 a_13666_25802.n13 GND 0.01fF
C2446 a_13666_25802.n14 GND 0.01fF
C2447 a_13666_25802.n15 GND 0.00fF
C2448 a_13666_25802.n16 GND 0.00fF
C2449 a_13666_25802.n17 GND 0.00fF
C2450 a_13666_25802.t0 GND 0.02fF $ **FLOATING
C2451 a_13666_25802.n18 GND 0.07fF
C2452 a_13666_25802.n19 GND 0.02fF
C2453 a_13666_25802.n20 GND 0.05fF
C2454 a_13666_25802.n22 GND 0.04fF
C2455 a_13666_25802.n23 GND 0.04fF
C2456 a_13666_25802.n24 GND 0.00fF
C2457 a_13666_25802.n25 GND 0.00fF
C2458 a_13666_25802.t1 GND 0.02fF $ **FLOATING
C2459 a_13666_25802.n26 GND 0.07fF
C2460 a_13666_25802.n27 GND 0.02fF
C2461 a_13666_25802.n28 GND 0.05fF
C2462 a_13666_25802.n30 GND 0.01fF
C2463 a_13666_25802.n31 GND 0.00fF
C2464 a_13666_25802.n32 GND 0.00fF
C2465 a_13666_25802.n33 GND 0.00fF
C2466 a_13666_25802.n34 GND 0.00fF
C2467 a_13666_25802.n35 GND 0.00fF
C2468 a_13666_25802.n36 GND 0.00fF
C2469 a_13666_25802.n38 GND 0.08fF
C2470 a_13666_25802.t2 GND 4.19fF $ **FLOATING
C2471 a_13666_25802.n39 GND 0.61fF
C2472 a_13666_25802.t3 GND 0.26fF $ **FLOATING
C2473 a_13376_25726.n0 GND 0.01fF
C2474 a_13376_25726.n1 GND 0.01fF
C2475 a_13376_25726.n2 GND 0.00fF
C2476 a_13376_25726.n3 GND 0.00fF
C2477 a_13376_25726.n4 GND 0.00fF
C2478 a_13376_25726.n5 GND 0.00fF
C2479 a_13376_25726.n6 GND 0.00fF
C2480 a_13376_25726.n7 GND 0.00fF
C2481 a_13376_25726.n8 GND 0.00fF
C2482 a_13376_25726.n9 GND 0.00fF
C2483 a_13376_25726.t1 GND 0.02fF $ **FLOATING
C2484 a_13376_25726.t0 GND 0.02fF $ **FLOATING
C2485 a_13376_25726.n10 GND 0.05fF
C2486 a_13376_25726.n11 GND 0.00fF
C2487 a_13376_25726.n12 GND 0.00fF
C2488 a_13376_25726.n13 GND 0.02fF
C2489 a_13376_25726.n14 GND 0.04fF
C2490 a_13376_25726.n15 GND 0.12fF
C2491 a_13376_25726.n16 GND 0.01fF
C2492 a_13376_25726.n17 GND 0.12fF
C2493 a_13376_25726.t2 GND 3.87fF $ **FLOATING
C2494 a_13376_25726.n18 GND 0.52fF
C2495 a_13376_25726.t3 GND 0.24fF $ **FLOATING
C2496 a_59376_55366.n0 GND 0.01fF
C2497 a_59376_55366.n1 GND 0.01fF
C2498 a_59376_55366.n2 GND 0.00fF
C2499 a_59376_55366.n3 GND 0.00fF
C2500 a_59376_55366.n4 GND 0.00fF
C2501 a_59376_55366.n5 GND 0.00fF
C2502 a_59376_55366.n6 GND 0.00fF
C2503 a_59376_55366.n7 GND 0.00fF
C2504 a_59376_55366.n8 GND 0.00fF
C2505 a_59376_55366.n9 GND 0.00fF
C2506 a_59376_55366.t1 GND 0.02fF $ **FLOATING
C2507 a_59376_55366.t0 GND 0.02fF $ **FLOATING
C2508 a_59376_55366.n10 GND 0.05fF
C2509 a_59376_55366.n11 GND 0.00fF
C2510 a_59376_55366.n12 GND 0.00fF
C2511 a_59376_55366.n13 GND 0.02fF
C2512 a_59376_55366.n14 GND 0.04fF
C2513 a_59376_55366.n15 GND 0.12fF
C2514 a_59376_55366.n16 GND 0.01fF
C2515 a_59376_55366.n17 GND 0.12fF
C2516 a_59376_55366.t2 GND 3.87fF $ **FLOATING
C2517 a_59376_55366.n18 GND 0.52fF
C2518 a_59376_55366.t3 GND 0.24fF $ **FLOATING
C2519 a_59376_15846.n0 GND 0.01fF
C2520 a_59376_15846.n1 GND 0.01fF
C2521 a_59376_15846.n2 GND 0.00fF
C2522 a_59376_15846.n3 GND 0.00fF
C2523 a_59376_15846.n4 GND 0.00fF
C2524 a_59376_15846.n5 GND 0.00fF
C2525 a_59376_15846.n6 GND 0.00fF
C2526 a_59376_15846.n7 GND 0.00fF
C2527 a_59376_15846.n8 GND 0.00fF
C2528 a_59376_15846.n9 GND 0.00fF
C2529 a_59376_15846.t0 GND 0.02fF $ **FLOATING
C2530 a_59376_15846.t1 GND 0.02fF $ **FLOATING
C2531 a_59376_15846.n10 GND 0.05fF
C2532 a_59376_15846.n11 GND 0.00fF
C2533 a_59376_15846.n12 GND 0.00fF
C2534 a_59376_15846.n13 GND 0.02fF
C2535 a_59376_15846.n14 GND 0.04fF
C2536 a_59376_15846.n15 GND 0.12fF
C2537 a_59376_15846.n16 GND 0.01fF
C2538 a_59376_15846.n17 GND 0.12fF
C2539 a_59376_15846.t3 GND 3.87fF $ **FLOATING
C2540 a_59376_15846.n18 GND 0.52fF
C2541 a_59376_15846.t2 GND 0.24fF $ **FLOATING
C2542 a_59666_15922.n0 GND 0.00fF
C2543 a_59666_15922.n1 GND 0.00fF
C2544 a_59666_15922.n2 GND 0.01fF
C2545 a_59666_15922.n3 GND 0.01fF
C2546 a_59666_15922.n4 GND 0.00fF
C2547 a_59666_15922.n5 GND 0.00fF
C2548 a_59666_15922.n6 GND 0.00fF
C2549 a_59666_15922.n7 GND 0.00fF
C2550 a_59666_15922.n8 GND 0.00fF
C2551 a_59666_15922.n9 GND 0.00fF
C2552 a_59666_15922.n10 GND 0.09fF
C2553 a_59666_15922.n11 GND 0.00fF
C2554 a_59666_15922.n12 GND 0.01fF
C2555 a_59666_15922.n13 GND 0.01fF
C2556 a_59666_15922.n14 GND 0.01fF
C2557 a_59666_15922.n15 GND 0.00fF
C2558 a_59666_15922.n16 GND 0.00fF
C2559 a_59666_15922.n17 GND 0.00fF
C2560 a_59666_15922.t2 GND 0.02fF $ **FLOATING
C2561 a_59666_15922.n18 GND 0.07fF
C2562 a_59666_15922.n19 GND 0.02fF
C2563 a_59666_15922.n20 GND 0.05fF
C2564 a_59666_15922.n22 GND 0.04fF
C2565 a_59666_15922.n23 GND 0.04fF
C2566 a_59666_15922.n24 GND 0.00fF
C2567 a_59666_15922.n25 GND 0.00fF
C2568 a_59666_15922.t1 GND 0.02fF $ **FLOATING
C2569 a_59666_15922.n26 GND 0.07fF
C2570 a_59666_15922.n27 GND 0.02fF
C2571 a_59666_15922.n28 GND 0.05fF
C2572 a_59666_15922.n30 GND 0.01fF
C2573 a_59666_15922.n31 GND 0.00fF
C2574 a_59666_15922.n32 GND 0.00fF
C2575 a_59666_15922.n33 GND 0.00fF
C2576 a_59666_15922.n34 GND 0.00fF
C2577 a_59666_15922.n35 GND 0.00fF
C2578 a_59666_15922.n36 GND 0.00fF
C2579 a_59666_15922.n38 GND 0.08fF
C2580 a_59666_15922.t3 GND 4.19fF $ **FLOATING
C2581 a_59666_15922.n39 GND 0.61fF
C2582 a_59666_15922.t0 GND 0.26fF $ **FLOATING
C2583 a_50176_35606.n0 GND 0.01fF
C2584 a_50176_35606.n1 GND 0.01fF
C2585 a_50176_35606.n2 GND 0.00fF
C2586 a_50176_35606.n3 GND 0.00fF
C2587 a_50176_35606.n4 GND 0.00fF
C2588 a_50176_35606.n5 GND 0.00fF
C2589 a_50176_35606.n6 GND 0.00fF
C2590 a_50176_35606.n7 GND 0.00fF
C2591 a_50176_35606.n8 GND 0.00fF
C2592 a_50176_35606.n9 GND 0.00fF
C2593 a_50176_35606.t1 GND 0.02fF $ **FLOATING
C2594 a_50176_35606.t0 GND 0.02fF $ **FLOATING
C2595 a_50176_35606.n10 GND 0.05fF
C2596 a_50176_35606.n11 GND 0.00fF
C2597 a_50176_35606.n12 GND 0.00fF
C2598 a_50176_35606.n13 GND 0.02fF
C2599 a_50176_35606.n14 GND 0.04fF
C2600 a_50176_35606.n15 GND 0.12fF
C2601 a_50176_35606.n16 GND 0.01fF
C2602 a_50176_35606.n17 GND 0.12fF
C2603 a_50176_35606.t2 GND 3.87fF $ **FLOATING
C2604 a_50176_35606.n18 GND 0.52fF
C2605 a_50176_35606.t3 GND 0.24fF $ **FLOATING
C2606 a_32066_25802.n0 GND 0.00fF
C2607 a_32066_25802.n1 GND 0.00fF
C2608 a_32066_25802.n2 GND 0.01fF
C2609 a_32066_25802.n3 GND 0.01fF
C2610 a_32066_25802.n4 GND 0.00fF
C2611 a_32066_25802.n5 GND 0.00fF
C2612 a_32066_25802.n6 GND 0.00fF
C2613 a_32066_25802.n7 GND 0.00fF
C2614 a_32066_25802.n8 GND 0.00fF
C2615 a_32066_25802.n9 GND 0.00fF
C2616 a_32066_25802.n10 GND 0.09fF
C2617 a_32066_25802.n11 GND 0.00fF
C2618 a_32066_25802.n12 GND 0.01fF
C2619 a_32066_25802.n13 GND 0.01fF
C2620 a_32066_25802.n14 GND 0.01fF
C2621 a_32066_25802.n15 GND 0.00fF
C2622 a_32066_25802.n16 GND 0.00fF
C2623 a_32066_25802.n17 GND 0.00fF
C2624 a_32066_25802.t0 GND 0.02fF $ **FLOATING
C2625 a_32066_25802.n18 GND 0.07fF
C2626 a_32066_25802.n19 GND 0.02fF
C2627 a_32066_25802.n20 GND 0.05fF
C2628 a_32066_25802.n22 GND 0.04fF
C2629 a_32066_25802.n23 GND 0.04fF
C2630 a_32066_25802.n24 GND 0.00fF
C2631 a_32066_25802.n25 GND 0.00fF
C2632 a_32066_25802.t1 GND 0.02fF $ **FLOATING
C2633 a_32066_25802.n26 GND 0.07fF
C2634 a_32066_25802.n27 GND 0.02fF
C2635 a_32066_25802.n28 GND 0.05fF
C2636 a_32066_25802.n30 GND 0.01fF
C2637 a_32066_25802.n31 GND 0.00fF
C2638 a_32066_25802.n32 GND 0.00fF
C2639 a_32066_25802.n33 GND 0.00fF
C2640 a_32066_25802.n34 GND 0.00fF
C2641 a_32066_25802.n35 GND 0.00fF
C2642 a_32066_25802.n36 GND 0.00fF
C2643 a_32066_25802.n38 GND 0.08fF
C2644 a_32066_25802.t2 GND 4.19fF $ **FLOATING
C2645 a_32066_25802.n39 GND 0.61fF
C2646 a_32066_25802.t3 GND 0.26fF $ **FLOATING
C2647 a_22866_15922.n0 GND 0.00fF
C2648 a_22866_15922.n1 GND 0.00fF
C2649 a_22866_15922.n2 GND 0.01fF
C2650 a_22866_15922.n3 GND 0.01fF
C2651 a_22866_15922.n4 GND 0.00fF
C2652 a_22866_15922.n5 GND 0.00fF
C2653 a_22866_15922.n6 GND 0.00fF
C2654 a_22866_15922.n7 GND 0.00fF
C2655 a_22866_15922.n8 GND 0.00fF
C2656 a_22866_15922.n9 GND 0.00fF
C2657 a_22866_15922.n10 GND 0.09fF
C2658 a_22866_15922.n11 GND 0.00fF
C2659 a_22866_15922.n12 GND 0.01fF
C2660 a_22866_15922.n13 GND 0.01fF
C2661 a_22866_15922.n14 GND 0.01fF
C2662 a_22866_15922.n15 GND 0.00fF
C2663 a_22866_15922.n16 GND 0.00fF
C2664 a_22866_15922.n17 GND 0.00fF
C2665 a_22866_15922.t1 GND 0.02fF $ **FLOATING
C2666 a_22866_15922.n18 GND 0.07fF
C2667 a_22866_15922.n19 GND 0.02fF
C2668 a_22866_15922.n20 GND 0.05fF
C2669 a_22866_15922.n22 GND 0.04fF
C2670 a_22866_15922.n23 GND 0.04fF
C2671 a_22866_15922.n24 GND 0.00fF
C2672 a_22866_15922.n25 GND 0.00fF
C2673 a_22866_15922.t0 GND 0.02fF $ **FLOATING
C2674 a_22866_15922.n26 GND 0.07fF
C2675 a_22866_15922.n27 GND 0.02fF
C2676 a_22866_15922.n28 GND 0.05fF
C2677 a_22866_15922.n30 GND 0.01fF
C2678 a_22866_15922.n31 GND 0.00fF
C2679 a_22866_15922.n32 GND 0.00fF
C2680 a_22866_15922.n33 GND 0.00fF
C2681 a_22866_15922.n34 GND 0.00fF
C2682 a_22866_15922.n35 GND 0.00fF
C2683 a_22866_15922.n36 GND 0.00fF
C2684 a_22866_15922.n38 GND 0.08fF
C2685 a_22866_15922.t3 GND 4.19fF $ **FLOATING
C2686 a_22866_15922.n39 GND 0.61fF
C2687 a_22866_15922.t2 GND 0.26fF $ **FLOATING
C2688 a_13666_65322.n0 GND 0.00fF
C2689 a_13666_65322.n1 GND 0.00fF
C2690 a_13666_65322.n2 GND 0.01fF
C2691 a_13666_65322.n3 GND 0.01fF
C2692 a_13666_65322.n4 GND 0.00fF
C2693 a_13666_65322.n5 GND 0.00fF
C2694 a_13666_65322.n6 GND 0.00fF
C2695 a_13666_65322.n7 GND 0.00fF
C2696 a_13666_65322.n8 GND 0.00fF
C2697 a_13666_65322.n9 GND 0.00fF
C2698 a_13666_65322.n10 GND 0.09fF
C2699 a_13666_65322.n11 GND 0.00fF
C2700 a_13666_65322.n12 GND 0.01fF
C2701 a_13666_65322.n13 GND 0.01fF
C2702 a_13666_65322.n14 GND 0.01fF
C2703 a_13666_65322.n15 GND 0.00fF
C2704 a_13666_65322.n16 GND 0.00fF
C2705 a_13666_65322.n17 GND 0.00fF
C2706 a_13666_65322.t3 GND 0.02fF $ **FLOATING
C2707 a_13666_65322.n18 GND 0.07fF
C2708 a_13666_65322.n19 GND 0.02fF
C2709 a_13666_65322.n20 GND 0.05fF
C2710 a_13666_65322.n22 GND 0.04fF
C2711 a_13666_65322.n23 GND 0.04fF
C2712 a_13666_65322.n24 GND 0.00fF
C2713 a_13666_65322.n25 GND 0.00fF
C2714 a_13666_65322.t0 GND 0.02fF $ **FLOATING
C2715 a_13666_65322.n26 GND 0.07fF
C2716 a_13666_65322.n27 GND 0.02fF
C2717 a_13666_65322.n28 GND 0.05fF
C2718 a_13666_65322.n30 GND 0.01fF
C2719 a_13666_65322.n31 GND 0.00fF
C2720 a_13666_65322.n32 GND 0.00fF
C2721 a_13666_65322.n33 GND 0.00fF
C2722 a_13666_65322.n34 GND 0.00fF
C2723 a_13666_65322.n35 GND 0.00fF
C2724 a_13666_65322.n36 GND 0.00fF
C2725 a_13666_65322.n38 GND 0.08fF
C2726 a_13666_65322.t2 GND 4.19fF $ **FLOATING
C2727 a_13666_65322.n39 GND 0.61fF
C2728 a_13666_65322.t1 GND 0.26fF $ **FLOATING
C2729 a_22866_6042.n0 GND 0.00fF
C2730 a_22866_6042.n1 GND 0.00fF
C2731 a_22866_6042.n2 GND 0.01fF
C2732 a_22866_6042.n3 GND 0.01fF
C2733 a_22866_6042.n4 GND 0.00fF
C2734 a_22866_6042.n5 GND 0.00fF
C2735 a_22866_6042.n6 GND 0.00fF
C2736 a_22866_6042.n7 GND 0.00fF
C2737 a_22866_6042.n8 GND 0.00fF
C2738 a_22866_6042.n9 GND 0.00fF
C2739 a_22866_6042.n10 GND 0.09fF
C2740 a_22866_6042.n11 GND 0.00fF
C2741 a_22866_6042.n12 GND 0.01fF
C2742 a_22866_6042.n13 GND 0.01fF
C2743 a_22866_6042.n14 GND 0.01fF
C2744 a_22866_6042.n15 GND 0.00fF
C2745 a_22866_6042.n16 GND 0.00fF
C2746 a_22866_6042.n17 GND 0.00fF
C2747 a_22866_6042.t0 GND 0.02fF $ **FLOATING
C2748 a_22866_6042.n18 GND 0.07fF
C2749 a_22866_6042.n19 GND 0.02fF
C2750 a_22866_6042.n20 GND 0.05fF
C2751 a_22866_6042.n22 GND 0.04fF
C2752 a_22866_6042.n23 GND 0.04fF
C2753 a_22866_6042.n24 GND 0.00fF
C2754 a_22866_6042.n25 GND 0.00fF
C2755 a_22866_6042.t1 GND 0.02fF $ **FLOATING
C2756 a_22866_6042.n26 GND 0.07fF
C2757 a_22866_6042.n27 GND 0.02fF
C2758 a_22866_6042.n28 GND 0.05fF
C2759 a_22866_6042.n30 GND 0.01fF
C2760 a_22866_6042.n31 GND 0.00fF
C2761 a_22866_6042.n32 GND 0.00fF
C2762 a_22866_6042.n33 GND 0.00fF
C2763 a_22866_6042.n34 GND 0.00fF
C2764 a_22866_6042.n35 GND 0.00fF
C2765 a_22866_6042.n36 GND 0.00fF
C2766 a_22866_6042.n38 GND 0.08fF
C2767 a_22866_6042.t3 GND 4.19fF $ **FLOATING
C2768 a_22866_6042.n39 GND 0.61fF
C2769 a_22866_6042.t2 GND 0.26fF $ **FLOATING
C2770 a_22576_5966.n0 GND 0.01fF
C2771 a_22576_5966.n1 GND 0.01fF
C2772 a_22576_5966.n2 GND 0.00fF
C2773 a_22576_5966.n3 GND 0.00fF
C2774 a_22576_5966.n4 GND 0.00fF
C2775 a_22576_5966.n5 GND 0.00fF
C2776 a_22576_5966.n6 GND 0.00fF
C2777 a_22576_5966.n7 GND 0.00fF
C2778 a_22576_5966.n8 GND 0.00fF
C2779 a_22576_5966.n9 GND 0.00fF
C2780 a_22576_5966.t1 GND 0.02fF $ **FLOATING
C2781 a_22576_5966.t0 GND 0.02fF $ **FLOATING
C2782 a_22576_5966.n10 GND 0.05fF
C2783 a_22576_5966.n11 GND 0.00fF
C2784 a_22576_5966.n12 GND 0.00fF
C2785 a_22576_5966.n13 GND 0.02fF
C2786 a_22576_5966.n14 GND 0.04fF
C2787 a_22576_5966.n15 GND 0.12fF
C2788 a_22576_5966.n16 GND 0.01fF
C2789 a_22576_5966.n17 GND 0.12fF
C2790 a_22576_5966.t2 GND 3.87fF $ **FLOATING
C2791 a_22576_5966.n18 GND 0.52fF
C2792 a_22576_5966.t3 GND 0.24fF $ **FLOATING
C2793 a_13376_45486.n0 GND 0.01fF
C2794 a_13376_45486.n1 GND 0.01fF
C2795 a_13376_45486.n2 GND 0.00fF
C2796 a_13376_45486.n3 GND 0.00fF
C2797 a_13376_45486.n4 GND 0.00fF
C2798 a_13376_45486.n5 GND 0.00fF
C2799 a_13376_45486.n6 GND 0.00fF
C2800 a_13376_45486.n7 GND 0.00fF
C2801 a_13376_45486.n8 GND 0.00fF
C2802 a_13376_45486.n9 GND 0.00fF
C2803 a_13376_45486.t1 GND 0.02fF $ **FLOATING
C2804 a_13376_45486.t0 GND 0.02fF $ **FLOATING
C2805 a_13376_45486.n10 GND 0.05fF
C2806 a_13376_45486.n11 GND 0.00fF
C2807 a_13376_45486.n12 GND 0.00fF
C2808 a_13376_45486.n13 GND 0.02fF
C2809 a_13376_45486.n14 GND 0.04fF
C2810 a_13376_45486.n15 GND 0.12fF
C2811 a_13376_45486.n16 GND 0.01fF
C2812 a_13376_45486.n17 GND 0.12fF
C2813 a_13376_45486.t3 GND 3.87fF $ **FLOATING
C2814 a_13376_45486.n18 GND 0.52fF
C2815 a_13376_45486.t2 GND 0.24fF $ **FLOATING
C2816 a_50466_15922.n0 GND 0.00fF
C2817 a_50466_15922.n1 GND 0.00fF
C2818 a_50466_15922.n2 GND 0.01fF
C2819 a_50466_15922.n3 GND 0.01fF
C2820 a_50466_15922.n4 GND 0.00fF
C2821 a_50466_15922.n5 GND 0.00fF
C2822 a_50466_15922.n6 GND 0.00fF
C2823 a_50466_15922.n7 GND 0.00fF
C2824 a_50466_15922.n8 GND 0.00fF
C2825 a_50466_15922.n9 GND 0.00fF
C2826 a_50466_15922.n10 GND 0.09fF
C2827 a_50466_15922.n11 GND 0.00fF
C2828 a_50466_15922.n12 GND 0.01fF
C2829 a_50466_15922.n13 GND 0.01fF
C2830 a_50466_15922.n14 GND 0.01fF
C2831 a_50466_15922.n15 GND 0.00fF
C2832 a_50466_15922.n16 GND 0.00fF
C2833 a_50466_15922.n17 GND 0.00fF
C2834 a_50466_15922.t0 GND 0.02fF $ **FLOATING
C2835 a_50466_15922.n18 GND 0.07fF
C2836 a_50466_15922.n19 GND 0.02fF
C2837 a_50466_15922.n20 GND 0.05fF
C2838 a_50466_15922.n22 GND 0.04fF
C2839 a_50466_15922.n23 GND 0.04fF
C2840 a_50466_15922.n24 GND 0.00fF
C2841 a_50466_15922.n25 GND 0.00fF
C2842 a_50466_15922.t1 GND 0.02fF $ **FLOATING
C2843 a_50466_15922.n26 GND 0.07fF
C2844 a_50466_15922.n27 GND 0.02fF
C2845 a_50466_15922.n28 GND 0.05fF
C2846 a_50466_15922.n30 GND 0.01fF
C2847 a_50466_15922.n31 GND 0.00fF
C2848 a_50466_15922.n32 GND 0.00fF
C2849 a_50466_15922.n33 GND 0.00fF
C2850 a_50466_15922.n34 GND 0.00fF
C2851 a_50466_15922.n35 GND 0.00fF
C2852 a_50466_15922.n36 GND 0.00fF
C2853 a_50466_15922.n38 GND 0.08fF
C2854 a_50466_15922.t2 GND 4.19fF $ **FLOATING
C2855 a_50466_15922.n39 GND 0.61fF
C2856 a_50466_15922.t3 GND 0.26fF $ **FLOATING
C2857 a_50176_15846.n0 GND 0.01fF
C2858 a_50176_15846.n1 GND 0.01fF
C2859 a_50176_15846.n2 GND 0.00fF
C2860 a_50176_15846.n3 GND 0.00fF
C2861 a_50176_15846.n4 GND 0.00fF
C2862 a_50176_15846.n5 GND 0.00fF
C2863 a_50176_15846.n6 GND 0.00fF
C2864 a_50176_15846.n7 GND 0.00fF
C2865 a_50176_15846.n8 GND 0.00fF
C2866 a_50176_15846.n9 GND 0.00fF
C2867 a_50176_15846.t1 GND 0.02fF $ **FLOATING
C2868 a_50176_15846.t0 GND 0.02fF $ **FLOATING
C2869 a_50176_15846.n10 GND 0.05fF
C2870 a_50176_15846.n11 GND 0.00fF
C2871 a_50176_15846.n12 GND 0.00fF
C2872 a_50176_15846.n13 GND 0.02fF
C2873 a_50176_15846.n14 GND 0.04fF
C2874 a_50176_15846.n15 GND 0.12fF
C2875 a_50176_15846.n16 GND 0.01fF
C2876 a_50176_15846.n17 GND 0.12fF
C2877 a_50176_15846.t2 GND 3.87fF $ **FLOATING
C2878 a_50176_15846.n18 GND 0.52fF
C2879 a_50176_15846.t3 GND 0.24fF $ **FLOATING
C2880 a_40976_55366.n0 GND 0.01fF
C2881 a_40976_55366.n1 GND 0.01fF
C2882 a_40976_55366.n2 GND 0.00fF
C2883 a_40976_55366.n3 GND 0.00fF
C2884 a_40976_55366.n4 GND 0.00fF
C2885 a_40976_55366.n5 GND 0.00fF
C2886 a_40976_55366.n6 GND 0.00fF
C2887 a_40976_55366.n7 GND 0.00fF
C2888 a_40976_55366.n8 GND 0.00fF
C2889 a_40976_55366.n9 GND 0.00fF
C2890 a_40976_55366.t0 GND 0.02fF $ **FLOATING
C2891 a_40976_55366.t1 GND 0.02fF $ **FLOATING
C2892 a_40976_55366.n10 GND 0.05fF
C2893 a_40976_55366.n11 GND 0.00fF
C2894 a_40976_55366.n12 GND 0.00fF
C2895 a_40976_55366.n13 GND 0.02fF
C2896 a_40976_55366.n14 GND 0.04fF
C2897 a_40976_55366.n15 GND 0.12fF
C2898 a_40976_55366.n16 GND 0.01fF
C2899 a_40976_55366.n17 GND 0.12fF
C2900 a_40976_55366.t3 GND 3.87fF $ **FLOATING
C2901 a_40976_55366.n18 GND 0.52fF
C2902 a_40976_55366.t2 GND 0.24fF $ **FLOATING
C2903 a_41266_55442.n0 GND 0.00fF
C2904 a_41266_55442.n1 GND 0.00fF
C2905 a_41266_55442.n2 GND 0.01fF
C2906 a_41266_55442.n3 GND 0.01fF
C2907 a_41266_55442.n4 GND 0.00fF
C2908 a_41266_55442.n5 GND 0.00fF
C2909 a_41266_55442.n6 GND 0.00fF
C2910 a_41266_55442.n7 GND 0.00fF
C2911 a_41266_55442.n8 GND 0.00fF
C2912 a_41266_55442.n9 GND 0.00fF
C2913 a_41266_55442.n10 GND 0.09fF
C2914 a_41266_55442.n11 GND 0.00fF
C2915 a_41266_55442.n12 GND 0.01fF
C2916 a_41266_55442.n13 GND 0.01fF
C2917 a_41266_55442.n14 GND 0.01fF
C2918 a_41266_55442.n15 GND 0.00fF
C2919 a_41266_55442.n16 GND 0.00fF
C2920 a_41266_55442.n17 GND 0.00fF
C2921 a_41266_55442.t0 GND 0.02fF $ **FLOATING
C2922 a_41266_55442.n18 GND 0.07fF
C2923 a_41266_55442.n19 GND 0.02fF
C2924 a_41266_55442.n20 GND 0.05fF
C2925 a_41266_55442.n22 GND 0.04fF
C2926 a_41266_55442.n23 GND 0.04fF
C2927 a_41266_55442.n24 GND 0.00fF
C2928 a_41266_55442.n25 GND 0.00fF
C2929 a_41266_55442.t1 GND 0.02fF $ **FLOATING
C2930 a_41266_55442.n26 GND 0.07fF
C2931 a_41266_55442.n27 GND 0.02fF
C2932 a_41266_55442.n28 GND 0.05fF
C2933 a_41266_55442.n30 GND 0.01fF
C2934 a_41266_55442.n31 GND 0.00fF
C2935 a_41266_55442.n32 GND 0.00fF
C2936 a_41266_55442.n33 GND 0.00fF
C2937 a_41266_55442.n34 GND 0.00fF
C2938 a_41266_55442.n35 GND 0.00fF
C2939 a_41266_55442.n36 GND 0.00fF
C2940 a_41266_55442.n38 GND 0.08fF
C2941 a_41266_55442.t2 GND 4.19fF $ **FLOATING
C2942 a_41266_55442.n39 GND 0.61fF
C2943 a_41266_55442.t3 GND 0.26fF $ **FLOATING
C2944 a_22576_35606.n0 GND 0.01fF
C2945 a_22576_35606.n1 GND 0.01fF
C2946 a_22576_35606.n2 GND 0.00fF
C2947 a_22576_35606.n3 GND 0.00fF
C2948 a_22576_35606.n4 GND 0.00fF
C2949 a_22576_35606.n5 GND 0.00fF
C2950 a_22576_35606.n6 GND 0.00fF
C2951 a_22576_35606.n7 GND 0.00fF
C2952 a_22576_35606.n8 GND 0.00fF
C2953 a_22576_35606.n9 GND 0.00fF
C2954 a_22576_35606.t0 GND 0.02fF $ **FLOATING
C2955 a_22576_35606.t1 GND 0.02fF $ **FLOATING
C2956 a_22576_35606.n10 GND 0.05fF
C2957 a_22576_35606.n11 GND 0.00fF
C2958 a_22576_35606.n12 GND 0.00fF
C2959 a_22576_35606.n13 GND 0.02fF
C2960 a_22576_35606.n14 GND 0.04fF
C2961 a_22576_35606.n15 GND 0.12fF
C2962 a_22576_35606.n16 GND 0.01fF
C2963 a_22576_35606.n17 GND 0.12fF
C2964 a_22576_35606.t3 GND 3.87fF $ **FLOATING
C2965 a_22576_35606.n18 GND 0.52fF
C2966 a_22576_35606.t2 GND 0.24fF $ **FLOATING
C2967 a_22866_55442.n0 GND 0.00fF
C2968 a_22866_55442.n1 GND 0.00fF
C2969 a_22866_55442.n2 GND 0.01fF
C2970 a_22866_55442.n3 GND 0.01fF
C2971 a_22866_55442.n4 GND 0.00fF
C2972 a_22866_55442.n5 GND 0.00fF
C2973 a_22866_55442.n6 GND 0.00fF
C2974 a_22866_55442.n7 GND 0.00fF
C2975 a_22866_55442.n8 GND 0.00fF
C2976 a_22866_55442.n9 GND 0.00fF
C2977 a_22866_55442.n10 GND 0.09fF
C2978 a_22866_55442.n11 GND 0.00fF
C2979 a_22866_55442.n12 GND 0.01fF
C2980 a_22866_55442.n13 GND 0.01fF
C2981 a_22866_55442.n14 GND 0.01fF
C2982 a_22866_55442.n15 GND 0.00fF
C2983 a_22866_55442.n16 GND 0.00fF
C2984 a_22866_55442.n17 GND 0.00fF
C2985 a_22866_55442.t2 GND 0.02fF $ **FLOATING
C2986 a_22866_55442.n18 GND 0.07fF
C2987 a_22866_55442.n19 GND 0.02fF
C2988 a_22866_55442.n20 GND 0.05fF
C2989 a_22866_55442.n22 GND 0.04fF
C2990 a_22866_55442.n23 GND 0.04fF
C2991 a_22866_55442.n24 GND 0.00fF
C2992 a_22866_55442.n25 GND 0.00fF
C2993 a_22866_55442.t1 GND 0.02fF $ **FLOATING
C2994 a_22866_55442.n26 GND 0.07fF
C2995 a_22866_55442.n27 GND 0.02fF
C2996 a_22866_55442.n28 GND 0.05fF
C2997 a_22866_55442.n30 GND 0.01fF
C2998 a_22866_55442.n31 GND 0.00fF
C2999 a_22866_55442.n32 GND 0.00fF
C3000 a_22866_55442.n33 GND 0.00fF
C3001 a_22866_55442.n34 GND 0.00fF
C3002 a_22866_55442.n35 GND 0.00fF
C3003 a_22866_55442.n36 GND 0.00fF
C3004 a_22866_55442.n38 GND 0.08fF
C3005 a_22866_55442.t3 GND 4.19fF $ **FLOATING
C3006 a_22866_55442.n39 GND 0.61fF
C3007 a_22866_55442.t0 GND 0.26fF $ **FLOATING
C3008 a_32066_6042.n0 GND 0.00fF
C3009 a_32066_6042.n1 GND 0.00fF
C3010 a_32066_6042.n2 GND 0.01fF
C3011 a_32066_6042.n3 GND 0.01fF
C3012 a_32066_6042.n4 GND 0.00fF
C3013 a_32066_6042.n5 GND 0.00fF
C3014 a_32066_6042.n6 GND 0.00fF
C3015 a_32066_6042.n7 GND 0.00fF
C3016 a_32066_6042.n8 GND 0.00fF
C3017 a_32066_6042.n9 GND 0.00fF
C3018 a_32066_6042.n10 GND 0.09fF
C3019 a_32066_6042.n11 GND 0.00fF
C3020 a_32066_6042.n12 GND 0.01fF
C3021 a_32066_6042.n13 GND 0.01fF
C3022 a_32066_6042.n14 GND 0.01fF
C3023 a_32066_6042.n15 GND 0.00fF
C3024 a_32066_6042.n16 GND 0.00fF
C3025 a_32066_6042.n17 GND 0.00fF
C3026 a_32066_6042.t0 GND 0.02fF $ **FLOATING
C3027 a_32066_6042.n18 GND 0.07fF
C3028 a_32066_6042.n19 GND 0.02fF
C3029 a_32066_6042.n20 GND 0.05fF
C3030 a_32066_6042.n22 GND 0.04fF
C3031 a_32066_6042.n23 GND 0.04fF
C3032 a_32066_6042.n24 GND 0.00fF
C3033 a_32066_6042.n25 GND 0.00fF
C3034 a_32066_6042.t1 GND 0.02fF $ **FLOATING
C3035 a_32066_6042.n26 GND 0.07fF
C3036 a_32066_6042.n27 GND 0.02fF
C3037 a_32066_6042.n28 GND 0.05fF
C3038 a_32066_6042.n30 GND 0.01fF
C3039 a_32066_6042.n31 GND 0.00fF
C3040 a_32066_6042.n32 GND 0.00fF
C3041 a_32066_6042.n33 GND 0.00fF
C3042 a_32066_6042.n34 GND 0.00fF
C3043 a_32066_6042.n35 GND 0.00fF
C3044 a_32066_6042.n36 GND 0.00fF
C3045 a_32066_6042.n38 GND 0.08fF
C3046 a_32066_6042.t3 GND 4.19fF $ **FLOATING
C3047 a_32066_6042.n39 GND 0.61fF
C3048 a_32066_6042.t2 GND 0.26fF $ **FLOATING
C3049 a_68576_35606.n0 GND 0.01fF
C3050 a_68576_35606.n1 GND 0.01fF
C3051 a_68576_35606.n2 GND 0.00fF
C3052 a_68576_35606.n3 GND 0.00fF
C3053 a_68576_35606.n4 GND 0.00fF
C3054 a_68576_35606.n5 GND 0.00fF
C3055 a_68576_35606.n6 GND 0.00fF
C3056 a_68576_35606.n7 GND 0.00fF
C3057 a_68576_35606.n8 GND 0.00fF
C3058 a_68576_35606.n9 GND 0.00fF
C3059 a_68576_35606.t2 GND 0.02fF $ **FLOATING
C3060 a_68576_35606.t1 GND 0.02fF $ **FLOATING
C3061 a_68576_35606.n10 GND 0.05fF
C3062 a_68576_35606.n11 GND 0.00fF
C3063 a_68576_35606.n12 GND 0.00fF
C3064 a_68576_35606.n13 GND 0.02fF
C3065 a_68576_35606.n14 GND 0.04fF
C3066 a_68576_35606.n15 GND 0.12fF
C3067 a_68576_35606.n16 GND 0.01fF
C3068 a_68576_35606.n17 GND 0.12fF
C3069 a_68576_35606.t3 GND 3.87fF $ **FLOATING
C3070 a_68576_35606.n18 GND 0.52fF
C3071 a_68576_35606.t0 GND 0.24fF $ **FLOATING
C3072 a_40976_25726.n0 GND 0.01fF
C3073 a_40976_25726.n1 GND 0.01fF
C3074 a_40976_25726.n2 GND 0.00fF
C3075 a_40976_25726.n3 GND 0.00fF
C3076 a_40976_25726.n4 GND 0.00fF
C3077 a_40976_25726.n5 GND 0.00fF
C3078 a_40976_25726.n6 GND 0.00fF
C3079 a_40976_25726.n7 GND 0.00fF
C3080 a_40976_25726.n8 GND 0.00fF
C3081 a_40976_25726.n9 GND 0.00fF
C3082 a_40976_25726.t2 GND 0.02fF $ **FLOATING
C3083 a_40976_25726.t1 GND 0.02fF $ **FLOATING
C3084 a_40976_25726.n10 GND 0.05fF
C3085 a_40976_25726.n11 GND 0.00fF
C3086 a_40976_25726.n12 GND 0.00fF
C3087 a_40976_25726.n13 GND 0.02fF
C3088 a_40976_25726.n14 GND 0.04fF
C3089 a_40976_25726.n15 GND 0.12fF
C3090 a_40976_25726.n16 GND 0.01fF
C3091 a_40976_25726.n17 GND 0.12fF
C3092 a_40976_25726.t3 GND 3.87fF $ **FLOATING
C3093 a_40976_25726.n18 GND 0.52fF
C3094 a_40976_25726.t0 GND 0.24fF $ **FLOATING
C3095 a_4466_6042.n0 GND 0.00fF
C3096 a_4466_6042.n1 GND 0.00fF
C3097 a_4466_6042.n2 GND 0.01fF
C3098 a_4466_6042.n3 GND 0.01fF
C3099 a_4466_6042.n4 GND 0.00fF
C3100 a_4466_6042.n5 GND 0.00fF
C3101 a_4466_6042.n6 GND 0.00fF
C3102 a_4466_6042.n7 GND 0.00fF
C3103 a_4466_6042.n8 GND 0.00fF
C3104 a_4466_6042.n9 GND 0.00fF
C3105 a_4466_6042.n10 GND 0.09fF
C3106 a_4466_6042.n11 GND 0.00fF
C3107 a_4466_6042.n12 GND 0.01fF
C3108 a_4466_6042.n13 GND 0.01fF
C3109 a_4466_6042.n14 GND 0.01fF
C3110 a_4466_6042.n15 GND 0.00fF
C3111 a_4466_6042.n16 GND 0.00fF
C3112 a_4466_6042.n17 GND 0.00fF
C3113 a_4466_6042.t1 GND 0.02fF $ **FLOATING
C3114 a_4466_6042.n18 GND 0.07fF
C3115 a_4466_6042.n19 GND 0.02fF
C3116 a_4466_6042.n20 GND 0.05fF
C3117 a_4466_6042.n22 GND 0.04fF
C3118 a_4466_6042.n23 GND 0.04fF
C3119 a_4466_6042.n24 GND 0.00fF
C3120 a_4466_6042.n25 GND 0.00fF
C3121 a_4466_6042.t2 GND 0.02fF $ **FLOATING
C3122 a_4466_6042.n26 GND 0.07fF
C3123 a_4466_6042.n27 GND 0.02fF
C3124 a_4466_6042.n28 GND 0.05fF
C3125 a_4466_6042.n30 GND 0.01fF
C3126 a_4466_6042.n31 GND 0.00fF
C3127 a_4466_6042.n32 GND 0.00fF
C3128 a_4466_6042.n33 GND 0.00fF
C3129 a_4466_6042.n34 GND 0.00fF
C3130 a_4466_6042.n35 GND 0.00fF
C3131 a_4466_6042.n36 GND 0.00fF
C3132 a_4466_6042.n38 GND 0.08fF
C3133 a_4466_6042.t3 GND 4.19fF $ **FLOATING
C3134 a_4466_6042.n39 GND 0.61fF
C3135 a_4466_6042.t0 GND 0.26fF $ **FLOATING
C3136 a_13376_55366.n0 GND 0.01fF
C3137 a_13376_55366.n1 GND 0.01fF
C3138 a_13376_55366.n2 GND 0.00fF
C3139 a_13376_55366.n3 GND 0.00fF
C3140 a_13376_55366.n4 GND 0.00fF
C3141 a_13376_55366.n5 GND 0.00fF
C3142 a_13376_55366.n6 GND 0.00fF
C3143 a_13376_55366.n7 GND 0.00fF
C3144 a_13376_55366.n8 GND 0.00fF
C3145 a_13376_55366.n9 GND 0.00fF
C3146 a_13376_55366.t0 GND 0.02fF $ **FLOATING
C3147 a_13376_55366.t1 GND 0.02fF $ **FLOATING
C3148 a_13376_55366.n10 GND 0.05fF
C3149 a_13376_55366.n11 GND 0.00fF
C3150 a_13376_55366.n12 GND 0.00fF
C3151 a_13376_55366.n13 GND 0.02fF
C3152 a_13376_55366.n14 GND 0.04fF
C3153 a_13376_55366.n15 GND 0.12fF
C3154 a_13376_55366.n16 GND 0.01fF
C3155 a_13376_55366.n17 GND 0.12fF
C3156 a_13376_55366.t3 GND 3.87fF $ **FLOATING
C3157 a_13376_55366.n18 GND 0.52fF
C3158 a_13376_55366.t2 GND 0.24fF $ **FLOATING
C3159 a_13666_55442.n0 GND 0.00fF
C3160 a_13666_55442.n1 GND 0.00fF
C3161 a_13666_55442.n2 GND 0.01fF
C3162 a_13666_55442.n3 GND 0.01fF
C3163 a_13666_55442.n4 GND 0.00fF
C3164 a_13666_55442.n5 GND 0.00fF
C3165 a_13666_55442.n6 GND 0.00fF
C3166 a_13666_55442.n7 GND 0.00fF
C3167 a_13666_55442.n8 GND 0.00fF
C3168 a_13666_55442.n9 GND 0.00fF
C3169 a_13666_55442.n10 GND 0.09fF
C3170 a_13666_55442.n11 GND 0.00fF
C3171 a_13666_55442.n12 GND 0.01fF
C3172 a_13666_55442.n13 GND 0.01fF
C3173 a_13666_55442.n14 GND 0.01fF
C3174 a_13666_55442.n15 GND 0.00fF
C3175 a_13666_55442.n16 GND 0.00fF
C3176 a_13666_55442.n17 GND 0.00fF
C3177 a_13666_55442.t1 GND 0.02fF $ **FLOATING
C3178 a_13666_55442.n18 GND 0.07fF
C3179 a_13666_55442.n19 GND 0.02fF
C3180 a_13666_55442.n20 GND 0.05fF
C3181 a_13666_55442.n22 GND 0.04fF
C3182 a_13666_55442.n23 GND 0.04fF
C3183 a_13666_55442.n24 GND 0.00fF
C3184 a_13666_55442.n25 GND 0.00fF
C3185 a_13666_55442.t2 GND 0.02fF $ **FLOATING
C3186 a_13666_55442.n26 GND 0.07fF
C3187 a_13666_55442.n27 GND 0.02fF
C3188 a_13666_55442.n28 GND 0.05fF
C3189 a_13666_55442.n30 GND 0.01fF
C3190 a_13666_55442.n31 GND 0.00fF
C3191 a_13666_55442.n32 GND 0.00fF
C3192 a_13666_55442.n33 GND 0.00fF
C3193 a_13666_55442.n34 GND 0.00fF
C3194 a_13666_55442.n35 GND 0.00fF
C3195 a_13666_55442.n36 GND 0.00fF
C3196 a_13666_55442.n38 GND 0.08fF
C3197 a_13666_55442.t3 GND 4.19fF $ **FLOATING
C3198 a_13666_55442.n39 GND 0.61fF
C3199 a_13666_55442.t0 GND 0.26fF $ **FLOATING
C3200 a_32066_45562.n0 GND 0.00fF
C3201 a_32066_45562.n1 GND 0.00fF
C3202 a_32066_45562.n2 GND 0.01fF
C3203 a_32066_45562.n3 GND 0.01fF
C3204 a_32066_45562.n4 GND 0.00fF
C3205 a_32066_45562.n5 GND 0.00fF
C3206 a_32066_45562.n6 GND 0.00fF
C3207 a_32066_45562.n7 GND 0.00fF
C3208 a_32066_45562.n8 GND 0.00fF
C3209 a_32066_45562.n9 GND 0.00fF
C3210 a_32066_45562.n10 GND 0.09fF
C3211 a_32066_45562.n11 GND 0.00fF
C3212 a_32066_45562.n12 GND 0.01fF
C3213 a_32066_45562.n13 GND 0.01fF
C3214 a_32066_45562.n14 GND 0.01fF
C3215 a_32066_45562.n15 GND 0.00fF
C3216 a_32066_45562.n16 GND 0.00fF
C3217 a_32066_45562.n17 GND 0.00fF
C3218 a_32066_45562.t1 GND 0.02fF $ **FLOATING
C3219 a_32066_45562.n18 GND 0.07fF
C3220 a_32066_45562.n19 GND 0.02fF
C3221 a_32066_45562.n20 GND 0.05fF
C3222 a_32066_45562.n22 GND 0.04fF
C3223 a_32066_45562.n23 GND 0.04fF
C3224 a_32066_45562.n24 GND 0.00fF
C3225 a_32066_45562.n25 GND 0.00fF
C3226 a_32066_45562.t2 GND 0.02fF $ **FLOATING
C3227 a_32066_45562.n26 GND 0.07fF
C3228 a_32066_45562.n27 GND 0.02fF
C3229 a_32066_45562.n28 GND 0.05fF
C3230 a_32066_45562.n30 GND 0.01fF
C3231 a_32066_45562.n31 GND 0.00fF
C3232 a_32066_45562.n32 GND 0.00fF
C3233 a_32066_45562.n33 GND 0.00fF
C3234 a_32066_45562.n34 GND 0.00fF
C3235 a_32066_45562.n35 GND 0.00fF
C3236 a_32066_45562.n36 GND 0.00fF
C3237 a_32066_45562.n38 GND 0.08fF
C3238 a_32066_45562.t3 GND 4.19fF $ **FLOATING
C3239 a_32066_45562.n39 GND 0.61fF
C3240 a_32066_45562.t0 GND 0.26fF $ **FLOATING
C3241 a_13376_65246.n0 GND 0.01fF
C3242 a_13376_65246.n1 GND 0.01fF
C3243 a_13376_65246.n2 GND 0.00fF
C3244 a_13376_65246.n3 GND 0.00fF
C3245 a_13376_65246.n4 GND 0.00fF
C3246 a_13376_65246.n5 GND 0.00fF
C3247 a_13376_65246.n6 GND 0.00fF
C3248 a_13376_65246.n7 GND 0.00fF
C3249 a_13376_65246.n8 GND 0.00fF
C3250 a_13376_65246.n9 GND 0.00fF
C3251 a_13376_65246.t0 GND 0.02fF $ **FLOATING
C3252 a_13376_65246.t3 GND 0.02fF $ **FLOATING
C3253 a_13376_65246.n10 GND 0.05fF
C3254 a_13376_65246.n11 GND 0.00fF
C3255 a_13376_65246.n12 GND 0.00fF
C3256 a_13376_65246.n13 GND 0.02fF
C3257 a_13376_65246.n14 GND 0.04fF
C3258 a_13376_65246.n15 GND 0.12fF
C3259 a_13376_65246.n16 GND 0.01fF
C3260 a_13376_65246.n17 GND 0.12fF
C3261 a_13376_65246.t2 GND 3.87fF $ **FLOATING
C3262 a_13376_65246.n18 GND 0.52fF
C3263 a_13376_65246.t1 GND 0.24fF $ **FLOATING
C3264 a_4466_94962.n0 GND 0.00fF
C3265 a_4466_94962.n1 GND 0.00fF
C3266 a_4466_94962.n2 GND 0.01fF
C3267 a_4466_94962.n3 GND 0.01fF
C3268 a_4466_94962.n4 GND 0.00fF
C3269 a_4466_94962.n5 GND 0.00fF
C3270 a_4466_94962.n6 GND 0.00fF
C3271 a_4466_94962.n7 GND 0.00fF
C3272 a_4466_94962.n8 GND 0.00fF
C3273 a_4466_94962.n9 GND 0.00fF
C3274 a_4466_94962.n10 GND 0.09fF
C3275 a_4466_94962.n11 GND 0.00fF
C3276 a_4466_94962.n12 GND 0.01fF
C3277 a_4466_94962.n13 GND 0.01fF
C3278 a_4466_94962.n14 GND 0.01fF
C3279 a_4466_94962.n15 GND 0.00fF
C3280 a_4466_94962.n16 GND 0.00fF
C3281 a_4466_94962.n17 GND 0.00fF
C3282 a_4466_94962.t1 GND 0.02fF $ **FLOATING
C3283 a_4466_94962.n18 GND 0.07fF
C3284 a_4466_94962.n19 GND 0.02fF
C3285 a_4466_94962.n20 GND 0.05fF
C3286 a_4466_94962.n22 GND 0.04fF
C3287 a_4466_94962.n23 GND 0.04fF
C3288 a_4466_94962.n24 GND 0.00fF
C3289 a_4466_94962.n25 GND 0.00fF
C3290 a_4466_94962.t0 GND 0.02fF $ **FLOATING
C3291 a_4466_94962.n26 GND 0.07fF
C3292 a_4466_94962.n27 GND 0.02fF
C3293 a_4466_94962.n28 GND 0.05fF
C3294 a_4466_94962.n30 GND 0.01fF
C3295 a_4466_94962.n31 GND 0.00fF
C3296 a_4466_94962.n32 GND 0.00fF
C3297 a_4466_94962.n33 GND 0.00fF
C3298 a_4466_94962.n34 GND 0.00fF
C3299 a_4466_94962.n35 GND 0.00fF
C3300 a_4466_94962.n36 GND 0.00fF
C3301 a_4466_94962.n38 GND 0.08fF
C3302 a_4466_94962.t2 GND 4.19fF $ **FLOATING
C3303 a_4466_94962.n39 GND 0.61fF
C3304 a_4466_94962.t3 GND 0.26fF $ **FLOATING
C3305 a_4466_75202.n0 GND 0.00fF
C3306 a_4466_75202.n1 GND 0.00fF
C3307 a_4466_75202.n2 GND 0.01fF
C3308 a_4466_75202.n3 GND 0.01fF
C3309 a_4466_75202.n4 GND 0.00fF
C3310 a_4466_75202.n5 GND 0.00fF
C3311 a_4466_75202.n6 GND 0.00fF
C3312 a_4466_75202.n7 GND 0.00fF
C3313 a_4466_75202.n8 GND 0.00fF
C3314 a_4466_75202.n9 GND 0.00fF
C3315 a_4466_75202.n10 GND 0.09fF
C3316 a_4466_75202.n11 GND 0.00fF
C3317 a_4466_75202.n12 GND 0.01fF
C3318 a_4466_75202.n13 GND 0.01fF
C3319 a_4466_75202.n14 GND 0.01fF
C3320 a_4466_75202.n15 GND 0.00fF
C3321 a_4466_75202.n16 GND 0.00fF
C3322 a_4466_75202.n17 GND 0.00fF
C3323 a_4466_75202.t0 GND 0.02fF $ **FLOATING
C3324 a_4466_75202.n18 GND 0.07fF
C3325 a_4466_75202.n19 GND 0.02fF
C3326 a_4466_75202.n20 GND 0.05fF
C3327 a_4466_75202.n22 GND 0.04fF
C3328 a_4466_75202.n23 GND 0.04fF
C3329 a_4466_75202.n24 GND 0.00fF
C3330 a_4466_75202.n25 GND 0.00fF
C3331 a_4466_75202.t1 GND 0.02fF $ **FLOATING
C3332 a_4466_75202.n26 GND 0.07fF
C3333 a_4466_75202.n27 GND 0.02fF
C3334 a_4466_75202.n28 GND 0.05fF
C3335 a_4466_75202.n30 GND 0.01fF
C3336 a_4466_75202.n31 GND 0.00fF
C3337 a_4466_75202.n32 GND 0.00fF
C3338 a_4466_75202.n33 GND 0.00fF
C3339 a_4466_75202.n34 GND 0.00fF
C3340 a_4466_75202.n35 GND 0.00fF
C3341 a_4466_75202.n36 GND 0.00fF
C3342 a_4466_75202.n38 GND 0.08fF
C3343 a_4466_75202.t2 GND 4.19fF $ **FLOATING
C3344 a_4466_75202.n39 GND 0.61fF
C3345 a_4466_75202.t3 GND 0.26fF $ **FLOATING
C3346 a_4176_75126.n0 GND 0.01fF
C3347 a_4176_75126.n1 GND 0.01fF
C3348 a_4176_75126.n2 GND 0.00fF
C3349 a_4176_75126.n3 GND 0.00fF
C3350 a_4176_75126.n4 GND 0.00fF
C3351 a_4176_75126.n5 GND 0.00fF
C3352 a_4176_75126.n6 GND 0.00fF
C3353 a_4176_75126.n7 GND 0.00fF
C3354 a_4176_75126.n8 GND 0.00fF
C3355 a_4176_75126.n9 GND 0.00fF
C3356 a_4176_75126.t1 GND 0.02fF $ **FLOATING
C3357 a_4176_75126.t0 GND 0.02fF $ **FLOATING
C3358 a_4176_75126.n10 GND 0.05fF
C3359 a_4176_75126.n11 GND 0.00fF
C3360 a_4176_75126.n12 GND 0.00fF
C3361 a_4176_75126.n13 GND 0.02fF
C3362 a_4176_75126.n14 GND 0.04fF
C3363 a_4176_75126.n15 GND 0.12fF
C3364 a_4176_75126.n16 GND 0.01fF
C3365 a_4176_75126.n17 GND 0.12fF
C3366 a_4176_75126.t2 GND 3.87fF $ **FLOATING
C3367 a_4176_75126.n18 GND 0.52fF
C3368 a_4176_75126.t3 GND 0.24fF $ **FLOATING
C3369 bit2.t2 GND 0.02fF $ **FLOATING
C3370 bit2.n0 GND 0.01fF
C3371 bit2.n1 GND 0.00fF
C3372 bit2.t7 GND 0.02fF $ **FLOATING
C3373 bit2.n2 GND 0.01fF
C3374 bit2.n3 GND 0.00fF
C3375 bit2.n4 GND 0.00fF
C3376 bit2.n5 GND 0.00fF
C3377 bit2.n6 GND 0.07fF
C3378 bit2.t4 GND 0.02fF $ **FLOATING
C3379 bit2.n7 GND 0.01fF
C3380 bit2.n8 GND 0.00fF
C3381 bit2.t6 GND 0.02fF $ **FLOATING
C3382 bit2.n9 GND 0.01fF
C3383 bit2.n10 GND 0.00fF
C3384 bit2.n11 GND 0.00fF
C3385 bit2.n12 GND 0.00fF
C3386 bit2.n13 GND 0.07fF
C3387 bit2.t3 GND 0.02fF $ **FLOATING
C3388 bit2.n14 GND 0.01fF
C3389 bit2.n15 GND 0.00fF
C3390 bit2.t8 GND 0.02fF $ **FLOATING
C3391 bit2.n16 GND 0.01fF
C3392 bit2.n17 GND 0.00fF
C3393 bit2.n18 GND 0.00fF
C3394 bit2.n19 GND 0.00fF
C3395 bit2.n20 GND 0.07fF
C3396 bit2.n21 GND 0.00fF
C3397 bit2.n22 GND 0.00fF
C3398 bit2.t5 GND 0.02fF $ **FLOATING
C3399 bit2.n23 GND 0.01fF
C3400 bit2.n24 GND 0.00fF
C3401 bit2.t0 GND 0.02fF $ **FLOATING
C3402 bit2.n25 GND 0.01fF
C3403 bit2.n26 GND 0.00fF
C3404 bit2.n27 GND 0.07fF
C3405 bit2.t9 GND 0.01fF $ **FLOATING
C3406 bit2.t1 GND 0.01fF $ **FLOATING
C3407 bit2.n28 GND 0.02fF
C3408 bit2.n29 GND 17.50fF
C3409 bit2.n30 GND 17.17fF
C3410 bit2.n31 GND 17.17fF
C3411 bit2.n32 GND 55.56fF
C3412 a_22866_25802.n0 GND 0.00fF
C3413 a_22866_25802.n1 GND 0.00fF
C3414 a_22866_25802.n2 GND 0.01fF
C3415 a_22866_25802.n3 GND 0.01fF
C3416 a_22866_25802.n4 GND 0.00fF
C3417 a_22866_25802.n5 GND 0.00fF
C3418 a_22866_25802.n6 GND 0.00fF
C3419 a_22866_25802.n7 GND 0.00fF
C3420 a_22866_25802.n8 GND 0.00fF
C3421 a_22866_25802.n9 GND 0.00fF
C3422 a_22866_25802.n10 GND 0.09fF
C3423 a_22866_25802.n11 GND 0.00fF
C3424 a_22866_25802.n12 GND 0.01fF
C3425 a_22866_25802.n13 GND 0.01fF
C3426 a_22866_25802.n14 GND 0.01fF
C3427 a_22866_25802.n15 GND 0.00fF
C3428 a_22866_25802.n16 GND 0.00fF
C3429 a_22866_25802.n17 GND 0.00fF
C3430 a_22866_25802.t1 GND 0.02fF $ **FLOATING
C3431 a_22866_25802.n18 GND 0.07fF
C3432 a_22866_25802.n19 GND 0.02fF
C3433 a_22866_25802.n20 GND 0.05fF
C3434 a_22866_25802.n22 GND 0.04fF
C3435 a_22866_25802.n23 GND 0.04fF
C3436 a_22866_25802.n24 GND 0.00fF
C3437 a_22866_25802.n25 GND 0.00fF
C3438 a_22866_25802.t2 GND 0.02fF $ **FLOATING
C3439 a_22866_25802.n26 GND 0.07fF
C3440 a_22866_25802.n27 GND 0.02fF
C3441 a_22866_25802.n28 GND 0.05fF
C3442 a_22866_25802.n30 GND 0.01fF
C3443 a_22866_25802.n31 GND 0.00fF
C3444 a_22866_25802.n32 GND 0.00fF
C3445 a_22866_25802.n33 GND 0.00fF
C3446 a_22866_25802.n34 GND 0.00fF
C3447 a_22866_25802.n35 GND 0.00fF
C3448 a_22866_25802.n36 GND 0.00fF
C3449 a_22866_25802.n38 GND 0.08fF
C3450 a_22866_25802.t3 GND 4.19fF $ **FLOATING
C3451 a_22866_25802.n39 GND 0.61fF
C3452 a_22866_25802.t0 GND 0.26fF $ **FLOATING
C3453 a_22576_25726.n0 GND 0.01fF
C3454 a_22576_25726.n1 GND 0.01fF
C3455 a_22576_25726.n2 GND 0.00fF
C3456 a_22576_25726.n3 GND 0.00fF
C3457 a_22576_25726.n4 GND 0.00fF
C3458 a_22576_25726.n5 GND 0.00fF
C3459 a_22576_25726.n6 GND 0.00fF
C3460 a_22576_25726.n7 GND 0.00fF
C3461 a_22576_25726.n8 GND 0.00fF
C3462 a_22576_25726.n9 GND 0.00fF
C3463 a_22576_25726.t1 GND 0.02fF $ **FLOATING
C3464 a_22576_25726.t0 GND 0.02fF $ **FLOATING
C3465 a_22576_25726.n10 GND 0.05fF
C3466 a_22576_25726.n11 GND 0.00fF
C3467 a_22576_25726.n12 GND 0.00fF
C3468 a_22576_25726.n13 GND 0.02fF
C3469 a_22576_25726.n14 GND 0.04fF
C3470 a_22576_25726.n15 GND 0.12fF
C3471 a_22576_25726.n16 GND 0.01fF
C3472 a_22576_25726.n17 GND 0.12fF
C3473 a_22576_25726.t2 GND 3.87fF $ **FLOATING
C3474 a_22576_25726.n18 GND 0.52fF
C3475 a_22576_25726.t3 GND 0.24fF $ **FLOATING
C3476 a_4176_35606.n0 GND 0.01fF
C3477 a_4176_35606.n1 GND 0.01fF
C3478 a_4176_35606.n2 GND 0.00fF
C3479 a_4176_35606.n3 GND 0.00fF
C3480 a_4176_35606.n4 GND 0.00fF
C3481 a_4176_35606.n5 GND 0.00fF
C3482 a_4176_35606.n6 GND 0.00fF
C3483 a_4176_35606.n7 GND 0.00fF
C3484 a_4176_35606.n8 GND 0.00fF
C3485 a_4176_35606.n9 GND 0.00fF
C3486 a_4176_35606.t0 GND 0.02fF $ **FLOATING
C3487 a_4176_35606.t1 GND 0.02fF $ **FLOATING
C3488 a_4176_35606.n10 GND 0.05fF
C3489 a_4176_35606.n11 GND 0.00fF
C3490 a_4176_35606.n12 GND 0.00fF
C3491 a_4176_35606.n13 GND 0.02fF
C3492 a_4176_35606.n14 GND 0.04fF
C3493 a_4176_35606.n15 GND 0.12fF
C3494 a_4176_35606.n16 GND 0.01fF
C3495 a_4176_35606.n17 GND 0.12fF
C3496 a_4176_35606.t2 GND 3.87fF $ **FLOATING
C3497 a_4176_35606.n18 GND 0.52fF
C3498 a_4176_35606.t3 GND 0.24fF $ **FLOATING
C3499 a_4466_35682.n0 GND 0.00fF
C3500 a_4466_35682.n1 GND 0.00fF
C3501 a_4466_35682.n2 GND 0.01fF
C3502 a_4466_35682.n3 GND 0.01fF
C3503 a_4466_35682.n4 GND 0.00fF
C3504 a_4466_35682.n5 GND 0.00fF
C3505 a_4466_35682.n6 GND 0.00fF
C3506 a_4466_35682.n7 GND 0.00fF
C3507 a_4466_35682.n8 GND 0.00fF
C3508 a_4466_35682.n9 GND 0.00fF
C3509 a_4466_35682.n10 GND 0.09fF
C3510 a_4466_35682.n11 GND 0.00fF
C3511 a_4466_35682.n12 GND 0.01fF
C3512 a_4466_35682.n13 GND 0.01fF
C3513 a_4466_35682.n14 GND 0.01fF
C3514 a_4466_35682.n15 GND 0.00fF
C3515 a_4466_35682.n16 GND 0.00fF
C3516 a_4466_35682.n17 GND 0.00fF
C3517 a_4466_35682.t1 GND 0.02fF $ **FLOATING
C3518 a_4466_35682.n18 GND 0.07fF
C3519 a_4466_35682.n19 GND 0.02fF
C3520 a_4466_35682.n20 GND 0.05fF
C3521 a_4466_35682.n22 GND 0.04fF
C3522 a_4466_35682.n23 GND 0.04fF
C3523 a_4466_35682.n24 GND 0.00fF
C3524 a_4466_35682.n25 GND 0.00fF
C3525 a_4466_35682.t0 GND 0.02fF $ **FLOATING
C3526 a_4466_35682.n26 GND 0.07fF
C3527 a_4466_35682.n27 GND 0.02fF
C3528 a_4466_35682.n28 GND 0.05fF
C3529 a_4466_35682.n30 GND 0.01fF
C3530 a_4466_35682.n31 GND 0.00fF
C3531 a_4466_35682.n32 GND 0.00fF
C3532 a_4466_35682.n33 GND 0.00fF
C3533 a_4466_35682.n34 GND 0.00fF
C3534 a_4466_35682.n35 GND 0.00fF
C3535 a_4466_35682.n36 GND 0.00fF
C3536 a_4466_35682.n38 GND 0.08fF
C3537 a_4466_35682.t3 GND 4.19fF $ **FLOATING
C3538 a_4466_35682.n39 GND 0.61fF
C3539 a_4466_35682.t2 GND 0.26fF $ **FLOATING
C3540 a_4466_55442.n0 GND 0.00fF
C3541 a_4466_55442.n1 GND 0.00fF
C3542 a_4466_55442.n2 GND 0.01fF
C3543 a_4466_55442.n3 GND 0.01fF
C3544 a_4466_55442.n4 GND 0.00fF
C3545 a_4466_55442.n5 GND 0.00fF
C3546 a_4466_55442.n6 GND 0.00fF
C3547 a_4466_55442.n7 GND 0.00fF
C3548 a_4466_55442.n8 GND 0.00fF
C3549 a_4466_55442.n9 GND 0.00fF
C3550 a_4466_55442.n10 GND 0.09fF
C3551 a_4466_55442.n11 GND 0.00fF
C3552 a_4466_55442.n12 GND 0.01fF
C3553 a_4466_55442.n13 GND 0.01fF
C3554 a_4466_55442.n14 GND 0.01fF
C3555 a_4466_55442.n15 GND 0.00fF
C3556 a_4466_55442.n16 GND 0.00fF
C3557 a_4466_55442.n17 GND 0.00fF
C3558 a_4466_55442.t1 GND 0.02fF $ **FLOATING
C3559 a_4466_55442.n18 GND 0.07fF
C3560 a_4466_55442.n19 GND 0.02fF
C3561 a_4466_55442.n20 GND 0.05fF
C3562 a_4466_55442.n22 GND 0.04fF
C3563 a_4466_55442.n23 GND 0.04fF
C3564 a_4466_55442.n24 GND 0.00fF
C3565 a_4466_55442.n25 GND 0.00fF
C3566 a_4466_55442.t0 GND 0.02fF $ **FLOATING
C3567 a_4466_55442.n26 GND 0.07fF
C3568 a_4466_55442.n27 GND 0.02fF
C3569 a_4466_55442.n28 GND 0.05fF
C3570 a_4466_55442.n30 GND 0.01fF
C3571 a_4466_55442.n31 GND 0.00fF
C3572 a_4466_55442.n32 GND 0.00fF
C3573 a_4466_55442.n33 GND 0.00fF
C3574 a_4466_55442.n34 GND 0.00fF
C3575 a_4466_55442.n35 GND 0.00fF
C3576 a_4466_55442.n36 GND 0.00fF
C3577 a_4466_55442.n38 GND 0.08fF
C3578 a_4466_55442.t2 GND 4.19fF $ **FLOATING
C3579 a_4466_55442.n39 GND 0.61fF
C3580 a_4466_55442.t3 GND 0.26fF $ **FLOATING
C3581 a_50466_65322.n0 GND 0.00fF
C3582 a_50466_65322.n1 GND 0.00fF
C3583 a_50466_65322.n2 GND 0.01fF
C3584 a_50466_65322.n3 GND 0.01fF
C3585 a_50466_65322.n4 GND 0.00fF
C3586 a_50466_65322.n5 GND 0.00fF
C3587 a_50466_65322.n6 GND 0.00fF
C3588 a_50466_65322.n7 GND 0.00fF
C3589 a_50466_65322.n8 GND 0.00fF
C3590 a_50466_65322.n9 GND 0.00fF
C3591 a_50466_65322.n10 GND 0.09fF
C3592 a_50466_65322.n11 GND 0.00fF
C3593 a_50466_65322.n12 GND 0.01fF
C3594 a_50466_65322.n13 GND 0.01fF
C3595 a_50466_65322.n14 GND 0.01fF
C3596 a_50466_65322.n15 GND 0.00fF
C3597 a_50466_65322.n16 GND 0.00fF
C3598 a_50466_65322.n17 GND 0.00fF
C3599 a_50466_65322.t2 GND 0.02fF $ **FLOATING
C3600 a_50466_65322.n18 GND 0.07fF
C3601 a_50466_65322.n19 GND 0.02fF
C3602 a_50466_65322.n20 GND 0.05fF
C3603 a_50466_65322.n22 GND 0.04fF
C3604 a_50466_65322.n23 GND 0.04fF
C3605 a_50466_65322.n24 GND 0.00fF
C3606 a_50466_65322.n25 GND 0.00fF
C3607 a_50466_65322.t0 GND 0.02fF $ **FLOATING
C3608 a_50466_65322.n26 GND 0.07fF
C3609 a_50466_65322.n27 GND 0.02fF
C3610 a_50466_65322.n28 GND 0.05fF
C3611 a_50466_65322.n30 GND 0.01fF
C3612 a_50466_65322.n31 GND 0.00fF
C3613 a_50466_65322.n32 GND 0.00fF
C3614 a_50466_65322.n33 GND 0.00fF
C3615 a_50466_65322.n34 GND 0.00fF
C3616 a_50466_65322.n35 GND 0.00fF
C3617 a_50466_65322.n36 GND 0.00fF
C3618 a_50466_65322.n38 GND 0.08fF
C3619 a_50466_65322.t1 GND 4.19fF $ **FLOATING
C3620 a_50466_65322.n39 GND 0.61fF
C3621 a_50466_65322.t3 GND 0.26fF $ **FLOATING
C3622 a_22576_55366.n0 GND 0.01fF
C3623 a_22576_55366.n1 GND 0.01fF
C3624 a_22576_55366.n2 GND 0.00fF
C3625 a_22576_55366.n3 GND 0.00fF
C3626 a_22576_55366.n4 GND 0.00fF
C3627 a_22576_55366.n5 GND 0.00fF
C3628 a_22576_55366.n6 GND 0.00fF
C3629 a_22576_55366.n7 GND 0.00fF
C3630 a_22576_55366.n8 GND 0.00fF
C3631 a_22576_55366.n9 GND 0.00fF
C3632 a_22576_55366.t0 GND 0.02fF $ **FLOATING
C3633 a_22576_55366.t1 GND 0.02fF $ **FLOATING
C3634 a_22576_55366.n10 GND 0.05fF
C3635 a_22576_55366.n11 GND 0.00fF
C3636 a_22576_55366.n12 GND 0.00fF
C3637 a_22576_55366.n13 GND 0.02fF
C3638 a_22576_55366.n14 GND 0.04fF
C3639 a_22576_55366.n15 GND 0.12fF
C3640 a_22576_55366.n16 GND 0.01fF
C3641 a_22576_55366.n17 GND 0.12fF
C3642 a_22576_55366.t3 GND 3.87fF $ **FLOATING
C3643 a_22576_55366.n18 GND 0.52fF
C3644 a_22576_55366.t2 GND 0.24fF $ **FLOATING
C3645 a_n436_64726.t9 GND 0.04fF $ **FLOATING
C3646 a_n436_64726.t3 GND 0.07fF $ **FLOATING
C3647 a_n436_64726.t5 GND 0.07fF $ **FLOATING
C3648 a_n436_64726.t8 GND 0.07fF $ **FLOATING
C3649 a_n436_64726.t4 GND 0.07fF $ **FLOATING
C3650 a_n436_64726.t10 GND 0.07fF $ **FLOATING
C3651 a_n436_64726.t13 GND 0.07fF $ **FLOATING
C3652 a_n436_64726.t12 GND 0.07fF $ **FLOATING
C3653 a_n436_64726.t14 GND 0.07fF $ **FLOATING
C3654 a_n436_64726.t6 GND 0.07fF $ **FLOATING
C3655 a_n436_64726.t1 GND 0.07fF $ **FLOATING
C3656 a_n436_64726.t11 GND 0.07fF $ **FLOATING
C3657 a_n436_64726.t15 GND 0.07fF $ **FLOATING
C3658 a_n436_64726.t16 GND 0.07fF $ **FLOATING
C3659 a_n436_64726.t0 GND 0.07fF $ **FLOATING
C3660 a_n436_64726.t17 GND 0.07fF $ **FLOATING
C3661 a_n436_64726.t7 GND 0.12fF $ **FLOATING
C3662 a_n436_64726.n0 GND 21.26fF
C3663 a_n436_64726.n1 GND 10.63fF
C3664 a_n436_64726.n2 GND 10.63fF
C3665 a_n436_64726.n3 GND 10.63fF
C3666 a_n436_64726.n4 GND 10.63fF
C3667 a_n436_64726.n5 GND 10.63fF
C3668 a_n436_64726.n6 GND 10.63fF
C3669 a_n436_64726.n7 GND 10.63fF
C3670 a_n436_64726.n8 GND 10.63fF
C3671 a_n436_64726.n9 GND 10.63fF
C3672 a_n436_64726.n10 GND 10.63fF
C3673 a_n436_64726.n11 GND 10.63fF
C3674 a_n436_64726.n12 GND 10.63fF
C3675 a_n436_64726.n13 GND 10.63fF
C3676 a_n436_64726.n14 GND 12.04fF
C3677 a_n436_64726.n15 GND 0.06fF
C3678 a_n436_64726.t2 GND 0.09fF $ **FLOATING
C3679 a_4466_65322.n0 GND 0.00fF
C3680 a_4466_65322.n1 GND 0.00fF
C3681 a_4466_65322.n2 GND 0.01fF
C3682 a_4466_65322.n3 GND 0.01fF
C3683 a_4466_65322.n4 GND 0.00fF
C3684 a_4466_65322.n5 GND 0.00fF
C3685 a_4466_65322.n6 GND 0.00fF
C3686 a_4466_65322.n7 GND 0.00fF
C3687 a_4466_65322.n8 GND 0.00fF
C3688 a_4466_65322.n9 GND 0.00fF
C3689 a_4466_65322.n10 GND 0.09fF
C3690 a_4466_65322.n11 GND 0.00fF
C3691 a_4466_65322.n12 GND 0.01fF
C3692 a_4466_65322.n13 GND 0.01fF
C3693 a_4466_65322.n14 GND 0.01fF
C3694 a_4466_65322.n15 GND 0.00fF
C3695 a_4466_65322.n16 GND 0.00fF
C3696 a_4466_65322.n17 GND 0.00fF
C3697 a_4466_65322.t3 GND 0.02fF $ **FLOATING
C3698 a_4466_65322.n18 GND 0.07fF
C3699 a_4466_65322.n19 GND 0.02fF
C3700 a_4466_65322.n20 GND 0.05fF
C3701 a_4466_65322.n22 GND 0.04fF
C3702 a_4466_65322.n23 GND 0.04fF
C3703 a_4466_65322.n24 GND 0.00fF
C3704 a_4466_65322.n25 GND 0.00fF
C3705 a_4466_65322.t0 GND 0.02fF $ **FLOATING
C3706 a_4466_65322.n26 GND 0.07fF
C3707 a_4466_65322.n27 GND 0.02fF
C3708 a_4466_65322.n28 GND 0.05fF
C3709 a_4466_65322.n30 GND 0.01fF
C3710 a_4466_65322.n31 GND 0.00fF
C3711 a_4466_65322.n32 GND 0.00fF
C3712 a_4466_65322.n33 GND 0.00fF
C3713 a_4466_65322.n34 GND 0.00fF
C3714 a_4466_65322.n35 GND 0.00fF
C3715 a_4466_65322.n36 GND 0.00fF
C3716 a_4466_65322.n38 GND 0.08fF
C3717 a_4466_65322.t2 GND 4.19fF $ **FLOATING
C3718 a_4466_65322.n39 GND 0.61fF
C3719 a_4466_65322.t1 GND 0.26fF $ **FLOATING
C3720 a_31776_55366.n0 GND 0.01fF
C3721 a_31776_55366.n1 GND 0.01fF
C3722 a_31776_55366.n2 GND 0.00fF
C3723 a_31776_55366.n3 GND 0.00fF
C3724 a_31776_55366.n4 GND 0.00fF
C3725 a_31776_55366.n5 GND 0.00fF
C3726 a_31776_55366.n6 GND 0.00fF
C3727 a_31776_55366.n7 GND 0.00fF
C3728 a_31776_55366.n8 GND 0.00fF
C3729 a_31776_55366.n9 GND 0.00fF
C3730 a_31776_55366.t0 GND 0.02fF $ **FLOATING
C3731 a_31776_55366.t1 GND 0.02fF $ **FLOATING
C3732 a_31776_55366.n10 GND 0.05fF
C3733 a_31776_55366.n11 GND 0.00fF
C3734 a_31776_55366.n12 GND 0.00fF
C3735 a_31776_55366.n13 GND 0.02fF
C3736 a_31776_55366.n14 GND 0.04fF
C3737 a_31776_55366.n15 GND 0.12fF
C3738 a_31776_55366.n16 GND 0.01fF
C3739 a_31776_55366.n17 GND 0.12fF
C3740 a_31776_55366.t3 GND 3.87fF $ **FLOATING
C3741 a_31776_55366.n18 GND 0.52fF
C3742 a_31776_55366.t2 GND 0.24fF $ **FLOATING
C3743 a_32066_55442.n0 GND 0.00fF
C3744 a_32066_55442.n1 GND 0.00fF
C3745 a_32066_55442.n2 GND 0.01fF
C3746 a_32066_55442.n3 GND 0.01fF
C3747 a_32066_55442.n4 GND 0.00fF
C3748 a_32066_55442.n5 GND 0.00fF
C3749 a_32066_55442.n6 GND 0.00fF
C3750 a_32066_55442.n7 GND 0.00fF
C3751 a_32066_55442.n8 GND 0.00fF
C3752 a_32066_55442.n9 GND 0.00fF
C3753 a_32066_55442.n10 GND 0.09fF
C3754 a_32066_55442.n11 GND 0.00fF
C3755 a_32066_55442.n12 GND 0.01fF
C3756 a_32066_55442.n13 GND 0.01fF
C3757 a_32066_55442.n14 GND 0.01fF
C3758 a_32066_55442.n15 GND 0.00fF
C3759 a_32066_55442.n16 GND 0.00fF
C3760 a_32066_55442.n17 GND 0.00fF
C3761 a_32066_55442.t1 GND 0.02fF $ **FLOATING
C3762 a_32066_55442.n18 GND 0.07fF
C3763 a_32066_55442.n19 GND 0.02fF
C3764 a_32066_55442.n20 GND 0.05fF
C3765 a_32066_55442.n22 GND 0.04fF
C3766 a_32066_55442.n23 GND 0.04fF
C3767 a_32066_55442.n24 GND 0.00fF
C3768 a_32066_55442.n25 GND 0.00fF
C3769 a_32066_55442.t2 GND 0.02fF $ **FLOATING
C3770 a_32066_55442.n26 GND 0.07fF
C3771 a_32066_55442.n27 GND 0.02fF
C3772 a_32066_55442.n28 GND 0.05fF
C3773 a_32066_55442.n30 GND 0.01fF
C3774 a_32066_55442.n31 GND 0.00fF
C3775 a_32066_55442.n32 GND 0.00fF
C3776 a_32066_55442.n33 GND 0.00fF
C3777 a_32066_55442.n34 GND 0.00fF
C3778 a_32066_55442.n35 GND 0.00fF
C3779 a_32066_55442.n36 GND 0.00fF
C3780 a_32066_55442.n38 GND 0.08fF
C3781 a_32066_55442.t3 GND 4.19fF $ **FLOATING
C3782 a_32066_55442.n39 GND 0.61fF
C3783 a_32066_55442.t0 GND 0.26fF $ **FLOATING
C3784 a_41266_15922.n0 GND 0.00fF
C3785 a_41266_15922.n1 GND 0.00fF
C3786 a_41266_15922.n2 GND 0.01fF
C3787 a_41266_15922.n3 GND 0.01fF
C3788 a_41266_15922.n4 GND 0.00fF
C3789 a_41266_15922.n5 GND 0.00fF
C3790 a_41266_15922.n6 GND 0.00fF
C3791 a_41266_15922.n7 GND 0.00fF
C3792 a_41266_15922.n8 GND 0.00fF
C3793 a_41266_15922.n9 GND 0.00fF
C3794 a_41266_15922.n10 GND 0.09fF
C3795 a_41266_15922.n11 GND 0.00fF
C3796 a_41266_15922.n12 GND 0.01fF
C3797 a_41266_15922.n13 GND 0.01fF
C3798 a_41266_15922.n14 GND 0.01fF
C3799 a_41266_15922.n15 GND 0.00fF
C3800 a_41266_15922.n16 GND 0.00fF
C3801 a_41266_15922.n17 GND 0.00fF
C3802 a_41266_15922.t1 GND 0.02fF $ **FLOATING
C3803 a_41266_15922.n18 GND 0.07fF
C3804 a_41266_15922.n19 GND 0.02fF
C3805 a_41266_15922.n20 GND 0.05fF
C3806 a_41266_15922.n22 GND 0.04fF
C3807 a_41266_15922.n23 GND 0.04fF
C3808 a_41266_15922.n24 GND 0.00fF
C3809 a_41266_15922.n25 GND 0.00fF
C3810 a_41266_15922.t2 GND 0.02fF $ **FLOATING
C3811 a_41266_15922.n26 GND 0.07fF
C3812 a_41266_15922.n27 GND 0.02fF
C3813 a_41266_15922.n28 GND 0.05fF
C3814 a_41266_15922.n30 GND 0.01fF
C3815 a_41266_15922.n31 GND 0.00fF
C3816 a_41266_15922.n32 GND 0.00fF
C3817 a_41266_15922.n33 GND 0.00fF
C3818 a_41266_15922.n34 GND 0.00fF
C3819 a_41266_15922.n35 GND 0.00fF
C3820 a_41266_15922.n36 GND 0.00fF
C3821 a_41266_15922.n38 GND 0.08fF
C3822 a_41266_15922.t3 GND 4.19fF $ **FLOATING
C3823 a_41266_15922.n39 GND 0.61fF
C3824 a_41266_15922.t0 GND 0.26fF $ **FLOATING
C3825 a_40976_15846.n0 GND 0.01fF
C3826 a_40976_15846.n1 GND 0.01fF
C3827 a_40976_15846.n2 GND 0.00fF
C3828 a_40976_15846.n3 GND 0.00fF
C3829 a_40976_15846.n4 GND 0.00fF
C3830 a_40976_15846.n5 GND 0.00fF
C3831 a_40976_15846.n6 GND 0.00fF
C3832 a_40976_15846.n7 GND 0.00fF
C3833 a_40976_15846.n8 GND 0.00fF
C3834 a_40976_15846.n9 GND 0.00fF
C3835 a_40976_15846.t1 GND 0.02fF $ **FLOATING
C3836 a_40976_15846.t0 GND 0.02fF $ **FLOATING
C3837 a_40976_15846.n10 GND 0.05fF
C3838 a_40976_15846.n11 GND 0.00fF
C3839 a_40976_15846.n12 GND 0.00fF
C3840 a_40976_15846.n13 GND 0.02fF
C3841 a_40976_15846.n14 GND 0.04fF
C3842 a_40976_15846.n15 GND 0.12fF
C3843 a_40976_15846.n16 GND 0.01fF
C3844 a_40976_15846.n17 GND 0.12fF
C3845 a_40976_15846.t2 GND 3.87fF $ **FLOATING
C3846 a_40976_15846.n18 GND 0.52fF
C3847 a_40976_15846.t3 GND 0.24fF $ **FLOATING
C3848 a_13376_35606.n0 GND 0.01fF
C3849 a_13376_35606.n1 GND 0.01fF
C3850 a_13376_35606.n2 GND 0.00fF
C3851 a_13376_35606.n3 GND 0.00fF
C3852 a_13376_35606.n4 GND 0.00fF
C3853 a_13376_35606.n5 GND 0.00fF
C3854 a_13376_35606.n6 GND 0.00fF
C3855 a_13376_35606.n7 GND 0.00fF
C3856 a_13376_35606.n8 GND 0.00fF
C3857 a_13376_35606.n9 GND 0.00fF
C3858 a_13376_35606.t1 GND 0.02fF $ **FLOATING
C3859 a_13376_35606.t0 GND 0.02fF $ **FLOATING
C3860 a_13376_35606.n10 GND 0.05fF
C3861 a_13376_35606.n11 GND 0.00fF
C3862 a_13376_35606.n12 GND 0.00fF
C3863 a_13376_35606.n13 GND 0.02fF
C3864 a_13376_35606.n14 GND 0.04fF
C3865 a_13376_35606.n15 GND 0.12fF
C3866 a_13376_35606.n16 GND 0.01fF
C3867 a_13376_35606.n17 GND 0.12fF
C3868 a_13376_35606.t2 GND 3.87fF $ **FLOATING
C3869 a_13376_35606.n18 GND 0.52fF
C3870 a_13376_35606.t3 GND 0.24fF $ **FLOATING
C3871 a_59666_55442.n0 GND 0.00fF
C3872 a_59666_55442.n1 GND 0.00fF
C3873 a_59666_55442.n2 GND 0.01fF
C3874 a_59666_55442.n3 GND 0.01fF
C3875 a_59666_55442.n4 GND 0.00fF
C3876 a_59666_55442.n5 GND 0.00fF
C3877 a_59666_55442.n6 GND 0.00fF
C3878 a_59666_55442.n7 GND 0.00fF
C3879 a_59666_55442.n8 GND 0.00fF
C3880 a_59666_55442.n9 GND 0.00fF
C3881 a_59666_55442.n10 GND 0.09fF
C3882 a_59666_55442.n11 GND 0.00fF
C3883 a_59666_55442.n12 GND 0.01fF
C3884 a_59666_55442.n13 GND 0.01fF
C3885 a_59666_55442.n14 GND 0.01fF
C3886 a_59666_55442.n15 GND 0.00fF
C3887 a_59666_55442.n16 GND 0.00fF
C3888 a_59666_55442.n17 GND 0.00fF
C3889 a_59666_55442.t1 GND 0.02fF $ **FLOATING
C3890 a_59666_55442.n18 GND 0.07fF
C3891 a_59666_55442.n19 GND 0.02fF
C3892 a_59666_55442.n20 GND 0.05fF
C3893 a_59666_55442.n22 GND 0.04fF
C3894 a_59666_55442.n23 GND 0.04fF
C3895 a_59666_55442.n24 GND 0.00fF
C3896 a_59666_55442.n25 GND 0.00fF
C3897 a_59666_55442.t2 GND 0.02fF $ **FLOATING
C3898 a_59666_55442.n26 GND 0.07fF
C3899 a_59666_55442.n27 GND 0.02fF
C3900 a_59666_55442.n28 GND 0.05fF
C3901 a_59666_55442.n30 GND 0.01fF
C3902 a_59666_55442.n31 GND 0.00fF
C3903 a_59666_55442.n32 GND 0.00fF
C3904 a_59666_55442.n33 GND 0.00fF
C3905 a_59666_55442.n34 GND 0.00fF
C3906 a_59666_55442.n35 GND 0.00fF
C3907 a_59666_55442.n36 GND 0.00fF
C3908 a_59666_55442.n38 GND 0.08fF
C3909 a_59666_55442.t3 GND 4.19fF $ **FLOATING
C3910 a_59666_55442.n39 GND 0.61fF
C3911 a_59666_55442.t0 GND 0.26fF $ **FLOATING
C3912 a_31776_45486.n0 GND 0.01fF
C3913 a_31776_45486.n1 GND 0.01fF
C3914 a_31776_45486.n2 GND 0.00fF
C3915 a_31776_45486.n3 GND 0.00fF
C3916 a_31776_45486.n4 GND 0.00fF
C3917 a_31776_45486.n5 GND 0.00fF
C3918 a_31776_45486.n6 GND 0.00fF
C3919 a_31776_45486.n7 GND 0.00fF
C3920 a_31776_45486.n8 GND 0.00fF
C3921 a_31776_45486.n9 GND 0.00fF
C3922 a_31776_45486.t2 GND 0.02fF $ **FLOATING
C3923 a_31776_45486.t1 GND 0.02fF $ **FLOATING
C3924 a_31776_45486.n10 GND 0.05fF
C3925 a_31776_45486.n11 GND 0.00fF
C3926 a_31776_45486.n12 GND 0.00fF
C3927 a_31776_45486.n13 GND 0.02fF
C3928 a_31776_45486.n14 GND 0.04fF
C3929 a_31776_45486.n15 GND 0.12fF
C3930 a_31776_45486.n16 GND 0.01fF
C3931 a_31776_45486.n17 GND 0.12fF
C3932 a_31776_45486.t3 GND 3.87fF $ **FLOATING
C3933 a_31776_45486.n18 GND 0.52fF
C3934 a_31776_45486.t0 GND 0.24fF $ **FLOATING
C3935 a_68866_35682.n0 GND 0.00fF
C3936 a_68866_35682.n1 GND 0.00fF
C3937 a_68866_35682.n2 GND 0.01fF
C3938 a_68866_35682.n3 GND 0.01fF
C3939 a_68866_35682.n4 GND 0.00fF
C3940 a_68866_35682.n5 GND 0.00fF
C3941 a_68866_35682.n6 GND 0.00fF
C3942 a_68866_35682.n7 GND 0.00fF
C3943 a_68866_35682.n8 GND 0.00fF
C3944 a_68866_35682.n9 GND 0.00fF
C3945 a_68866_35682.n10 GND 0.09fF
C3946 a_68866_35682.n11 GND 0.00fF
C3947 a_68866_35682.n12 GND 0.01fF
C3948 a_68866_35682.n13 GND 0.01fF
C3949 a_68866_35682.n14 GND 0.01fF
C3950 a_68866_35682.n15 GND 0.00fF
C3951 a_68866_35682.n16 GND 0.00fF
C3952 a_68866_35682.n17 GND 0.00fF
C3953 a_68866_35682.t1 GND 0.02fF $ **FLOATING
C3954 a_68866_35682.n18 GND 0.07fF
C3955 a_68866_35682.n19 GND 0.02fF
C3956 a_68866_35682.n20 GND 0.05fF
C3957 a_68866_35682.n22 GND 0.04fF
C3958 a_68866_35682.n23 GND 0.04fF
C3959 a_68866_35682.n24 GND 0.00fF
C3960 a_68866_35682.n25 GND 0.00fF
C3961 a_68866_35682.t0 GND 0.02fF $ **FLOATING
C3962 a_68866_35682.n26 GND 0.07fF
C3963 a_68866_35682.n27 GND 0.02fF
C3964 a_68866_35682.n28 GND 0.05fF
C3965 a_68866_35682.n30 GND 0.01fF
C3966 a_68866_35682.n31 GND 0.00fF
C3967 a_68866_35682.n32 GND 0.00fF
C3968 a_68866_35682.n33 GND 0.00fF
C3969 a_68866_35682.n34 GND 0.00fF
C3970 a_68866_35682.n35 GND 0.00fF
C3971 a_68866_35682.n36 GND 0.00fF
C3972 a_68866_35682.n38 GND 0.08fF
C3973 a_68866_35682.t2 GND 4.19fF $ **FLOATING
C3974 a_68866_35682.n39 GND 0.61fF
C3975 a_68866_35682.t3 GND 0.26fF $ **FLOATING
C3976 OUT_N.t13 GND 0.48fF $ **FLOATING
C3977 OUT_N.t51 GND 0.48fF $ **FLOATING
C3978 OUT_N.t25 GND 0.48fF $ **FLOATING
C3979 OUT_N.t0 GND 0.48fF $ **FLOATING
C3980 OUT_N.t48 GND 0.48fF $ **FLOATING
C3981 OUT_N.t19 GND 0.48fF $ **FLOATING
C3982 OUT_N.t9 GND 3.91fF $ **FLOATING
C3983 OUT_N.n0 GND 14.21fF
C3984 OUT_N.n1 GND 12.29fF
C3985 OUT_N.n2 GND 12.29fF
C3986 OUT_N.n3 GND 12.29fF
C3987 OUT_N.n4 GND 12.29fF
C3988 OUT_N.n5 GND 32.90fF
C3989 OUT_N.t26 GND 0.48fF $ **FLOATING
C3990 OUT_N.t1 GND 0.48fF $ **FLOATING
C3991 OUT_N.t42 GND 0.48fF $ **FLOATING
C3992 OUT_N.t14 GND 0.48fF $ **FLOATING
C3993 OUT_N.t58 GND 0.48fF $ **FLOATING
C3994 OUT_N.t35 GND 0.48fF $ **FLOATING
C3995 OUT_N.t36 GND 3.91fF $ **FLOATING
C3996 OUT_N.n6 GND 14.21fF
C3997 OUT_N.n7 GND 12.29fF
C3998 OUT_N.n8 GND 12.29fF
C3999 OUT_N.n9 GND 12.29fF
C4000 OUT_N.n10 GND 12.29fF
C4001 OUT_N.n11 GND 32.90fF
C4002 OUT_N.t2 GND 0.48fF $ **FLOATING
C4003 OUT_N.t43 GND 0.48fF $ **FLOATING
C4004 OUT_N.t16 GND 0.48fF $ **FLOATING
C4005 OUT_N.t55 GND 0.48fF $ **FLOATING
C4006 OUT_N.t37 GND 0.48fF $ **FLOATING
C4007 OUT_N.t8 GND 0.48fF $ **FLOATING
C4008 OUT_N.t30 GND 3.91fF $ **FLOATING
C4009 OUT_N.n12 GND 14.21fF
C4010 OUT_N.n13 GND 12.29fF
C4011 OUT_N.n14 GND 12.29fF
C4012 OUT_N.n15 GND 12.29fF
C4013 OUT_N.n16 GND 12.29fF
C4014 OUT_N.n17 GND 32.91fF
C4015 OUT_N.t46 GND 0.48fF $ **FLOATING
C4016 OUT_N.t18 GND 0.48fF $ **FLOATING
C4017 OUT_N.t56 GND 0.48fF $ **FLOATING
C4018 OUT_N.t32 GND 0.48fF $ **FLOATING
C4019 OUT_N.t10 GND 0.48fF $ **FLOATING
C4020 OUT_N.t50 GND 0.48fF $ **FLOATING
C4021 OUT_N.t24 GND 3.91fF $ **FLOATING
C4022 OUT_N.n18 GND 14.21fF
C4023 OUT_N.n19 GND 12.29fF
C4024 OUT_N.n20 GND 12.29fF
C4025 OUT_N.n21 GND 12.29fF
C4026 OUT_N.n22 GND 12.29fF
C4027 OUT_N.n23 GND 32.91fF
C4028 OUT_N.t15 GND 0.48fF $ **FLOATING
C4029 OUT_N.t54 GND 0.48fF $ **FLOATING
C4030 OUT_N.t29 GND 0.48fF $ **FLOATING
C4031 OUT_N.t5 GND 0.48fF $ **FLOATING
C4032 OUT_N.t45 GND 0.48fF $ **FLOATING
C4033 OUT_N.t22 GND 0.48fF $ **FLOATING
C4034 OUT_N.t61 GND 0.48fF $ **FLOATING
C4035 OUT_N.t33 GND 3.91fF $ **FLOATING
C4036 OUT_N.n24 GND 14.21fF
C4037 OUT_N.n25 GND 12.29fF
C4038 OUT_N.n26 GND 12.29fF
C4039 OUT_N.n27 GND 12.29fF
C4040 OUT_N.n28 GND 12.29fF
C4041 OUT_N.n29 GND 12.29fF
C4042 OUT_N.n30 GND 26.78fF
C4043 OUT_N.t57 GND 0.48fF $ **FLOATING
C4044 OUT_N.t31 GND 0.48fF $ **FLOATING
C4045 OUT_N.t6 GND 0.48fF $ **FLOATING
C4046 OUT_N.t47 GND 0.48fF $ **FLOATING
C4047 OUT_N.t20 GND 0.48fF $ **FLOATING
C4048 OUT_N.t62 GND 0.48fF $ **FLOATING
C4049 OUT_N.t39 GND 0.48fF $ **FLOATING
C4050 OUT_N.t27 GND 3.91fF $ **FLOATING
C4051 OUT_N.n31 GND 14.21fF
C4052 OUT_N.n32 GND 12.29fF
C4053 OUT_N.n33 GND 12.29fF
C4054 OUT_N.n34 GND 12.29fF
C4055 OUT_N.n35 GND 12.29fF
C4056 OUT_N.n36 GND 12.29fF
C4057 OUT_N.n37 GND 26.78fF
C4058 OUT_N.t52 GND 0.48fF $ **FLOATING
C4059 OUT_N.t34 GND 0.48fF $ **FLOATING
C4060 OUT_N.t7 GND 0.48fF $ **FLOATING
C4061 OUT_N.t49 GND 0.48fF $ **FLOATING
C4062 OUT_N.t21 GND 0.48fF $ **FLOATING
C4063 OUT_N.t59 GND 0.48fF $ **FLOATING
C4064 OUT_N.t40 GND 0.48fF $ **FLOATING
C4065 OUT_N.t11 GND 0.48fF $ **FLOATING
C4066 OUT_N.t23 GND 3.91fF $ **FLOATING
C4067 OUT_N.n38 GND 14.21fF
C4068 OUT_N.n39 GND 12.29fF
C4069 OUT_N.n40 GND 12.29fF
C4070 OUT_N.n41 GND 12.29fF
C4071 OUT_N.n42 GND 12.29fF
C4072 OUT_N.n43 GND 12.29fF
C4073 OUT_N.n44 GND 12.29fF
C4074 OUT_N.n45 GND 20.66fF
C4075 OUT_N.t4 GND 0.48fF $ **FLOATING
C4076 OUT_N.t12 GND 0.48fF $ **FLOATING
C4077 OUT_N.t53 GND 0.48fF $ **FLOATING
C4078 OUT_N.t28 GND 0.48fF $ **FLOATING
C4079 OUT_N.t3 GND 0.48fF $ **FLOATING
C4080 OUT_N.t44 GND 0.48fF $ **FLOATING
C4081 OUT_N.t17 GND 0.48fF $ **FLOATING
C4082 OUT_N.t60 GND 0.48fF $ **FLOATING
C4083 OUT_N.t38 GND 0.48fF $ **FLOATING
C4084 OUT_N.t41 GND 3.91fF $ **FLOATING
C4085 OUT_N.n46 GND 14.21fF
C4086 OUT_N.n47 GND 12.29fF
C4087 OUT_N.n48 GND 12.29fF
C4088 OUT_N.n49 GND 12.29fF
C4089 OUT_N.n50 GND 12.29fF
C4090 OUT_N.n51 GND 12.29fF
C4091 OUT_N.n52 GND 12.29fF
C4092 OUT_N.n53 GND 12.29fF
C4093 OUT_N.n54 GND 26.86fF
C4094 OUT_N.n55 GND 46.56fF
C4095 OUT_N.n56 GND 34.52fF
C4096 OUT_N.n57 GND 34.52fF
C4097 OUT_N.n58 GND 40.64fF
C4098 OUT_N.n59 GND 40.64fF
C4099 OUT_N.n60 GND 40.63fF
C4100 OUT_N.n61 GND 41.75fF
C4101 a_50176_55366.n0 GND 0.01fF
C4102 a_50176_55366.n1 GND 0.01fF
C4103 a_50176_55366.n2 GND 0.00fF
C4104 a_50176_55366.n3 GND 0.00fF
C4105 a_50176_55366.n4 GND 0.00fF
C4106 a_50176_55366.n5 GND 0.00fF
C4107 a_50176_55366.n6 GND 0.00fF
C4108 a_50176_55366.n7 GND 0.00fF
C4109 a_50176_55366.n8 GND 0.00fF
C4110 a_50176_55366.n9 GND 0.00fF
C4111 a_50176_55366.t0 GND 0.02fF $ **FLOATING
C4112 a_50176_55366.t1 GND 0.02fF $ **FLOATING
C4113 a_50176_55366.n10 GND 0.05fF
C4114 a_50176_55366.n11 GND 0.00fF
C4115 a_50176_55366.n12 GND 0.00fF
C4116 a_50176_55366.n13 GND 0.02fF
C4117 a_50176_55366.n14 GND 0.04fF
C4118 a_50176_55366.n15 GND 0.12fF
C4119 a_50176_55366.n16 GND 0.01fF
C4120 a_50176_55366.n17 GND 0.12fF
C4121 a_50176_55366.t3 GND 3.87fF $ **FLOATING
C4122 a_50176_55366.n18 GND 0.52fF
C4123 a_50176_55366.t2 GND 0.24fF $ **FLOATING
C4124 a_50176_45486.n0 GND 0.01fF
C4125 a_50176_45486.n1 GND 0.01fF
C4126 a_50176_45486.n2 GND 0.00fF
C4127 a_50176_45486.n3 GND 0.00fF
C4128 a_50176_45486.n4 GND 0.00fF
C4129 a_50176_45486.n5 GND 0.00fF
C4130 a_50176_45486.n6 GND 0.00fF
C4131 a_50176_45486.n7 GND 0.00fF
C4132 a_50176_45486.n8 GND 0.00fF
C4133 a_50176_45486.n9 GND 0.00fF
C4134 a_50176_45486.t0 GND 0.02fF $ **FLOATING
C4135 a_50176_45486.t1 GND 0.02fF $ **FLOATING
C4136 a_50176_45486.n10 GND 0.05fF
C4137 a_50176_45486.n11 GND 0.00fF
C4138 a_50176_45486.n12 GND 0.00fF
C4139 a_50176_45486.n13 GND 0.02fF
C4140 a_50176_45486.n14 GND 0.04fF
C4141 a_50176_45486.n15 GND 0.12fF
C4142 a_50176_45486.n16 GND 0.01fF
C4143 a_50176_45486.n17 GND 0.12fF
C4144 a_50176_45486.t2 GND 3.87fF $ **FLOATING
C4145 a_50176_45486.n18 GND 0.52fF
C4146 a_50176_45486.t3 GND 0.24fF $ **FLOATING
C4147 a_50466_45562.n0 GND 0.00fF
C4148 a_50466_45562.n1 GND 0.00fF
C4149 a_50466_45562.n2 GND 0.01fF
C4150 a_50466_45562.n3 GND 0.01fF
C4151 a_50466_45562.n4 GND 0.00fF
C4152 a_50466_45562.n5 GND 0.00fF
C4153 a_50466_45562.n6 GND 0.00fF
C4154 a_50466_45562.n7 GND 0.00fF
C4155 a_50466_45562.n8 GND 0.00fF
C4156 a_50466_45562.n9 GND 0.00fF
C4157 a_50466_45562.n10 GND 0.09fF
C4158 a_50466_45562.n11 GND 0.00fF
C4159 a_50466_45562.n12 GND 0.01fF
C4160 a_50466_45562.n13 GND 0.01fF
C4161 a_50466_45562.n14 GND 0.01fF
C4162 a_50466_45562.n15 GND 0.00fF
C4163 a_50466_45562.n16 GND 0.00fF
C4164 a_50466_45562.n17 GND 0.00fF
C4165 a_50466_45562.t1 GND 0.02fF $ **FLOATING
C4166 a_50466_45562.n18 GND 0.07fF
C4167 a_50466_45562.n19 GND 0.02fF
C4168 a_50466_45562.n20 GND 0.05fF
C4169 a_50466_45562.n22 GND 0.04fF
C4170 a_50466_45562.n23 GND 0.04fF
C4171 a_50466_45562.n24 GND 0.00fF
C4172 a_50466_45562.n25 GND 0.00fF
C4173 a_50466_45562.t0 GND 0.02fF $ **FLOATING
C4174 a_50466_45562.n26 GND 0.07fF
C4175 a_50466_45562.n27 GND 0.02fF
C4176 a_50466_45562.n28 GND 0.05fF
C4177 a_50466_45562.n30 GND 0.01fF
C4178 a_50466_45562.n31 GND 0.00fF
C4179 a_50466_45562.n32 GND 0.00fF
C4180 a_50466_45562.n33 GND 0.00fF
C4181 a_50466_45562.n34 GND 0.00fF
C4182 a_50466_45562.n35 GND 0.00fF
C4183 a_50466_45562.n36 GND 0.00fF
C4184 a_50466_45562.n38 GND 0.08fF
C4185 a_50466_45562.t3 GND 4.19fF $ **FLOATING
C4186 a_50466_45562.n39 GND 0.61fF
C4187 a_50466_45562.t2 GND 0.26fF $ **FLOATING
C4188 a_n436_44966.t8 GND 0.04fF $ **FLOATING
C4189 a_n436_44966.t13 GND 0.07fF $ **FLOATING
C4190 a_n436_44966.t20 GND 0.07fF $ **FLOATING
C4191 a_n436_44966.t14 GND 0.07fF $ **FLOATING
C4192 a_n436_44966.t28 GND 0.07fF $ **FLOATING
C4193 a_n436_44966.t26 GND 0.07fF $ **FLOATING
C4194 a_n436_44966.t0 GND 0.07fF $ **FLOATING
C4195 a_n436_44966.t3 GND 0.07fF $ **FLOATING
C4196 a_n436_44966.t2 GND 0.07fF $ **FLOATING
C4197 a_n436_44966.t27 GND 0.07fF $ **FLOATING
C4198 a_n436_44966.t12 GND 0.07fF $ **FLOATING
C4199 a_n436_44966.t30 GND 0.07fF $ **FLOATING
C4200 a_n436_44966.t16 GND 0.07fF $ **FLOATING
C4201 a_n436_44966.t22 GND 0.07fF $ **FLOATING
C4202 a_n436_44966.t10 GND 0.07fF $ **FLOATING
C4203 a_n436_44966.t24 GND 0.07fF $ **FLOATING
C4204 a_n436_44966.t33 GND 0.07fF $ **FLOATING
C4205 a_n436_44966.t1 GND 0.07fF $ **FLOATING
C4206 a_n436_44966.t31 GND 0.07fF $ **FLOATING
C4207 a_n436_44966.t6 GND 0.07fF $ **FLOATING
C4208 a_n436_44966.t29 GND 0.07fF $ **FLOATING
C4209 a_n436_44966.t25 GND 0.07fF $ **FLOATING
C4210 a_n436_44966.t17 GND 0.07fF $ **FLOATING
C4211 a_n436_44966.t23 GND 0.07fF $ **FLOATING
C4212 a_n436_44966.t19 GND 0.07fF $ **FLOATING
C4213 a_n436_44966.t5 GND 0.07fF $ **FLOATING
C4214 a_n436_44966.t18 GND 0.07fF $ **FLOATING
C4215 a_n436_44966.t4 GND 0.07fF $ **FLOATING
C4216 a_n436_44966.t15 GND 0.07fF $ **FLOATING
C4217 a_n436_44966.t7 GND 0.07fF $ **FLOATING
C4218 a_n436_44966.t11 GND 0.07fF $ **FLOATING
C4219 a_n436_44966.t32 GND 0.07fF $ **FLOATING
C4220 a_n436_44966.t21 GND 0.12fF $ **FLOATING
C4221 a_n436_44966.n0 GND 20.98fF
C4222 a_n436_44966.n1 GND 10.54fF
C4223 a_n436_44966.n2 GND 10.54fF
C4224 a_n436_44966.n3 GND 10.54fF
C4225 a_n436_44966.n4 GND 10.54fF
C4226 a_n436_44966.n5 GND 10.54fF
C4227 a_n436_44966.n6 GND 10.54fF
C4228 a_n436_44966.n7 GND 10.54fF
C4229 a_n436_44966.n8 GND 10.54fF
C4230 a_n436_44966.n9 GND 10.54fF
C4231 a_n436_44966.n10 GND 10.54fF
C4232 a_n436_44966.n11 GND 10.54fF
C4233 a_n436_44966.n12 GND 10.54fF
C4234 a_n436_44966.n13 GND 10.54fF
C4235 a_n436_44966.n14 GND 28.75fF
C4236 a_n436_44966.n15 GND 28.75fF
C4237 a_n436_44966.n16 GND 10.54fF
C4238 a_n436_44966.n17 GND 10.54fF
C4239 a_n436_44966.n18 GND 10.54fF
C4240 a_n436_44966.n19 GND 10.54fF
C4241 a_n436_44966.n20 GND 10.54fF
C4242 a_n436_44966.n21 GND 10.54fF
C4243 a_n436_44966.n22 GND 10.54fF
C4244 a_n436_44966.n23 GND 10.54fF
C4245 a_n436_44966.n24 GND 10.54fF
C4246 a_n436_44966.n25 GND 10.54fF
C4247 a_n436_44966.n26 GND 10.54fF
C4248 a_n436_44966.n27 GND 10.54fF
C4249 a_n436_44966.n28 GND 10.54fF
C4250 a_n436_44966.n29 GND 10.54fF
C4251 a_n436_44966.n30 GND 11.93fF
C4252 a_n436_44966.n31 GND 0.06fF
C4253 a_n436_44966.t9 GND 0.08fF $ **FLOATING
C4254 a_68866_45562.n0 GND 0.00fF
C4255 a_68866_45562.n1 GND 0.00fF
C4256 a_68866_45562.n2 GND 0.01fF
C4257 a_68866_45562.n3 GND 0.01fF
C4258 a_68866_45562.n4 GND 0.00fF
C4259 a_68866_45562.n5 GND 0.00fF
C4260 a_68866_45562.n6 GND 0.00fF
C4261 a_68866_45562.n7 GND 0.00fF
C4262 a_68866_45562.n8 GND 0.00fF
C4263 a_68866_45562.n9 GND 0.00fF
C4264 a_68866_45562.n10 GND 0.09fF
C4265 a_68866_45562.n11 GND 0.00fF
C4266 a_68866_45562.n12 GND 0.01fF
C4267 a_68866_45562.n13 GND 0.01fF
C4268 a_68866_45562.n14 GND 0.01fF
C4269 a_68866_45562.n15 GND 0.00fF
C4270 a_68866_45562.n16 GND 0.00fF
C4271 a_68866_45562.n17 GND 0.00fF
C4272 a_68866_45562.t0 GND 0.02fF $ **FLOATING
C4273 a_68866_45562.n18 GND 0.07fF
C4274 a_68866_45562.n19 GND 0.02fF
C4275 a_68866_45562.n20 GND 0.05fF
C4276 a_68866_45562.n22 GND 0.04fF
C4277 a_68866_45562.n23 GND 0.04fF
C4278 a_68866_45562.n24 GND 0.00fF
C4279 a_68866_45562.n25 GND 0.00fF
C4280 a_68866_45562.t1 GND 0.02fF $ **FLOATING
C4281 a_68866_45562.n26 GND 0.07fF
C4282 a_68866_45562.n27 GND 0.02fF
C4283 a_68866_45562.n28 GND 0.05fF
C4284 a_68866_45562.n30 GND 0.01fF
C4285 a_68866_45562.n31 GND 0.00fF
C4286 a_68866_45562.n32 GND 0.00fF
C4287 a_68866_45562.n33 GND 0.00fF
C4288 a_68866_45562.n34 GND 0.00fF
C4289 a_68866_45562.n35 GND 0.00fF
C4290 a_68866_45562.n36 GND 0.00fF
C4291 a_68866_45562.n38 GND 0.08fF
C4292 a_68866_45562.t2 GND 4.19fF $ **FLOATING
C4293 a_68866_45562.n39 GND 0.61fF
C4294 a_68866_45562.t3 GND 0.26fF $ **FLOATING
C4295 a_31776_25726.n0 GND 0.01fF
C4296 a_31776_25726.n1 GND 0.01fF
C4297 a_31776_25726.n2 GND 0.00fF
C4298 a_31776_25726.n3 GND 0.00fF
C4299 a_31776_25726.n4 GND 0.00fF
C4300 a_31776_25726.n5 GND 0.00fF
C4301 a_31776_25726.n6 GND 0.00fF
C4302 a_31776_25726.n7 GND 0.00fF
C4303 a_31776_25726.n8 GND 0.00fF
C4304 a_31776_25726.n9 GND 0.00fF
C4305 a_31776_25726.t1 GND 0.02fF $ **FLOATING
C4306 a_31776_25726.t0 GND 0.02fF $ **FLOATING
C4307 a_31776_25726.n10 GND 0.05fF
C4308 a_31776_25726.n11 GND 0.00fF
C4309 a_31776_25726.n12 GND 0.00fF
C4310 a_31776_25726.n13 GND 0.02fF
C4311 a_31776_25726.n14 GND 0.04fF
C4312 a_31776_25726.n15 GND 0.12fF
C4313 a_31776_25726.n16 GND 0.01fF
C4314 a_31776_25726.n17 GND 0.12fF
C4315 a_31776_25726.t2 GND 3.87fF $ **FLOATING
C4316 a_31776_25726.n18 GND 0.52fF
C4317 a_31776_25726.t3 GND 0.24fF $ **FLOATING
C4318 a_n436_5446.t24 GND 0.04fF $ **FLOATING
C4319 a_n436_5446.t14 GND 0.07fF $ **FLOATING
C4320 a_n436_5446.t10 GND 0.07fF $ **FLOATING
C4321 a_n436_5446.t56 GND 0.07fF $ **FLOATING
C4322 a_n436_5446.t48 GND 0.07fF $ **FLOATING
C4323 a_n436_5446.t40 GND 0.07fF $ **FLOATING
C4324 a_n436_5446.t33 GND 0.07fF $ **FLOATING
C4325 a_n436_5446.t6 GND 0.07fF $ **FLOATING
C4326 a_n436_5446.t26 GND 0.07fF $ **FLOATING
C4327 a_n436_5446.t60 GND 0.07fF $ **FLOATING
C4328 a_n436_5446.t23 GND 0.07fF $ **FLOATING
C4329 a_n436_5446.t2 GND 0.07fF $ **FLOATING
C4330 a_n436_5446.t58 GND 0.07fF $ **FLOATING
C4331 a_n436_5446.t37 GND 0.07fF $ **FLOATING
C4332 a_n436_5446.t20 GND 0.07fF $ **FLOATING
C4333 a_n436_5446.t18 GND 0.07fF $ **FLOATING
C4334 a_n436_5446.t0 GND 0.07fF $ **FLOATING
C4335 a_n436_5446.t62 GND 0.07fF $ **FLOATING
C4336 a_n436_5446.t16 GND 0.07fF $ **FLOATING
C4337 a_n436_5446.t5 GND 0.07fF $ **FLOATING
C4338 a_n436_5446.t15 GND 0.07fF $ **FLOATING
C4339 a_n436_5446.t28 GND 0.07fF $ **FLOATING
C4340 a_n436_5446.t57 GND 0.07fF $ **FLOATING
C4341 a_n436_5446.t7 GND 0.07fF $ **FLOATING
C4342 a_n436_5446.t21 GND 0.07fF $ **FLOATING
C4343 a_n436_5446.t53 GND 0.07fF $ **FLOATING
C4344 a_n436_5446.t42 GND 0.07fF $ **FLOATING
C4345 a_n436_5446.t51 GND 0.07fF $ **FLOATING
C4346 a_n436_5446.t27 GND 0.07fF $ **FLOATING
C4347 a_n436_5446.t59 GND 0.07fF $ **FLOATING
C4348 a_n436_5446.t65 GND 0.07fF $ **FLOATING
C4349 a_n436_5446.t35 GND 0.07fF $ **FLOATING
C4350 a_n436_5446.t44 GND 0.12fF $ **FLOATING
C4351 a_n436_5446.n0 GND 21.02fF
C4352 a_n436_5446.n1 GND 10.56fF
C4353 a_n436_5446.n2 GND 10.56fF
C4354 a_n436_5446.n3 GND 10.56fF
C4355 a_n436_5446.n4 GND 10.56fF
C4356 a_n436_5446.n5 GND 10.56fF
C4357 a_n436_5446.n6 GND 10.56fF
C4358 a_n436_5446.n7 GND 10.56fF
C4359 a_n436_5446.n8 GND 10.56fF
C4360 a_n436_5446.n9 GND 10.56fF
C4361 a_n436_5446.n10 GND 10.56fF
C4362 a_n436_5446.n11 GND 10.56fF
C4363 a_n436_5446.n12 GND 10.56fF
C4364 a_n436_5446.n13 GND 10.56fF
C4365 a_n436_5446.n14 GND 19.39fF
C4366 a_n436_5446.t1 GND 0.07fF $ **FLOATING
C4367 a_n436_5446.t22 GND 0.07fF $ **FLOATING
C4368 a_n436_5446.t29 GND 0.07fF $ **FLOATING
C4369 a_n436_5446.t38 GND 0.07fF $ **FLOATING
C4370 a_n436_5446.t52 GND 0.07fF $ **FLOATING
C4371 a_n436_5446.t64 GND 0.07fF $ **FLOATING
C4372 a_n436_5446.t30 GND 0.07fF $ **FLOATING
C4373 a_n436_5446.t11 GND 0.07fF $ **FLOATING
C4374 a_n436_5446.t46 GND 0.07fF $ **FLOATING
C4375 a_n436_5446.t43 GND 0.07fF $ **FLOATING
C4376 a_n436_5446.t13 GND 0.07fF $ **FLOATING
C4377 a_n436_5446.t63 GND 0.07fF $ **FLOATING
C4378 a_n436_5446.t55 GND 0.07fF $ **FLOATING
C4379 a_n436_5446.t50 GND 0.07fF $ **FLOATING
C4380 a_n436_5446.t32 GND 0.07fF $ **FLOATING
C4381 a_n436_5446.t54 GND 0.12fF $ **FLOATING
C4382 a_n436_5446.n15 GND 21.02fF
C4383 a_n436_5446.n16 GND 10.56fF
C4384 a_n436_5446.n17 GND 10.56fF
C4385 a_n436_5446.n18 GND 10.56fF
C4386 a_n436_5446.n19 GND 10.56fF
C4387 a_n436_5446.n20 GND 10.56fF
C4388 a_n436_5446.n21 GND 10.56fF
C4389 a_n436_5446.n22 GND 10.56fF
C4390 a_n436_5446.n23 GND 10.56fF
C4391 a_n436_5446.n24 GND 10.56fF
C4392 a_n436_5446.n25 GND 10.56fF
C4393 a_n436_5446.n26 GND 10.56fF
C4394 a_n436_5446.n27 GND 10.56fF
C4395 a_n436_5446.n28 GND 10.56fF
C4396 a_n436_5446.n29 GND 9.17fF
C4397 a_n436_5446.n30 GND 38.07fF
C4398 a_n436_5446.t39 GND 0.07fF $ **FLOATING
C4399 a_n436_5446.t36 GND 0.07fF $ **FLOATING
C4400 a_n436_5446.t19 GND 0.07fF $ **FLOATING
C4401 a_n436_5446.t34 GND 0.07fF $ **FLOATING
C4402 a_n436_5446.t45 GND 0.07fF $ **FLOATING
C4403 a_n436_5446.t47 GND 0.07fF $ **FLOATING
C4404 a_n436_5446.t12 GND 0.07fF $ **FLOATING
C4405 a_n436_5446.t61 GND 0.07fF $ **FLOATING
C4406 a_n436_5446.t17 GND 0.07fF $ **FLOATING
C4407 a_n436_5446.t49 GND 0.07fF $ **FLOATING
C4408 a_n436_5446.t31 GND 0.07fF $ **FLOATING
C4409 a_n436_5446.t3 GND 0.07fF $ **FLOATING
C4410 a_n436_5446.t9 GND 0.07fF $ **FLOATING
C4411 a_n436_5446.t41 GND 0.07fF $ **FLOATING
C4412 a_n436_5446.t4 GND 0.07fF $ **FLOATING
C4413 a_n436_5446.t8 GND 0.12fF $ **FLOATING
C4414 a_n436_5446.n31 GND 21.02fF
C4415 a_n436_5446.n32 GND 10.56fF
C4416 a_n436_5446.n33 GND 10.56fF
C4417 a_n436_5446.n34 GND 10.56fF
C4418 a_n436_5446.n35 GND 10.56fF
C4419 a_n436_5446.n36 GND 10.56fF
C4420 a_n436_5446.n37 GND 10.56fF
C4421 a_n436_5446.n38 GND 10.56fF
C4422 a_n436_5446.n39 GND 10.56fF
C4423 a_n436_5446.n40 GND 10.56fF
C4424 a_n436_5446.n41 GND 10.56fF
C4425 a_n436_5446.n42 GND 10.56fF
C4426 a_n436_5446.n43 GND 10.56fF
C4427 a_n436_5446.n44 GND 10.56fF
C4428 a_n436_5446.n45 GND 9.17fF
C4429 a_n436_5446.n46 GND 38.07fF
C4430 a_n436_5446.n47 GND 19.39fF
C4431 a_n436_5446.n48 GND 10.56fF
C4432 a_n436_5446.n49 GND 10.56fF
C4433 a_n436_5446.n50 GND 10.56fF
C4434 a_n436_5446.n51 GND 10.56fF
C4435 a_n436_5446.n52 GND 10.56fF
C4436 a_n436_5446.n53 GND 10.56fF
C4437 a_n436_5446.n54 GND 10.56fF
C4438 a_n436_5446.n55 GND 10.56fF
C4439 a_n436_5446.n56 GND 10.56fF
C4440 a_n436_5446.n57 GND 10.56fF
C4441 a_n436_5446.n58 GND 10.56fF
C4442 a_n436_5446.n59 GND 10.56fF
C4443 a_n436_5446.n60 GND 10.56fF
C4444 a_n436_5446.n61 GND 10.56fF
C4445 a_n436_5446.n62 GND 11.95fF
C4446 a_n436_5446.n63 GND 0.06fF
C4447 a_n436_5446.t25 GND 0.08fF $ **FLOATING
C4448 a_4176_15846.n0 GND 0.01fF
C4449 a_4176_15846.n1 GND 0.01fF
C4450 a_4176_15846.n2 GND 0.00fF
C4451 a_4176_15846.n3 GND 0.00fF
C4452 a_4176_15846.n4 GND 0.00fF
C4453 a_4176_15846.n5 GND 0.00fF
C4454 a_4176_15846.n6 GND 0.00fF
C4455 a_4176_15846.n7 GND 0.00fF
C4456 a_4176_15846.n8 GND 0.00fF
C4457 a_4176_15846.n9 GND 0.00fF
C4458 a_4176_15846.t2 GND 0.02fF $ **FLOATING
C4459 a_4176_15846.t1 GND 0.02fF $ **FLOATING
C4460 a_4176_15846.n10 GND 0.05fF
C4461 a_4176_15846.n11 GND 0.00fF
C4462 a_4176_15846.n12 GND 0.00fF
C4463 a_4176_15846.n13 GND 0.02fF
C4464 a_4176_15846.n14 GND 0.04fF
C4465 a_4176_15846.n15 GND 0.12fF
C4466 a_4176_15846.n16 GND 0.01fF
C4467 a_4176_15846.n17 GND 0.12fF
C4468 a_4176_15846.t3 GND 3.87fF $ **FLOATING
C4469 a_4176_15846.n18 GND 0.52fF
C4470 a_4176_15846.t0 GND 0.24fF $ **FLOATING
C4471 a_13666_15922.n0 GND 0.00fF
C4472 a_13666_15922.n1 GND 0.00fF
C4473 a_13666_15922.n2 GND 0.01fF
C4474 a_13666_15922.n3 GND 0.01fF
C4475 a_13666_15922.n4 GND 0.00fF
C4476 a_13666_15922.n5 GND 0.00fF
C4477 a_13666_15922.n6 GND 0.00fF
C4478 a_13666_15922.n7 GND 0.00fF
C4479 a_13666_15922.n8 GND 0.00fF
C4480 a_13666_15922.n9 GND 0.00fF
C4481 a_13666_15922.n10 GND 0.09fF
C4482 a_13666_15922.n11 GND 0.00fF
C4483 a_13666_15922.n12 GND 0.01fF
C4484 a_13666_15922.n13 GND 0.01fF
C4485 a_13666_15922.n14 GND 0.01fF
C4486 a_13666_15922.n15 GND 0.00fF
C4487 a_13666_15922.n16 GND 0.00fF
C4488 a_13666_15922.n17 GND 0.00fF
C4489 a_13666_15922.t1 GND 0.02fF $ **FLOATING
C4490 a_13666_15922.n18 GND 0.07fF
C4491 a_13666_15922.n19 GND 0.02fF
C4492 a_13666_15922.n20 GND 0.05fF
C4493 a_13666_15922.n22 GND 0.04fF
C4494 a_13666_15922.n23 GND 0.04fF
C4495 a_13666_15922.n24 GND 0.00fF
C4496 a_13666_15922.n25 GND 0.00fF
C4497 a_13666_15922.t2 GND 0.02fF $ **FLOATING
C4498 a_13666_15922.n26 GND 0.07fF
C4499 a_13666_15922.n27 GND 0.02fF
C4500 a_13666_15922.n28 GND 0.05fF
C4501 a_13666_15922.n30 GND 0.01fF
C4502 a_13666_15922.n31 GND 0.00fF
C4503 a_13666_15922.n32 GND 0.00fF
C4504 a_13666_15922.n33 GND 0.00fF
C4505 a_13666_15922.n34 GND 0.00fF
C4506 a_13666_15922.n35 GND 0.00fF
C4507 a_13666_15922.n36 GND 0.00fF
C4508 a_13666_15922.n38 GND 0.08fF
C4509 a_13666_15922.t3 GND 4.19fF $ **FLOATING
C4510 a_13666_15922.n39 GND 0.61fF
C4511 a_13666_15922.t0 GND 0.26fF $ **FLOATING
C4512 a_13376_15846.n0 GND 0.01fF
C4513 a_13376_15846.n1 GND 0.01fF
C4514 a_13376_15846.n2 GND 0.00fF
C4515 a_13376_15846.n3 GND 0.00fF
C4516 a_13376_15846.n4 GND 0.00fF
C4517 a_13376_15846.n5 GND 0.00fF
C4518 a_13376_15846.n6 GND 0.00fF
C4519 a_13376_15846.n7 GND 0.00fF
C4520 a_13376_15846.n8 GND 0.00fF
C4521 a_13376_15846.n9 GND 0.00fF
C4522 a_13376_15846.t1 GND 0.02fF $ **FLOATING
C4523 a_13376_15846.t0 GND 0.02fF $ **FLOATING
C4524 a_13376_15846.n10 GND 0.05fF
C4525 a_13376_15846.n11 GND 0.00fF
C4526 a_13376_15846.n12 GND 0.00fF
C4527 a_13376_15846.n13 GND 0.02fF
C4528 a_13376_15846.n14 GND 0.04fF
C4529 a_13376_15846.n15 GND 0.12fF
C4530 a_13376_15846.n16 GND 0.01fF
C4531 a_13376_15846.n17 GND 0.12fF
C4532 a_13376_15846.t2 GND 3.87fF $ **FLOATING
C4533 a_13376_15846.n18 GND 0.52fF
C4534 a_13376_15846.t3 GND 0.24fF $ **FLOATING
C4535 a_4176_55366.n0 GND 0.01fF
C4536 a_4176_55366.n1 GND 0.01fF
C4537 a_4176_55366.n2 GND 0.00fF
C4538 a_4176_55366.n3 GND 0.00fF
C4539 a_4176_55366.n4 GND 0.00fF
C4540 a_4176_55366.n5 GND 0.00fF
C4541 a_4176_55366.n6 GND 0.00fF
C4542 a_4176_55366.n7 GND 0.00fF
C4543 a_4176_55366.n8 GND 0.00fF
C4544 a_4176_55366.n9 GND 0.00fF
C4545 a_4176_55366.t0 GND 0.02fF $ **FLOATING
C4546 a_4176_55366.t1 GND 0.02fF $ **FLOATING
C4547 a_4176_55366.n10 GND 0.05fF
C4548 a_4176_55366.n11 GND 0.00fF
C4549 a_4176_55366.n12 GND 0.00fF
C4550 a_4176_55366.n13 GND 0.02fF
C4551 a_4176_55366.n14 GND 0.04fF
C4552 a_4176_55366.n15 GND 0.12fF
C4553 a_4176_55366.n16 GND 0.01fF
C4554 a_4176_55366.n17 GND 0.12fF
C4555 a_4176_55366.t2 GND 3.87fF $ **FLOATING
C4556 a_4176_55366.n18 GND 0.52fF
C4557 a_4176_55366.t3 GND 0.24fF $ **FLOATING
C4558 a_n436_94366.t2 GND 0.04fF $ **FLOATING
C4559 a_n436_94366.t0 GND 0.07fF $ **FLOATING
C4560 a_n436_94366.t3 GND 0.13fF $ **FLOATING
C4561 a_n436_94366.n0 GND 23.88fF
C4562 a_n436_94366.n1 GND 0.06fF
C4563 a_n436_94366.t1 GND 0.09fF $ **FLOATING
C4564 a_4176_94886.n0 GND 0.01fF
C4565 a_4176_94886.n1 GND 0.01fF
C4566 a_4176_94886.n2 GND 0.00fF
C4567 a_4176_94886.n3 GND 0.00fF
C4568 a_4176_94886.n4 GND 0.00fF
C4569 a_4176_94886.n5 GND 0.00fF
C4570 a_4176_94886.n6 GND 0.00fF
C4571 a_4176_94886.n7 GND 0.00fF
C4572 a_4176_94886.n8 GND 0.00fF
C4573 a_4176_94886.n9 GND 0.00fF
C4574 a_4176_94886.t1 GND 0.02fF $ **FLOATING
C4575 a_4176_94886.t2 GND 0.02fF $ **FLOATING
C4576 a_4176_94886.n10 GND 0.05fF
C4577 a_4176_94886.n11 GND 0.00fF
C4578 a_4176_94886.n12 GND 0.00fF
C4579 a_4176_94886.n13 GND 0.02fF
C4580 a_4176_94886.n14 GND 0.04fF
C4581 a_4176_94886.n15 GND 0.12fF
C4582 a_4176_94886.n16 GND 0.01fF
C4583 a_4176_94886.n17 GND 0.12fF
C4584 a_4176_94886.t3 GND 3.87fF $ **FLOATING
C4585 a_4176_94886.n18 GND 0.52fF
C4586 a_4176_94886.t0 GND 0.24fF $ **FLOATING
C4587 a_50176_5966.n0 GND 0.01fF
C4588 a_50176_5966.n1 GND 0.01fF
C4589 a_50176_5966.n2 GND 0.00fF
C4590 a_50176_5966.n3 GND 0.00fF
C4591 a_50176_5966.n4 GND 0.00fF
C4592 a_50176_5966.n5 GND 0.00fF
C4593 a_50176_5966.n6 GND 0.00fF
C4594 a_50176_5966.n7 GND 0.00fF
C4595 a_50176_5966.n8 GND 0.00fF
C4596 a_50176_5966.n9 GND 0.00fF
C4597 a_50176_5966.t1 GND 0.02fF $ **FLOATING
C4598 a_50176_5966.t2 GND 0.02fF $ **FLOATING
C4599 a_50176_5966.n10 GND 0.05fF
C4600 a_50176_5966.n11 GND 0.00fF
C4601 a_50176_5966.n12 GND 0.00fF
C4602 a_50176_5966.n13 GND 0.02fF
C4603 a_50176_5966.n14 GND 0.04fF
C4604 a_50176_5966.n15 GND 0.12fF
C4605 a_50176_5966.n16 GND 0.01fF
C4606 a_50176_5966.n17 GND 0.12fF
C4607 a_50176_5966.t3 GND 3.87fF $ **FLOATING
C4608 a_50176_5966.n18 GND 0.52fF
C4609 a_50176_5966.t0 GND 0.24fF $ **FLOATING
C4610 a_50466_6042.n0 GND 0.00fF
C4611 a_50466_6042.n1 GND 0.00fF
C4612 a_50466_6042.n2 GND 0.01fF
C4613 a_50466_6042.n3 GND 0.01fF
C4614 a_50466_6042.n4 GND 0.00fF
C4615 a_50466_6042.n5 GND 0.00fF
C4616 a_50466_6042.n6 GND 0.00fF
C4617 a_50466_6042.n7 GND 0.00fF
C4618 a_50466_6042.n8 GND 0.00fF
C4619 a_50466_6042.n9 GND 0.00fF
C4620 a_50466_6042.n10 GND 0.09fF
C4621 a_50466_6042.n11 GND 0.00fF
C4622 a_50466_6042.n12 GND 0.01fF
C4623 a_50466_6042.n13 GND 0.01fF
C4624 a_50466_6042.n14 GND 0.01fF
C4625 a_50466_6042.n15 GND 0.00fF
C4626 a_50466_6042.n16 GND 0.00fF
C4627 a_50466_6042.n17 GND 0.00fF
C4628 a_50466_6042.t1 GND 0.02fF $ **FLOATING
C4629 a_50466_6042.n18 GND 0.07fF
C4630 a_50466_6042.n19 GND 0.02fF
C4631 a_50466_6042.n20 GND 0.05fF
C4632 a_50466_6042.n22 GND 0.04fF
C4633 a_50466_6042.n23 GND 0.04fF
C4634 a_50466_6042.n24 GND 0.00fF
C4635 a_50466_6042.n25 GND 0.00fF
C4636 a_50466_6042.t0 GND 0.02fF $ **FLOATING
C4637 a_50466_6042.n26 GND 0.07fF
C4638 a_50466_6042.n27 GND 0.02fF
C4639 a_50466_6042.n28 GND 0.05fF
C4640 a_50466_6042.n30 GND 0.01fF
C4641 a_50466_6042.n31 GND 0.00fF
C4642 a_50466_6042.n32 GND 0.00fF
C4643 a_50466_6042.n33 GND 0.00fF
C4644 a_50466_6042.n34 GND 0.00fF
C4645 a_50466_6042.n35 GND 0.00fF
C4646 a_50466_6042.n36 GND 0.00fF
C4647 a_50466_6042.n38 GND 0.08fF
C4648 a_50466_6042.t2 GND 4.19fF $ **FLOATING
C4649 a_50466_6042.n39 GND 0.61fF
C4650 a_50466_6042.t3 GND 0.26fF $ **FLOATING
C4651 bit5.t43 GND 0.03fF $ **FLOATING
C4652 bit5.n0 GND 0.01fF
C4653 bit5.n1 GND 0.00fF
C4654 bit5.t5 GND 0.03fF $ **FLOATING
C4655 bit5.n2 GND 0.01fF
C4656 bit5.n3 GND 0.00fF
C4657 bit5.n4 GND 0.00fF
C4658 bit5.n5 GND 0.00fF
C4659 bit5.n6 GND 0.07fF
C4660 bit5.t40 GND 0.03fF $ **FLOATING
C4661 bit5.n7 GND 0.01fF
C4662 bit5.n8 GND 0.00fF
C4663 bit5.t12 GND 0.03fF $ **FLOATING
C4664 bit5.n9 GND 0.01fF
C4665 bit5.n10 GND 0.00fF
C4666 bit5.n11 GND 0.00fF
C4667 bit5.n12 GND 0.00fF
C4668 bit5.n13 GND 0.07fF
C4669 bit5.t61 GND 0.03fF $ **FLOATING
C4670 bit5.n14 GND 0.01fF
C4671 bit5.n15 GND 0.00fF
C4672 bit5.t37 GND 0.03fF $ **FLOATING
C4673 bit5.n16 GND 0.01fF
C4674 bit5.n17 GND 0.00fF
C4675 bit5.n18 GND 0.00fF
C4676 bit5.n19 GND 0.00fF
C4677 bit5.n20 GND 0.07fF
C4678 bit5.t59 GND 0.03fF $ **FLOATING
C4679 bit5.n21 GND 0.01fF
C4680 bit5.n22 GND 0.00fF
C4681 bit5.t33 GND 0.03fF $ **FLOATING
C4682 bit5.n23 GND 0.01fF
C4683 bit5.n24 GND 0.00fF
C4684 bit5.n25 GND 0.00fF
C4685 bit5.n26 GND 0.00fF
C4686 bit5.n27 GND 0.07fF
C4687 bit5.t55 GND 0.03fF $ **FLOATING
C4688 bit5.n28 GND 0.01fF
C4689 bit5.n29 GND 0.00fF
C4690 bit5.t28 GND 0.03fF $ **FLOATING
C4691 bit5.n30 GND 0.01fF
C4692 bit5.n31 GND 0.00fF
C4693 bit5.n32 GND 0.00fF
C4694 bit5.n33 GND 0.00fF
C4695 bit5.n34 GND 0.07fF
C4696 bit5.t60 GND 0.03fF $ **FLOATING
C4697 bit5.n35 GND 0.01fF
C4698 bit5.n36 GND 0.00fF
C4699 bit5.t24 GND 0.03fF $ **FLOATING
C4700 bit5.n37 GND 0.01fF
C4701 bit5.n38 GND 0.00fF
C4702 bit5.n39 GND 0.00fF
C4703 bit5.n40 GND 0.00fF
C4704 bit5.n41 GND 0.07fF
C4705 bit5.t58 GND 0.03fF $ **FLOATING
C4706 bit5.n42 GND 0.01fF
C4707 bit5.n43 GND 0.00fF
C4708 bit5.t31 GND 0.03fF $ **FLOATING
C4709 bit5.n44 GND 0.01fF
C4710 bit5.n45 GND 0.00fF
C4711 bit5.n46 GND 0.00fF
C4712 bit5.n47 GND 0.00fF
C4713 bit5.n48 GND 0.07fF
C4714 bit5.n49 GND 0.00fF
C4715 bit5.n50 GND 0.00fF
C4716 bit5.t3 GND 0.03fF $ **FLOATING
C4717 bit5.n51 GND 0.01fF
C4718 bit5.n52 GND 0.00fF
C4719 bit5.t46 GND 0.03fF $ **FLOATING
C4720 bit5.n53 GND 0.01fF
C4721 bit5.n54 GND 0.00fF
C4722 bit5.n55 GND 11.99fF
C4723 bit5.n56 GND 24.30fF
C4724 bit5.n57 GND 18.13fF
C4725 bit5.n58 GND 18.13fF
C4726 bit5.n59 GND 18.13fF
C4727 bit5.n60 GND 18.13fF
C4728 bit5.n61 GND 18.13fF
C4729 bit5.n62 GND 29.05fF
C4730 bit5.t18 GND 0.03fF $ **FLOATING
C4731 bit5.n63 GND 0.01fF
C4732 bit5.n64 GND 0.00fF
C4733 bit5.t52 GND 0.03fF $ **FLOATING
C4734 bit5.n65 GND 0.01fF
C4735 bit5.n66 GND 0.00fF
C4736 bit5.n67 GND 0.00fF
C4737 bit5.n68 GND 0.00fF
C4738 bit5.n69 GND 0.07fF
C4739 bit5.t16 GND 0.03fF $ **FLOATING
C4740 bit5.n70 GND 0.01fF
C4741 bit5.n71 GND 0.00fF
C4742 bit5.t53 GND 0.03fF $ **FLOATING
C4743 bit5.n72 GND 0.01fF
C4744 bit5.n73 GND 0.00fF
C4745 bit5.n74 GND 0.00fF
C4746 bit5.n75 GND 0.00fF
C4747 bit5.n76 GND 0.07fF
C4748 bit5.t42 GND 0.03fF $ **FLOATING
C4749 bit5.n77 GND 0.01fF
C4750 bit5.n78 GND 0.00fF
C4751 bit5.t15 GND 0.03fF $ **FLOATING
C4752 bit5.n79 GND 0.01fF
C4753 bit5.n80 GND 0.00fF
C4754 bit5.n81 GND 0.00fF
C4755 bit5.n82 GND 0.00fF
C4756 bit5.n83 GND 0.07fF
C4757 bit5.t39 GND 0.03fF $ **FLOATING
C4758 bit5.n84 GND 0.01fF
C4759 bit5.n85 GND 0.00fF
C4760 bit5.t11 GND 0.03fF $ **FLOATING
C4761 bit5.n86 GND 0.01fF
C4762 bit5.n87 GND 0.00fF
C4763 bit5.n88 GND 0.00fF
C4764 bit5.n89 GND 0.00fF
C4765 bit5.n90 GND 0.07fF
C4766 bit5.t35 GND 0.03fF $ **FLOATING
C4767 bit5.n91 GND 0.01fF
C4768 bit5.n92 GND 0.00fF
C4769 bit5.t8 GND 0.03fF $ **FLOATING
C4770 bit5.n93 GND 0.01fF
C4771 bit5.n94 GND 0.00fF
C4772 bit5.n95 GND 0.00fF
C4773 bit5.n96 GND 0.00fF
C4774 bit5.n97 GND 0.07fF
C4775 bit5.t41 GND 0.03fF $ **FLOATING
C4776 bit5.n98 GND 0.01fF
C4777 bit5.n99 GND 0.00fF
C4778 bit5.t4 GND 0.03fF $ **FLOATING
C4779 bit5.n100 GND 0.01fF
C4780 bit5.n101 GND 0.00fF
C4781 bit5.n102 GND 0.00fF
C4782 bit5.n103 GND 0.00fF
C4783 bit5.n104 GND 0.07fF
C4784 bit5.t36 GND 0.03fF $ **FLOATING
C4785 bit5.n105 GND 0.01fF
C4786 bit5.n106 GND 0.00fF
C4787 bit5.t10 GND 0.03fF $ **FLOATING
C4788 bit5.n107 GND 0.01fF
C4789 bit5.n108 GND 0.00fF
C4790 bit5.n109 GND 0.00fF
C4791 bit5.n110 GND 0.00fF
C4792 bit5.n111 GND 0.07fF
C4793 bit5.t50 GND 0.03fF $ **FLOATING
C4794 bit5.n112 GND 0.01fF
C4795 bit5.n113 GND 0.00fF
C4796 bit5.t21 GND 0.03fF $ **FLOATING
C4797 bit5.n114 GND 0.01fF
C4798 bit5.n115 GND 0.00fF
C4799 bit5.n116 GND 0.00fF
C4800 bit5.n117 GND 0.00fF
C4801 bit5.n118 GND 11.99fF
C4802 bit5.n119 GND 24.30fF
C4803 bit5.n120 GND 18.13fF
C4804 bit5.n121 GND 18.13fF
C4805 bit5.n122 GND 18.13fF
C4806 bit5.n123 GND 18.13fF
C4807 bit5.n124 GND 18.13fF
C4808 bit5.n125 GND 20.51fF
C4809 bit5.n126 GND 41.49fF
C4810 bit5.t13 GND 0.03fF $ **FLOATING
C4811 bit5.n127 GND 0.01fF
C4812 bit5.n128 GND 0.00fF
C4813 bit5.t45 GND 0.03fF $ **FLOATING
C4814 bit5.n129 GND 0.01fF
C4815 bit5.n130 GND 0.00fF
C4816 bit5.n131 GND 0.00fF
C4817 bit5.n132 GND 0.00fF
C4818 bit5.n133 GND 0.07fF
C4819 bit5.t9 GND 0.03fF $ **FLOATING
C4820 bit5.n134 GND 0.01fF
C4821 bit5.n135 GND 0.00fF
C4822 bit5.t49 GND 0.03fF $ **FLOATING
C4823 bit5.n136 GND 0.01fF
C4824 bit5.n137 GND 0.00fF
C4825 bit5.n138 GND 0.00fF
C4826 bit5.n139 GND 0.00fF
C4827 bit5.n140 GND 0.07fF
C4828 bit5.t34 GND 0.03fF $ **FLOATING
C4829 bit5.n141 GND 0.01fF
C4830 bit5.n142 GND 0.00fF
C4831 bit5.t6 GND 0.03fF $ **FLOATING
C4832 bit5.n143 GND 0.01fF
C4833 bit5.n144 GND 0.00fF
C4834 bit5.n145 GND 0.00fF
C4835 bit5.n146 GND 0.00fF
C4836 bit5.n147 GND 0.07fF
C4837 bit5.t29 GND 0.03fF $ **FLOATING
C4838 bit5.n148 GND 0.01fF
C4839 bit5.n149 GND 0.00fF
C4840 bit5.t2 GND 0.03fF $ **FLOATING
C4841 bit5.n150 GND 0.01fF
C4842 bit5.n151 GND 0.00fF
C4843 bit5.n152 GND 0.00fF
C4844 bit5.n153 GND 0.00fF
C4845 bit5.n154 GND 0.07fF
C4846 bit5.t25 GND 0.03fF $ **FLOATING
C4847 bit5.n155 GND 0.01fF
C4848 bit5.n156 GND 0.00fF
C4849 bit5.t64 GND 0.03fF $ **FLOATING
C4850 bit5.n157 GND 0.01fF
C4851 bit5.n158 GND 0.00fF
C4852 bit5.n159 GND 0.00fF
C4853 bit5.n160 GND 0.00fF
C4854 bit5.n161 GND 0.07fF
C4855 bit5.t32 GND 0.03fF $ **FLOATING
C4856 bit5.n162 GND 0.01fF
C4857 bit5.n163 GND 0.00fF
C4858 bit5.t63 GND 0.03fF $ **FLOATING
C4859 bit5.n164 GND 0.01fF
C4860 bit5.n165 GND 0.00fF
C4861 bit5.n166 GND 0.00fF
C4862 bit5.n167 GND 0.00fF
C4863 bit5.n168 GND 0.07fF
C4864 bit5.t26 GND 0.03fF $ **FLOATING
C4865 bit5.n169 GND 0.01fF
C4866 bit5.n170 GND 0.00fF
C4867 bit5.t1 GND 0.03fF $ **FLOATING
C4868 bit5.n171 GND 0.01fF
C4869 bit5.n172 GND 0.00fF
C4870 bit5.n173 GND 0.00fF
C4871 bit5.n174 GND 0.00fF
C4872 bit5.n175 GND 0.07fF
C4873 bit5.t44 GND 0.03fF $ **FLOATING
C4874 bit5.n176 GND 0.01fF
C4875 bit5.n177 GND 0.00fF
C4876 bit5.t17 GND 0.03fF $ **FLOATING
C4877 bit5.n178 GND 0.01fF
C4878 bit5.n179 GND 0.00fF
C4879 bit5.n180 GND 0.00fF
C4880 bit5.n181 GND 0.00fF
C4881 bit5.n182 GND 11.99fF
C4882 bit5.n183 GND 24.30fF
C4883 bit5.n184 GND 18.13fF
C4884 bit5.n185 GND 18.13fF
C4885 bit5.n186 GND 18.13fF
C4886 bit5.n187 GND 18.13fF
C4887 bit5.n188 GND 18.13fF
C4888 bit5.n189 GND 20.51fF
C4889 bit5.n190 GND 28.89fF
C4890 bit5.t20 GND 0.03fF $ **FLOATING
C4891 bit5.n191 GND 0.01fF
C4892 bit5.n192 GND 0.00fF
C4893 bit5.t30 GND 0.03fF $ **FLOATING
C4894 bit5.n193 GND 0.01fF
C4895 bit5.n194 GND 0.00fF
C4896 bit5.n195 GND 0.00fF
C4897 bit5.n196 GND 0.00fF
C4898 bit5.n197 GND 0.07fF
C4899 bit5.t51 GND 0.03fF $ **FLOATING
C4900 bit5.n198 GND 0.01fF
C4901 bit5.n199 GND 0.00fF
C4902 bit5.t38 GND 0.03fF $ **FLOATING
C4903 bit5.n200 GND 0.01fF
C4904 bit5.n201 GND 0.00fF
C4905 bit5.n202 GND 0.00fF
C4906 bit5.n203 GND 0.00fF
C4907 bit5.n204 GND 0.07fF
C4908 bit5.t0 GND 0.03fF $ **FLOATING
C4909 bit5.n205 GND 0.01fF
C4910 bit5.n206 GND 0.00fF
C4911 bit5.t54 GND 0.03fF $ **FLOATING
C4912 bit5.n207 GND 0.01fF
C4913 bit5.n208 GND 0.00fF
C4914 bit5.n209 GND 0.00fF
C4915 bit5.n210 GND 0.00fF
C4916 bit5.n211 GND 0.07fF
C4917 bit5.t27 GND 0.03fF $ **FLOATING
C4918 bit5.n212 GND 0.01fF
C4919 bit5.n213 GND 0.00fF
C4920 bit5.t19 GND 0.03fF $ **FLOATING
C4921 bit5.n214 GND 0.01fF
C4922 bit5.n215 GND 0.00fF
C4923 bit5.n216 GND 0.00fF
C4924 bit5.n217 GND 0.00fF
C4925 bit5.n218 GND 0.07fF
C4926 bit5.t57 GND 0.03fF $ **FLOATING
C4927 bit5.n219 GND 0.01fF
C4928 bit5.n220 GND 0.00fF
C4929 bit5.t48 GND 0.03fF $ **FLOATING
C4930 bit5.n221 GND 0.01fF
C4931 bit5.n222 GND 0.00fF
C4932 bit5.n223 GND 0.00fF
C4933 bit5.n224 GND 0.00fF
C4934 bit5.n225 GND 0.07fF
C4935 bit5.t62 GND 0.03fF $ **FLOATING
C4936 bit5.n226 GND 0.01fF
C4937 bit5.n227 GND 0.00fF
C4938 bit5.t7 GND 0.03fF $ **FLOATING
C4939 bit5.n228 GND 0.01fF
C4940 bit5.n229 GND 0.00fF
C4941 bit5.n230 GND 0.00fF
C4942 bit5.n231 GND 0.00fF
C4943 bit5.n232 GND 0.07fF
C4944 bit5.t22 GND 0.03fF $ **FLOATING
C4945 bit5.n233 GND 0.01fF
C4946 bit5.n234 GND 0.00fF
C4947 bit5.t14 GND 0.03fF $ **FLOATING
C4948 bit5.n235 GND 0.01fF
C4949 bit5.n236 GND 0.00fF
C4950 bit5.n237 GND 0.00fF
C4951 bit5.n238 GND 0.00fF
C4952 bit5.n239 GND 0.07fF
C4953 bit5.t56 GND 0.03fF $ **FLOATING
C4954 bit5.n240 GND 0.01fF
C4955 bit5.n241 GND 0.00fF
C4956 bit5.t47 GND 0.03fF $ **FLOATING
C4957 bit5.n242 GND 0.01fF
C4958 bit5.n243 GND 0.00fF
C4959 bit5.n244 GND 0.00fF
C4960 bit5.n245 GND 0.00fF
C4961 bit5.n246 GND 0.07fF
C4962 bit5.t65 GND 0.01fF $ **FLOATING
C4963 bit5.t23 GND 0.01fF $ **FLOATING
C4964 bit5.n247 GND 0.03fF
C4965 bit5.n248 GND 18.47fF
C4966 bit5.n249 GND 18.13fF
C4967 bit5.n250 GND 18.13fF
C4968 bit5.n251 GND 18.13fF
C4969 bit5.n252 GND 18.13fF
C4970 bit5.n253 GND 18.13fF
C4971 bit5.n254 GND 18.13fF
C4972 bit5.n255 GND 20.51fF
C4973 bit5.n256 GND 21.14fF
C4974 a_59376_45486.n0 GND 0.01fF
C4975 a_59376_45486.n1 GND 0.01fF
C4976 a_59376_45486.n2 GND 0.00fF
C4977 a_59376_45486.n3 GND 0.00fF
C4978 a_59376_45486.n4 GND 0.00fF
C4979 a_59376_45486.n5 GND 0.00fF
C4980 a_59376_45486.n6 GND 0.00fF
C4981 a_59376_45486.n7 GND 0.00fF
C4982 a_59376_45486.n8 GND 0.00fF
C4983 a_59376_45486.n9 GND 0.00fF
C4984 a_59376_45486.t1 GND 0.02fF $ **FLOATING
C4985 a_59376_45486.t0 GND 0.02fF $ **FLOATING
C4986 a_59376_45486.n10 GND 0.05fF
C4987 a_59376_45486.n11 GND 0.00fF
C4988 a_59376_45486.n12 GND 0.00fF
C4989 a_59376_45486.n13 GND 0.02fF
C4990 a_59376_45486.n14 GND 0.04fF
C4991 a_59376_45486.n15 GND 0.12fF
C4992 a_59376_45486.n16 GND 0.01fF
C4993 a_59376_45486.n17 GND 0.12fF
C4994 a_59376_45486.t2 GND 3.87fF $ **FLOATING
C4995 a_59376_45486.n18 GND 0.52fF
C4996 a_59376_45486.t3 GND 0.24fF $ **FLOATING
C4997 OUT_P.t2 GND 0.46fF $ **FLOATING
C4998 OUT_P.t9 GND 0.46fF $ **FLOATING
C4999 OUT_P.t52 GND 0.13fF $ **FLOATING
C5000 OUT_P.t26 GND 0.13fF $ **FLOATING
C5001 OUT_P.t1 GND 0.13fF $ **FLOATING
C5002 OUT_P.t40 GND 0.13fF $ **FLOATING
C5003 OUT_P.t15 GND 0.13fF $ **FLOATING
C5004 OUT_P.t58 GND 0.13fF $ **FLOATING
C5005 OUT_P.t32 GND 0.13fF $ **FLOATING
C5006 OUT_P.t48 GND 6.80fF $ **FLOATING
C5007 OUT_P.n0 GND 18.86fF
C5008 OUT_P.n1 GND 11.90fF
C5009 OUT_P.n2 GND 11.90fF
C5010 OUT_P.n3 GND 11.90fF
C5011 OUT_P.n4 GND 11.90fF
C5012 OUT_P.n5 GND 11.90fF
C5013 OUT_P.n6 GND 11.90fF
C5014 OUT_P.n7 GND 11.90fF
C5015 OUT_P.n8 GND 10.46fF
C5016 OUT_P.t51 GND 0.46fF $ **FLOATING
C5017 OUT_P.t31 GND 0.46fF $ **FLOATING
C5018 OUT_P.t6 GND 0.13fF $ **FLOATING
C5019 OUT_P.t46 GND 0.13fF $ **FLOATING
C5020 OUT_P.t21 GND 0.13fF $ **FLOATING
C5021 OUT_P.t57 GND 0.13fF $ **FLOATING
C5022 OUT_P.t35 GND 0.13fF $ **FLOATING
C5023 OUT_P.t8 GND 0.13fF $ **FLOATING
C5024 OUT_P.t36 GND 6.80fF $ **FLOATING
C5025 OUT_P.n9 GND 18.86fF
C5026 OUT_P.n10 GND 11.90fF
C5027 OUT_P.n11 GND 11.90fF
C5028 OUT_P.n12 GND 11.90fF
C5029 OUT_P.n13 GND 11.90fF
C5030 OUT_P.n14 GND 11.90fF
C5031 OUT_P.n15 GND 11.90fF
C5032 OUT_P.n16 GND 16.40fF
C5033 OUT_P.t55 GND 0.46fF $ **FLOATING
C5034 OUT_P.t30 GND 0.13fF $ **FLOATING
C5035 OUT_P.t5 GND 0.13fF $ **FLOATING
C5036 OUT_P.t45 GND 0.13fF $ **FLOATING
C5037 OUT_P.t18 GND 0.13fF $ **FLOATING
C5038 OUT_P.t61 GND 0.13fF $ **FLOATING
C5039 OUT_P.t34 GND 0.13fF $ **FLOATING
C5040 OUT_P.t37 GND 6.80fF $ **FLOATING
C5041 OUT_P.n17 GND 18.86fF
C5042 OUT_P.n18 GND 11.90fF
C5043 OUT_P.n19 GND 11.90fF
C5044 OUT_P.n20 GND 11.90fF
C5045 OUT_P.n21 GND 11.90fF
C5046 OUT_P.n22 GND 11.90fF
C5047 OUT_P.n23 GND 22.35fF
C5048 OUT_P.t14 GND 0.46fF $ **FLOATING
C5049 OUT_P.t54 GND 0.46fF $ **FLOATING
C5050 OUT_P.t29 GND 0.13fF $ **FLOATING
C5051 OUT_P.t4 GND 0.13fF $ **FLOATING
C5052 OUT_P.t43 GND 0.13fF $ **FLOATING
C5053 OUT_P.t23 GND 0.13fF $ **FLOATING
C5054 OUT_P.t60 GND 0.13fF $ **FLOATING
C5055 OUT_P.t42 GND 6.80fF $ **FLOATING
C5056 OUT_P.n24 GND 18.86fF
C5057 OUT_P.n25 GND 11.90fF
C5058 OUT_P.n26 GND 11.90fF
C5059 OUT_P.n27 GND 11.90fF
C5060 OUT_P.n28 GND 11.90fF
C5061 OUT_P.n29 GND 11.90fF
C5062 OUT_P.n30 GND 22.35fF
C5063 OUT_P.t38 GND 0.46fF $ **FLOATING
C5064 OUT_P.t12 GND 0.13fF $ **FLOATING
C5065 OUT_P.t53 GND 0.13fF $ **FLOATING
C5066 OUT_P.t27 GND 0.13fF $ **FLOATING
C5067 OUT_P.t7 GND 0.13fF $ **FLOATING
C5068 OUT_P.t47 GND 0.13fF $ **FLOATING
C5069 OUT_P.t17 GND 6.80fF $ **FLOATING
C5070 OUT_P.n31 GND 18.86fF
C5071 OUT_P.n32 GND 11.90fF
C5072 OUT_P.n33 GND 11.90fF
C5073 OUT_P.n34 GND 11.90fF
C5074 OUT_P.n35 GND 11.90fF
C5075 OUT_P.n36 GND 28.29fF
C5076 OUT_P.t28 GND 0.46fF $ **FLOATING
C5077 OUT_P.t3 GND 0.13fF $ **FLOATING
C5078 OUT_P.t41 GND 0.13fF $ **FLOATING
C5079 OUT_P.t16 GND 0.13fF $ **FLOATING
C5080 OUT_P.t59 GND 0.13fF $ **FLOATING
C5081 OUT_P.t33 GND 0.13fF $ **FLOATING
C5082 OUT_P.t10 GND 6.80fF $ **FLOATING
C5083 OUT_P.n37 GND 18.86fF
C5084 OUT_P.n38 GND 11.90fF
C5085 OUT_P.n39 GND 11.90fF
C5086 OUT_P.n40 GND 11.90fF
C5087 OUT_P.n41 GND 11.90fF
C5088 OUT_P.n42 GND 28.29fF
C5089 OUT_P.t50 GND 0.46fF $ **FLOATING
C5090 OUT_P.t25 GND 0.13fF $ **FLOATING
C5091 OUT_P.t0 GND 0.13fF $ **FLOATING
C5092 OUT_P.t39 GND 0.13fF $ **FLOATING
C5093 OUT_P.t22 GND 0.13fF $ **FLOATING
C5094 OUT_P.t56 GND 0.13fF $ **FLOATING
C5095 OUT_P.t13 GND 6.80fF $ **FLOATING
C5096 OUT_P.n43 GND 18.86fF
C5097 OUT_P.n44 GND 11.90fF
C5098 OUT_P.n45 GND 11.90fF
C5099 OUT_P.n46 GND 11.90fF
C5100 OUT_P.n47 GND 11.90fF
C5101 OUT_P.n48 GND 28.29fF
C5102 OUT_P.t11 GND 0.46fF $ **FLOATING
C5103 OUT_P.t49 GND 0.46fF $ **FLOATING
C5104 OUT_P.t24 GND 0.46fF $ **FLOATING
C5105 OUT_P.t62 GND 0.46fF $ **FLOATING
C5106 OUT_P.t44 GND 0.46fF $ **FLOATING
C5107 OUT_P.t19 GND 0.46fF $ **FLOATING
C5108 OUT_P.t20 GND 9.25fF $ **FLOATING
C5109 OUT_P.n49 GND 16.75fF
C5110 OUT_P.n50 GND 11.90fF
C5111 OUT_P.n51 GND 11.90fF
C5112 OUT_P.n52 GND 11.90fF
C5113 OUT_P.n53 GND 11.90fF
C5114 OUT_P.n54 GND 34.82fF
C5115 OUT_P.n55 GND 69.40fF
C5116 OUT_P.n56 GND 43.01fF
C5117 OUT_P.n57 GND 43.01fF
C5118 OUT_P.n58 GND 37.07fF
C5119 OUT_P.n59 GND 37.07fF
C5120 OUT_P.n60 GND 31.13fF
C5121 OUT_P.n61 GND 26.73fF
C5122 a_22576_45486.n0 GND 0.01fF
C5123 a_22576_45486.n1 GND 0.01fF
C5124 a_22576_45486.n2 GND 0.00fF
C5125 a_22576_45486.n3 GND 0.00fF
C5126 a_22576_45486.n4 GND 0.00fF
C5127 a_22576_45486.n5 GND 0.00fF
C5128 a_22576_45486.n6 GND 0.00fF
C5129 a_22576_45486.n7 GND 0.00fF
C5130 a_22576_45486.n8 GND 0.00fF
C5131 a_22576_45486.n9 GND 0.00fF
C5132 a_22576_45486.t0 GND 0.02fF $ **FLOATING
C5133 a_22576_45486.t1 GND 0.02fF $ **FLOATING
C5134 a_22576_45486.n10 GND 0.05fF
C5135 a_22576_45486.n11 GND 0.00fF
C5136 a_22576_45486.n12 GND 0.00fF
C5137 a_22576_45486.n13 GND 0.02fF
C5138 a_22576_45486.n14 GND 0.04fF
C5139 a_22576_45486.n15 GND 0.12fF
C5140 a_22576_45486.n16 GND 0.01fF
C5141 a_22576_45486.n17 GND 0.12fF
C5142 a_22576_45486.t2 GND 3.87fF $ **FLOATING
C5143 a_22576_45486.n18 GND 0.52fF
C5144 a_22576_45486.t3 GND 0.24fF $ **FLOATING
C5145 a_22866_45562.n0 GND 0.00fF
C5146 a_22866_45562.n1 GND 0.00fF
C5147 a_22866_45562.n2 GND 0.01fF
C5148 a_22866_45562.n3 GND 0.01fF
C5149 a_22866_45562.n4 GND 0.00fF
C5150 a_22866_45562.n5 GND 0.00fF
C5151 a_22866_45562.n6 GND 0.00fF
C5152 a_22866_45562.n7 GND 0.00fF
C5153 a_22866_45562.n8 GND 0.00fF
C5154 a_22866_45562.n9 GND 0.00fF
C5155 a_22866_45562.n10 GND 0.09fF
C5156 a_22866_45562.n11 GND 0.00fF
C5157 a_22866_45562.n12 GND 0.01fF
C5158 a_22866_45562.n13 GND 0.01fF
C5159 a_22866_45562.n14 GND 0.01fF
C5160 a_22866_45562.n15 GND 0.00fF
C5161 a_22866_45562.n16 GND 0.00fF
C5162 a_22866_45562.n17 GND 0.00fF
C5163 a_22866_45562.t2 GND 0.02fF $ **FLOATING
C5164 a_22866_45562.n18 GND 0.07fF
C5165 a_22866_45562.n19 GND 0.02fF
C5166 a_22866_45562.n20 GND 0.05fF
C5167 a_22866_45562.n22 GND 0.04fF
C5168 a_22866_45562.n23 GND 0.04fF
C5169 a_22866_45562.n24 GND 0.00fF
C5170 a_22866_45562.n25 GND 0.00fF
C5171 a_22866_45562.t1 GND 0.02fF $ **FLOATING
C5172 a_22866_45562.n26 GND 0.07fF
C5173 a_22866_45562.n27 GND 0.02fF
C5174 a_22866_45562.n28 GND 0.05fF
C5175 a_22866_45562.n30 GND 0.01fF
C5176 a_22866_45562.n31 GND 0.00fF
C5177 a_22866_45562.n32 GND 0.00fF
C5178 a_22866_45562.n33 GND 0.00fF
C5179 a_22866_45562.n34 GND 0.00fF
C5180 a_22866_45562.n35 GND 0.00fF
C5181 a_22866_45562.n36 GND 0.00fF
C5182 a_22866_45562.n38 GND 0.08fF
C5183 a_22866_45562.t3 GND 4.19fF $ **FLOATING
C5184 a_22866_45562.n39 GND 0.61fF
C5185 a_22866_45562.t0 GND 0.26fF $ **FLOATING
C5186 bit4.t28 GND 0.03fF $ **FLOATING
C5187 bit4.n0 GND 0.01fF
C5188 bit4.n1 GND 0.00fF
C5189 bit4.t11 GND 0.03fF $ **FLOATING
C5190 bit4.n2 GND 0.01fF
C5191 bit4.n3 GND 0.00fF
C5192 bit4.n4 GND 0.00fF
C5193 bit4.n5 GND 0.00fF
C5194 bit4.n6 GND 0.07fF
C5195 bit4.t26 GND 0.03fF $ **FLOATING
C5196 bit4.n7 GND 0.01fF
C5197 bit4.n8 GND 0.00fF
C5198 bit4.t12 GND 0.03fF $ **FLOATING
C5199 bit4.n9 GND 0.01fF
C5200 bit4.n10 GND 0.00fF
C5201 bit4.n11 GND 0.00fF
C5202 bit4.n12 GND 0.00fF
C5203 bit4.n13 GND 0.07fF
C5204 bit4.t6 GND 0.03fF $ **FLOATING
C5205 bit4.n14 GND 0.01fF
C5206 bit4.n15 GND 0.00fF
C5207 bit4.t25 GND 0.03fF $ **FLOATING
C5208 bit4.n16 GND 0.01fF
C5209 bit4.n17 GND 0.00fF
C5210 bit4.n18 GND 0.00fF
C5211 bit4.n19 GND 0.00fF
C5212 bit4.n20 GND 0.07fF
C5213 bit4.t4 GND 0.03fF $ **FLOATING
C5214 bit4.n21 GND 0.01fF
C5215 bit4.n22 GND 0.00fF
C5216 bit4.t23 GND 0.03fF $ **FLOATING
C5217 bit4.n23 GND 0.01fF
C5218 bit4.n24 GND 0.00fF
C5219 bit4.n25 GND 0.00fF
C5220 bit4.n26 GND 0.00fF
C5221 bit4.n27 GND 0.07fF
C5222 bit4.t2 GND 0.03fF $ **FLOATING
C5223 bit4.n28 GND 0.01fF
C5224 bit4.n29 GND 0.00fF
C5225 bit4.t20 GND 0.03fF $ **FLOATING
C5226 bit4.n30 GND 0.01fF
C5227 bit4.n31 GND 0.00fF
C5228 bit4.n32 GND 0.00fF
C5229 bit4.n33 GND 0.00fF
C5230 bit4.n34 GND 0.07fF
C5231 bit4.t5 GND 0.03fF $ **FLOATING
C5232 bit4.n35 GND 0.01fF
C5233 bit4.n36 GND 0.00fF
C5234 bit4.t17 GND 0.03fF $ **FLOATING
C5235 bit4.n37 GND 0.01fF
C5236 bit4.n38 GND 0.00fF
C5237 bit4.n39 GND 0.00fF
C5238 bit4.n40 GND 0.00fF
C5239 bit4.n41 GND 0.07fF
C5240 bit4.t3 GND 0.03fF $ **FLOATING
C5241 bit4.n42 GND 0.01fF
C5242 bit4.n43 GND 0.00fF
C5243 bit4.t22 GND 0.03fF $ **FLOATING
C5244 bit4.n44 GND 0.01fF
C5245 bit4.n45 GND 0.00fF
C5246 bit4.n46 GND 0.00fF
C5247 bit4.n47 GND 0.00fF
C5248 bit4.n48 GND 0.07fF
C5249 bit4.n49 GND 0.00fF
C5250 bit4.n50 GND 0.00fF
C5251 bit4.t10 GND 0.03fF $ **FLOATING
C5252 bit4.n51 GND 0.01fF
C5253 bit4.n52 GND 0.00fF
C5254 bit4.t29 GND 0.03fF $ **FLOATING
C5255 bit4.n53 GND 0.01fF
C5256 bit4.n54 GND 0.00fF
C5257 bit4.n55 GND 12.02fF
C5258 bit4.n56 GND 24.36fF
C5259 bit4.n57 GND 18.17fF
C5260 bit4.n58 GND 18.17fF
C5261 bit4.n59 GND 18.17fF
C5262 bit4.n60 GND 18.17fF
C5263 bit4.n61 GND 18.17fF
C5264 bit4.n62 GND 29.12fF
C5265 bit4.t24 GND 0.03fF $ **FLOATING
C5266 bit4.n63 GND 0.01fF
C5267 bit4.n64 GND 0.00fF
C5268 bit4.t8 GND 0.03fF $ **FLOATING
C5269 bit4.n65 GND 0.01fF
C5270 bit4.n66 GND 0.00fF
C5271 bit4.n67 GND 0.00fF
C5272 bit4.n68 GND 0.00fF
C5273 bit4.n69 GND 0.07fF
C5274 bit4.t21 GND 0.03fF $ **FLOATING
C5275 bit4.n70 GND 0.01fF
C5276 bit4.n71 GND 0.00fF
C5277 bit4.t9 GND 0.03fF $ **FLOATING
C5278 bit4.n72 GND 0.01fF
C5279 bit4.n73 GND 0.00fF
C5280 bit4.n74 GND 0.00fF
C5281 bit4.n75 GND 0.00fF
C5282 bit4.n76 GND 0.07fF
C5283 bit4.t1 GND 0.03fF $ **FLOATING
C5284 bit4.n77 GND 0.01fF
C5285 bit4.n78 GND 0.00fF
C5286 bit4.t18 GND 0.03fF $ **FLOATING
C5287 bit4.n79 GND 0.01fF
C5288 bit4.n80 GND 0.00fF
C5289 bit4.n81 GND 0.00fF
C5290 bit4.n82 GND 0.00fF
C5291 bit4.n83 GND 0.07fF
C5292 bit4.t33 GND 0.03fF $ **FLOATING
C5293 bit4.n84 GND 0.01fF
C5294 bit4.n85 GND 0.00fF
C5295 bit4.t16 GND 0.03fF $ **FLOATING
C5296 bit4.n86 GND 0.01fF
C5297 bit4.n87 GND 0.00fF
C5298 bit4.n88 GND 0.00fF
C5299 bit4.n89 GND 0.00fF
C5300 bit4.n90 GND 0.07fF
C5301 bit4.t31 GND 0.03fF $ **FLOATING
C5302 bit4.n91 GND 0.01fF
C5303 bit4.n92 GND 0.00fF
C5304 bit4.t14 GND 0.03fF $ **FLOATING
C5305 bit4.n93 GND 0.01fF
C5306 bit4.n94 GND 0.00fF
C5307 bit4.n95 GND 0.00fF
C5308 bit4.n96 GND 0.00fF
C5309 bit4.n97 GND 0.07fF
C5310 bit4.t0 GND 0.03fF $ **FLOATING
C5311 bit4.n98 GND 0.01fF
C5312 bit4.n99 GND 0.00fF
C5313 bit4.t13 GND 0.03fF $ **FLOATING
C5314 bit4.n100 GND 0.01fF
C5315 bit4.n101 GND 0.00fF
C5316 bit4.n102 GND 0.00fF
C5317 bit4.n103 GND 0.00fF
C5318 bit4.n104 GND 0.07fF
C5319 bit4.t32 GND 0.03fF $ **FLOATING
C5320 bit4.n105 GND 0.01fF
C5321 bit4.n106 GND 0.00fF
C5322 bit4.t15 GND 0.03fF $ **FLOATING
C5323 bit4.n107 GND 0.01fF
C5324 bit4.n108 GND 0.00fF
C5325 bit4.n109 GND 0.00fF
C5326 bit4.n110 GND 0.00fF
C5327 bit4.n111 GND 0.07fF
C5328 bit4.t7 GND 0.03fF $ **FLOATING
C5329 bit4.n112 GND 0.01fF
C5330 bit4.n113 GND 0.00fF
C5331 bit4.t27 GND 0.03fF $ **FLOATING
C5332 bit4.n114 GND 0.01fF
C5333 bit4.n115 GND 0.00fF
C5334 bit4.n116 GND 0.00fF
C5335 bit4.n117 GND 0.00fF
C5336 bit4.n118 GND 0.07fF
C5337 bit4.t19 GND 0.01fF $ **FLOATING
C5338 bit4.t30 GND 0.01fF $ **FLOATING
C5339 bit4.n119 GND 0.03fF
C5340 bit4.n120 GND 18.52fF
C5341 bit4.n121 GND 18.17fF
C5342 bit4.n122 GND 18.17fF
C5343 bit4.n123 GND 18.17fF
C5344 bit4.n124 GND 18.17fF
C5345 bit4.n125 GND 18.17fF
C5346 bit4.n126 GND 18.17fF
C5347 bit4.n127 GND 20.56fF
C5348 bit4.n128 GND 33.82fF
.ends
