magic
tech sky130B
magscale 1 2
timestamp 1654107163
<< nwell >>
rect -72 394 218 1236
<< pwell >>
rect -72 -120 216 348
<< psubdiff >>
rect -30 -64 168 -62
rect -30 -100 10 -64
rect 48 -100 108 -64
rect 144 -100 168 -64
rect -30 -102 168 -100
<< nsubdiff >>
rect -36 1192 174 1200
rect -36 1154 -12 1192
rect 36 1154 102 1192
rect 150 1154 174 1192
rect -36 1146 174 1154
<< psubdiffcont >>
rect 10 -100 48 -64
rect 108 -100 144 -64
<< nsubdiffcont >>
rect -12 1154 36 1192
rect 102 1154 150 1192
<< poly >>
rect 58 412 88 430
rect -72 372 88 412
rect 58 352 88 372
<< locali >>
rect -72 1192 216 1220
rect -72 1154 -12 1192
rect 36 1154 102 1192
rect 150 1154 216 1192
rect -72 1118 216 1154
rect 12 1060 46 1118
rect 100 412 134 452
rect 100 372 218 412
rect 100 330 134 372
rect 12 -42 46 22
rect -72 -64 216 -42
rect -72 -100 10 -64
rect 48 -100 108 -64
rect 144 -100 216 -64
rect -72 -120 216 -100
use sky130_fd_pr__nfet_01v8_S96UGK  sky130_fd_pr__nfet_01v8_S96UGK_0
timestamp 1654103908
transform 1 0 73 0 1 176
box -73 -176 73 176
use sky130_fd_pr__pfet_01v8_5EUT2B  sky130_fd_pr__pfet_01v8_5EUT2B_0
timestamp 1654103908
transform 1 0 73 0 1 756
box -109 -362 109 362
<< labels >>
flabel locali -72 1164 -72 1164 0 FreeSans 320 0 0 0 VDD
port 0 nsew
flabel locali -72 -78 -72 -78 0 FreeSans 320 0 0 0 GND
port 1 nsew
flabel poly -72 388 -72 388 0 FreeSans 320 0 0 0 IN
port 2 nsew
flabel locali 218 392 218 392 0 FreeSans 320 0 0 0 OUT
port 3 nsew
<< end >>
