magic
tech sky130B
magscale 1 2
timestamp 1654424809
<< nwell >>
rect -508 94734 -218 95576
rect -508 84854 -218 85696
rect -508 74974 -218 75816
rect -508 65094 -218 65936
rect -508 45334 -218 46176
rect -508 5814 -218 6656
<< pwell >>
rect 4124 94836 5034 96000
rect -506 94220 -218 94688
rect 4124 84956 5034 86120
rect 13324 84956 14234 86120
rect -506 84340 -218 84808
rect 4124 75076 5034 76240
rect 13324 75076 14234 76240
rect 22524 75076 23434 76240
rect 31724 75076 32634 76240
rect -506 74460 -218 74928
rect 4124 65196 5034 66360
rect 13324 65196 14234 66360
rect 22524 65196 23434 66360
rect 31724 65196 32634 66360
rect 40924 65196 41834 66360
rect 50124 65196 51034 66360
rect 59324 65196 60234 66360
rect 68524 65196 69434 66360
rect -506 64580 -218 65048
rect 4124 55316 5034 56480
rect 13324 55316 14234 56480
rect 22524 55316 23434 56480
rect 31724 55316 32634 56480
rect 40924 55316 41834 56480
rect 50124 55316 51034 56480
rect 59324 55316 60234 56480
rect 68524 55316 69434 56480
rect 4124 45436 5034 46600
rect 13324 45436 14234 46600
rect 22524 45436 23434 46600
rect 31724 45436 32634 46600
rect 40924 45436 41834 46600
rect 50124 45436 51034 46600
rect 59324 45436 60234 46600
rect 68524 45436 69434 46600
rect -506 44820 -218 45288
rect 4124 35556 5034 36720
rect 13324 35556 14234 36720
rect 22524 35556 23434 36720
rect 31724 35556 32634 36720
rect 40924 35556 41834 36720
rect 50124 35556 51034 36720
rect 59324 35556 60234 36720
rect 68524 35556 69434 36720
rect 4124 25676 5034 26840
rect 13324 25676 14234 26840
rect 22524 25676 23434 26840
rect 31724 25676 32634 26840
rect 40924 25676 41834 26840
rect 50124 25676 51034 26840
rect 59324 25676 60234 26840
rect 68524 25676 69434 26840
rect 4124 15796 5034 16960
rect 13324 15796 14234 16960
rect 22524 15796 23434 16960
rect 31724 15796 32634 16960
rect 40924 15796 41834 16960
rect 50124 15796 51034 16960
rect 59324 15796 60234 16960
rect 68524 15796 69434 16960
rect 4124 5916 5034 7080
rect 13324 5916 14234 7080
rect 22524 5916 23434 7080
rect 31724 5916 32634 7080
rect 40924 5916 41834 7080
rect 50124 5916 51034 7080
rect 59324 5916 60234 7080
rect 68524 5916 69434 7080
rect -506 5300 -218 5768
<< nmos >>
rect 4522 94962 4552 95292
rect 4608 94962 4638 95292
rect -378 94366 -348 94666
rect 4522 85082 4552 85412
rect 4608 85082 4638 85412
rect 13722 85082 13752 85412
rect 13808 85082 13838 85412
rect -378 84486 -348 84786
rect 4522 75202 4552 75532
rect 4608 75202 4638 75532
rect 13722 75202 13752 75532
rect 13808 75202 13838 75532
rect 22922 75202 22952 75532
rect 23008 75202 23038 75532
rect 32122 75202 32152 75532
rect 32208 75202 32238 75532
rect -378 74606 -348 74906
rect 4522 65322 4552 65652
rect 4608 65322 4638 65652
rect 13722 65322 13752 65652
rect 13808 65322 13838 65652
rect 22922 65322 22952 65652
rect 23008 65322 23038 65652
rect 32122 65322 32152 65652
rect 32208 65322 32238 65652
rect 41322 65322 41352 65652
rect 41408 65322 41438 65652
rect 50522 65322 50552 65652
rect 50608 65322 50638 65652
rect 59722 65322 59752 65652
rect 59808 65322 59838 65652
rect 68922 65322 68952 65652
rect 69008 65322 69038 65652
rect -378 64726 -348 65026
rect 4522 55442 4552 55772
rect 4608 55442 4638 55772
rect 13722 55442 13752 55772
rect 13808 55442 13838 55772
rect 22922 55442 22952 55772
rect 23008 55442 23038 55772
rect 32122 55442 32152 55772
rect 32208 55442 32238 55772
rect 41322 55442 41352 55772
rect 41408 55442 41438 55772
rect 50522 55442 50552 55772
rect 50608 55442 50638 55772
rect 59722 55442 59752 55772
rect 59808 55442 59838 55772
rect 68922 55442 68952 55772
rect 69008 55442 69038 55772
rect 4522 45562 4552 45892
rect 4608 45562 4638 45892
rect 13722 45562 13752 45892
rect 13808 45562 13838 45892
rect 22922 45562 22952 45892
rect 23008 45562 23038 45892
rect 32122 45562 32152 45892
rect 32208 45562 32238 45892
rect 41322 45562 41352 45892
rect 41408 45562 41438 45892
rect 50522 45562 50552 45892
rect 50608 45562 50638 45892
rect 59722 45562 59752 45892
rect 59808 45562 59838 45892
rect 68922 45562 68952 45892
rect 69008 45562 69038 45892
rect -378 44966 -348 45266
rect 4522 35682 4552 36012
rect 4608 35682 4638 36012
rect 13722 35682 13752 36012
rect 13808 35682 13838 36012
rect 22922 35682 22952 36012
rect 23008 35682 23038 36012
rect 32122 35682 32152 36012
rect 32208 35682 32238 36012
rect 41322 35682 41352 36012
rect 41408 35682 41438 36012
rect 50522 35682 50552 36012
rect 50608 35682 50638 36012
rect 59722 35682 59752 36012
rect 59808 35682 59838 36012
rect 68922 35682 68952 36012
rect 69008 35682 69038 36012
rect 4522 25802 4552 26132
rect 4608 25802 4638 26132
rect 13722 25802 13752 26132
rect 13808 25802 13838 26132
rect 22922 25802 22952 26132
rect 23008 25802 23038 26132
rect 32122 25802 32152 26132
rect 32208 25802 32238 26132
rect 41322 25802 41352 26132
rect 41408 25802 41438 26132
rect 50522 25802 50552 26132
rect 50608 25802 50638 26132
rect 59722 25802 59752 26132
rect 59808 25802 59838 26132
rect 68922 25802 68952 26132
rect 69008 25802 69038 26132
rect 4522 15922 4552 16252
rect 4608 15922 4638 16252
rect 13722 15922 13752 16252
rect 13808 15922 13838 16252
rect 22922 15922 22952 16252
rect 23008 15922 23038 16252
rect 32122 15922 32152 16252
rect 32208 15922 32238 16252
rect 41322 15922 41352 16252
rect 41408 15922 41438 16252
rect 50522 15922 50552 16252
rect 50608 15922 50638 16252
rect 59722 15922 59752 16252
rect 59808 15922 59838 16252
rect 68922 15922 68952 16252
rect 69008 15922 69038 16252
rect 4522 6042 4552 6372
rect 4608 6042 4638 6372
rect 13722 6042 13752 6372
rect 13808 6042 13838 6372
rect 22922 6042 22952 6372
rect 23008 6042 23038 6372
rect 32122 6042 32152 6372
rect 32208 6042 32238 6372
rect 41322 6042 41352 6372
rect 41408 6042 41438 6372
rect 50522 6042 50552 6372
rect 50608 6042 50638 6372
rect 59722 6042 59752 6372
rect 59808 6042 59838 6372
rect 68922 6042 68952 6372
rect 69008 6042 69038 6372
rect -378 5446 -348 5746
<< pmos >>
rect -378 94796 -348 95396
rect -378 84916 -348 85516
rect -378 75036 -348 75636
rect -378 65156 -348 65756
rect -378 45396 -348 45996
rect -378 5876 -348 6476
<< ndiff >>
rect 4466 95280 4522 95292
rect 4466 95246 4477 95280
rect 4511 95246 4522 95280
rect 4466 95212 4522 95246
rect 4466 95178 4477 95212
rect 4511 95178 4522 95212
rect 4466 95144 4522 95178
rect 4466 95110 4477 95144
rect 4511 95110 4522 95144
rect 4466 95076 4522 95110
rect 4466 95042 4477 95076
rect 4511 95042 4522 95076
rect 4466 95008 4522 95042
rect 4466 94974 4477 95008
rect 4511 94974 4522 95008
rect 4466 94962 4522 94974
rect 4552 95280 4608 95292
rect 4552 95246 4563 95280
rect 4597 95246 4608 95280
rect 4552 95212 4608 95246
rect 4552 95178 4563 95212
rect 4597 95178 4608 95212
rect 4552 95144 4608 95178
rect 4552 95110 4563 95144
rect 4597 95110 4608 95144
rect 4552 95076 4608 95110
rect 4552 95042 4563 95076
rect 4597 95042 4608 95076
rect 4552 95008 4608 95042
rect 4552 94974 4563 95008
rect 4597 94974 4608 95008
rect 4552 94962 4608 94974
rect 4638 95280 4694 95292
rect 4638 95246 4649 95280
rect 4683 95246 4694 95280
rect 4638 95212 4694 95246
rect 4638 95178 4649 95212
rect 4683 95178 4694 95212
rect 4638 95144 4694 95178
rect 4638 95110 4649 95144
rect 4683 95110 4694 95144
rect 4638 95076 4694 95110
rect 4638 95042 4649 95076
rect 4683 95042 4694 95076
rect 4638 95008 4694 95042
rect 4638 94974 4649 95008
rect 4683 94974 4694 95008
rect 4638 94962 4694 94974
rect -436 94654 -378 94666
rect -436 94378 -424 94654
rect -390 94378 -378 94654
rect -436 94366 -378 94378
rect -348 94654 -290 94666
rect -348 94378 -336 94654
rect -302 94378 -290 94654
rect -348 94366 -290 94378
rect 4466 85400 4522 85412
rect 4466 85366 4477 85400
rect 4511 85366 4522 85400
rect 4466 85332 4522 85366
rect 4466 85298 4477 85332
rect 4511 85298 4522 85332
rect 4466 85264 4522 85298
rect 4466 85230 4477 85264
rect 4511 85230 4522 85264
rect 4466 85196 4522 85230
rect 4466 85162 4477 85196
rect 4511 85162 4522 85196
rect 4466 85128 4522 85162
rect 4466 85094 4477 85128
rect 4511 85094 4522 85128
rect 4466 85082 4522 85094
rect 4552 85400 4608 85412
rect 4552 85366 4563 85400
rect 4597 85366 4608 85400
rect 4552 85332 4608 85366
rect 4552 85298 4563 85332
rect 4597 85298 4608 85332
rect 4552 85264 4608 85298
rect 4552 85230 4563 85264
rect 4597 85230 4608 85264
rect 4552 85196 4608 85230
rect 4552 85162 4563 85196
rect 4597 85162 4608 85196
rect 4552 85128 4608 85162
rect 4552 85094 4563 85128
rect 4597 85094 4608 85128
rect 4552 85082 4608 85094
rect 4638 85400 4694 85412
rect 4638 85366 4649 85400
rect 4683 85366 4694 85400
rect 4638 85332 4694 85366
rect 4638 85298 4649 85332
rect 4683 85298 4694 85332
rect 4638 85264 4694 85298
rect 4638 85230 4649 85264
rect 4683 85230 4694 85264
rect 4638 85196 4694 85230
rect 4638 85162 4649 85196
rect 4683 85162 4694 85196
rect 4638 85128 4694 85162
rect 4638 85094 4649 85128
rect 4683 85094 4694 85128
rect 4638 85082 4694 85094
rect 13666 85400 13722 85412
rect 13666 85366 13677 85400
rect 13711 85366 13722 85400
rect 13666 85332 13722 85366
rect 13666 85298 13677 85332
rect 13711 85298 13722 85332
rect 13666 85264 13722 85298
rect 13666 85230 13677 85264
rect 13711 85230 13722 85264
rect 13666 85196 13722 85230
rect 13666 85162 13677 85196
rect 13711 85162 13722 85196
rect 13666 85128 13722 85162
rect 13666 85094 13677 85128
rect 13711 85094 13722 85128
rect 13666 85082 13722 85094
rect 13752 85400 13808 85412
rect 13752 85366 13763 85400
rect 13797 85366 13808 85400
rect 13752 85332 13808 85366
rect 13752 85298 13763 85332
rect 13797 85298 13808 85332
rect 13752 85264 13808 85298
rect 13752 85230 13763 85264
rect 13797 85230 13808 85264
rect 13752 85196 13808 85230
rect 13752 85162 13763 85196
rect 13797 85162 13808 85196
rect 13752 85128 13808 85162
rect 13752 85094 13763 85128
rect 13797 85094 13808 85128
rect 13752 85082 13808 85094
rect 13838 85400 13894 85412
rect 13838 85366 13849 85400
rect 13883 85366 13894 85400
rect 13838 85332 13894 85366
rect 13838 85298 13849 85332
rect 13883 85298 13894 85332
rect 13838 85264 13894 85298
rect 13838 85230 13849 85264
rect 13883 85230 13894 85264
rect 13838 85196 13894 85230
rect 13838 85162 13849 85196
rect 13883 85162 13894 85196
rect 13838 85128 13894 85162
rect 13838 85094 13849 85128
rect 13883 85094 13894 85128
rect 13838 85082 13894 85094
rect -436 84774 -378 84786
rect -436 84498 -424 84774
rect -390 84498 -378 84774
rect -436 84486 -378 84498
rect -348 84774 -290 84786
rect -348 84498 -336 84774
rect -302 84498 -290 84774
rect -348 84486 -290 84498
rect 4466 75520 4522 75532
rect 4466 75486 4477 75520
rect 4511 75486 4522 75520
rect 4466 75452 4522 75486
rect 4466 75418 4477 75452
rect 4511 75418 4522 75452
rect 4466 75384 4522 75418
rect 4466 75350 4477 75384
rect 4511 75350 4522 75384
rect 4466 75316 4522 75350
rect 4466 75282 4477 75316
rect 4511 75282 4522 75316
rect 4466 75248 4522 75282
rect 4466 75214 4477 75248
rect 4511 75214 4522 75248
rect 4466 75202 4522 75214
rect 4552 75520 4608 75532
rect 4552 75486 4563 75520
rect 4597 75486 4608 75520
rect 4552 75452 4608 75486
rect 4552 75418 4563 75452
rect 4597 75418 4608 75452
rect 4552 75384 4608 75418
rect 4552 75350 4563 75384
rect 4597 75350 4608 75384
rect 4552 75316 4608 75350
rect 4552 75282 4563 75316
rect 4597 75282 4608 75316
rect 4552 75248 4608 75282
rect 4552 75214 4563 75248
rect 4597 75214 4608 75248
rect 4552 75202 4608 75214
rect 4638 75520 4694 75532
rect 4638 75486 4649 75520
rect 4683 75486 4694 75520
rect 4638 75452 4694 75486
rect 4638 75418 4649 75452
rect 4683 75418 4694 75452
rect 4638 75384 4694 75418
rect 4638 75350 4649 75384
rect 4683 75350 4694 75384
rect 4638 75316 4694 75350
rect 4638 75282 4649 75316
rect 4683 75282 4694 75316
rect 4638 75248 4694 75282
rect 4638 75214 4649 75248
rect 4683 75214 4694 75248
rect 4638 75202 4694 75214
rect 13666 75520 13722 75532
rect 13666 75486 13677 75520
rect 13711 75486 13722 75520
rect 13666 75452 13722 75486
rect 13666 75418 13677 75452
rect 13711 75418 13722 75452
rect 13666 75384 13722 75418
rect 13666 75350 13677 75384
rect 13711 75350 13722 75384
rect 13666 75316 13722 75350
rect 13666 75282 13677 75316
rect 13711 75282 13722 75316
rect 13666 75248 13722 75282
rect 13666 75214 13677 75248
rect 13711 75214 13722 75248
rect 13666 75202 13722 75214
rect 13752 75520 13808 75532
rect 13752 75486 13763 75520
rect 13797 75486 13808 75520
rect 13752 75452 13808 75486
rect 13752 75418 13763 75452
rect 13797 75418 13808 75452
rect 13752 75384 13808 75418
rect 13752 75350 13763 75384
rect 13797 75350 13808 75384
rect 13752 75316 13808 75350
rect 13752 75282 13763 75316
rect 13797 75282 13808 75316
rect 13752 75248 13808 75282
rect 13752 75214 13763 75248
rect 13797 75214 13808 75248
rect 13752 75202 13808 75214
rect 13838 75520 13894 75532
rect 13838 75486 13849 75520
rect 13883 75486 13894 75520
rect 13838 75452 13894 75486
rect 13838 75418 13849 75452
rect 13883 75418 13894 75452
rect 13838 75384 13894 75418
rect 13838 75350 13849 75384
rect 13883 75350 13894 75384
rect 13838 75316 13894 75350
rect 13838 75282 13849 75316
rect 13883 75282 13894 75316
rect 13838 75248 13894 75282
rect 13838 75214 13849 75248
rect 13883 75214 13894 75248
rect 13838 75202 13894 75214
rect 22866 75520 22922 75532
rect 22866 75486 22877 75520
rect 22911 75486 22922 75520
rect 22866 75452 22922 75486
rect 22866 75418 22877 75452
rect 22911 75418 22922 75452
rect 22866 75384 22922 75418
rect 22866 75350 22877 75384
rect 22911 75350 22922 75384
rect 22866 75316 22922 75350
rect 22866 75282 22877 75316
rect 22911 75282 22922 75316
rect 22866 75248 22922 75282
rect 22866 75214 22877 75248
rect 22911 75214 22922 75248
rect 22866 75202 22922 75214
rect 22952 75520 23008 75532
rect 22952 75486 22963 75520
rect 22997 75486 23008 75520
rect 22952 75452 23008 75486
rect 22952 75418 22963 75452
rect 22997 75418 23008 75452
rect 22952 75384 23008 75418
rect 22952 75350 22963 75384
rect 22997 75350 23008 75384
rect 22952 75316 23008 75350
rect 22952 75282 22963 75316
rect 22997 75282 23008 75316
rect 22952 75248 23008 75282
rect 22952 75214 22963 75248
rect 22997 75214 23008 75248
rect 22952 75202 23008 75214
rect 23038 75520 23094 75532
rect 23038 75486 23049 75520
rect 23083 75486 23094 75520
rect 23038 75452 23094 75486
rect 23038 75418 23049 75452
rect 23083 75418 23094 75452
rect 23038 75384 23094 75418
rect 23038 75350 23049 75384
rect 23083 75350 23094 75384
rect 23038 75316 23094 75350
rect 23038 75282 23049 75316
rect 23083 75282 23094 75316
rect 23038 75248 23094 75282
rect 23038 75214 23049 75248
rect 23083 75214 23094 75248
rect 23038 75202 23094 75214
rect 32066 75520 32122 75532
rect 32066 75486 32077 75520
rect 32111 75486 32122 75520
rect 32066 75452 32122 75486
rect 32066 75418 32077 75452
rect 32111 75418 32122 75452
rect 32066 75384 32122 75418
rect 32066 75350 32077 75384
rect 32111 75350 32122 75384
rect 32066 75316 32122 75350
rect 32066 75282 32077 75316
rect 32111 75282 32122 75316
rect 32066 75248 32122 75282
rect 32066 75214 32077 75248
rect 32111 75214 32122 75248
rect 32066 75202 32122 75214
rect 32152 75520 32208 75532
rect 32152 75486 32163 75520
rect 32197 75486 32208 75520
rect 32152 75452 32208 75486
rect 32152 75418 32163 75452
rect 32197 75418 32208 75452
rect 32152 75384 32208 75418
rect 32152 75350 32163 75384
rect 32197 75350 32208 75384
rect 32152 75316 32208 75350
rect 32152 75282 32163 75316
rect 32197 75282 32208 75316
rect 32152 75248 32208 75282
rect 32152 75214 32163 75248
rect 32197 75214 32208 75248
rect 32152 75202 32208 75214
rect 32238 75520 32294 75532
rect 32238 75486 32249 75520
rect 32283 75486 32294 75520
rect 32238 75452 32294 75486
rect 32238 75418 32249 75452
rect 32283 75418 32294 75452
rect 32238 75384 32294 75418
rect 32238 75350 32249 75384
rect 32283 75350 32294 75384
rect 32238 75316 32294 75350
rect 32238 75282 32249 75316
rect 32283 75282 32294 75316
rect 32238 75248 32294 75282
rect 32238 75214 32249 75248
rect 32283 75214 32294 75248
rect 32238 75202 32294 75214
rect -436 74894 -378 74906
rect -436 74618 -424 74894
rect -390 74618 -378 74894
rect -436 74606 -378 74618
rect -348 74894 -290 74906
rect -348 74618 -336 74894
rect -302 74618 -290 74894
rect -348 74606 -290 74618
rect 4466 65640 4522 65652
rect 4466 65606 4477 65640
rect 4511 65606 4522 65640
rect 4466 65572 4522 65606
rect 4466 65538 4477 65572
rect 4511 65538 4522 65572
rect 4466 65504 4522 65538
rect 4466 65470 4477 65504
rect 4511 65470 4522 65504
rect 4466 65436 4522 65470
rect 4466 65402 4477 65436
rect 4511 65402 4522 65436
rect 4466 65368 4522 65402
rect 4466 65334 4477 65368
rect 4511 65334 4522 65368
rect 4466 65322 4522 65334
rect 4552 65640 4608 65652
rect 4552 65606 4563 65640
rect 4597 65606 4608 65640
rect 4552 65572 4608 65606
rect 4552 65538 4563 65572
rect 4597 65538 4608 65572
rect 4552 65504 4608 65538
rect 4552 65470 4563 65504
rect 4597 65470 4608 65504
rect 4552 65436 4608 65470
rect 4552 65402 4563 65436
rect 4597 65402 4608 65436
rect 4552 65368 4608 65402
rect 4552 65334 4563 65368
rect 4597 65334 4608 65368
rect 4552 65322 4608 65334
rect 4638 65640 4694 65652
rect 4638 65606 4649 65640
rect 4683 65606 4694 65640
rect 4638 65572 4694 65606
rect 4638 65538 4649 65572
rect 4683 65538 4694 65572
rect 4638 65504 4694 65538
rect 4638 65470 4649 65504
rect 4683 65470 4694 65504
rect 4638 65436 4694 65470
rect 4638 65402 4649 65436
rect 4683 65402 4694 65436
rect 4638 65368 4694 65402
rect 4638 65334 4649 65368
rect 4683 65334 4694 65368
rect 4638 65322 4694 65334
rect 13666 65640 13722 65652
rect 13666 65606 13677 65640
rect 13711 65606 13722 65640
rect 13666 65572 13722 65606
rect 13666 65538 13677 65572
rect 13711 65538 13722 65572
rect 13666 65504 13722 65538
rect 13666 65470 13677 65504
rect 13711 65470 13722 65504
rect 13666 65436 13722 65470
rect 13666 65402 13677 65436
rect 13711 65402 13722 65436
rect 13666 65368 13722 65402
rect 13666 65334 13677 65368
rect 13711 65334 13722 65368
rect 13666 65322 13722 65334
rect 13752 65640 13808 65652
rect 13752 65606 13763 65640
rect 13797 65606 13808 65640
rect 13752 65572 13808 65606
rect 13752 65538 13763 65572
rect 13797 65538 13808 65572
rect 13752 65504 13808 65538
rect 13752 65470 13763 65504
rect 13797 65470 13808 65504
rect 13752 65436 13808 65470
rect 13752 65402 13763 65436
rect 13797 65402 13808 65436
rect 13752 65368 13808 65402
rect 13752 65334 13763 65368
rect 13797 65334 13808 65368
rect 13752 65322 13808 65334
rect 13838 65640 13894 65652
rect 13838 65606 13849 65640
rect 13883 65606 13894 65640
rect 13838 65572 13894 65606
rect 13838 65538 13849 65572
rect 13883 65538 13894 65572
rect 13838 65504 13894 65538
rect 13838 65470 13849 65504
rect 13883 65470 13894 65504
rect 13838 65436 13894 65470
rect 13838 65402 13849 65436
rect 13883 65402 13894 65436
rect 13838 65368 13894 65402
rect 13838 65334 13849 65368
rect 13883 65334 13894 65368
rect 13838 65322 13894 65334
rect 22866 65640 22922 65652
rect 22866 65606 22877 65640
rect 22911 65606 22922 65640
rect 22866 65572 22922 65606
rect 22866 65538 22877 65572
rect 22911 65538 22922 65572
rect 22866 65504 22922 65538
rect 22866 65470 22877 65504
rect 22911 65470 22922 65504
rect 22866 65436 22922 65470
rect 22866 65402 22877 65436
rect 22911 65402 22922 65436
rect 22866 65368 22922 65402
rect 22866 65334 22877 65368
rect 22911 65334 22922 65368
rect 22866 65322 22922 65334
rect 22952 65640 23008 65652
rect 22952 65606 22963 65640
rect 22997 65606 23008 65640
rect 22952 65572 23008 65606
rect 22952 65538 22963 65572
rect 22997 65538 23008 65572
rect 22952 65504 23008 65538
rect 22952 65470 22963 65504
rect 22997 65470 23008 65504
rect 22952 65436 23008 65470
rect 22952 65402 22963 65436
rect 22997 65402 23008 65436
rect 22952 65368 23008 65402
rect 22952 65334 22963 65368
rect 22997 65334 23008 65368
rect 22952 65322 23008 65334
rect 23038 65640 23094 65652
rect 23038 65606 23049 65640
rect 23083 65606 23094 65640
rect 23038 65572 23094 65606
rect 23038 65538 23049 65572
rect 23083 65538 23094 65572
rect 23038 65504 23094 65538
rect 23038 65470 23049 65504
rect 23083 65470 23094 65504
rect 23038 65436 23094 65470
rect 23038 65402 23049 65436
rect 23083 65402 23094 65436
rect 23038 65368 23094 65402
rect 23038 65334 23049 65368
rect 23083 65334 23094 65368
rect 23038 65322 23094 65334
rect 32066 65640 32122 65652
rect 32066 65606 32077 65640
rect 32111 65606 32122 65640
rect 32066 65572 32122 65606
rect 32066 65538 32077 65572
rect 32111 65538 32122 65572
rect 32066 65504 32122 65538
rect 32066 65470 32077 65504
rect 32111 65470 32122 65504
rect 32066 65436 32122 65470
rect 32066 65402 32077 65436
rect 32111 65402 32122 65436
rect 32066 65368 32122 65402
rect 32066 65334 32077 65368
rect 32111 65334 32122 65368
rect 32066 65322 32122 65334
rect 32152 65640 32208 65652
rect 32152 65606 32163 65640
rect 32197 65606 32208 65640
rect 32152 65572 32208 65606
rect 32152 65538 32163 65572
rect 32197 65538 32208 65572
rect 32152 65504 32208 65538
rect 32152 65470 32163 65504
rect 32197 65470 32208 65504
rect 32152 65436 32208 65470
rect 32152 65402 32163 65436
rect 32197 65402 32208 65436
rect 32152 65368 32208 65402
rect 32152 65334 32163 65368
rect 32197 65334 32208 65368
rect 32152 65322 32208 65334
rect 32238 65640 32294 65652
rect 32238 65606 32249 65640
rect 32283 65606 32294 65640
rect 32238 65572 32294 65606
rect 32238 65538 32249 65572
rect 32283 65538 32294 65572
rect 32238 65504 32294 65538
rect 32238 65470 32249 65504
rect 32283 65470 32294 65504
rect 32238 65436 32294 65470
rect 32238 65402 32249 65436
rect 32283 65402 32294 65436
rect 32238 65368 32294 65402
rect 32238 65334 32249 65368
rect 32283 65334 32294 65368
rect 32238 65322 32294 65334
rect 41266 65640 41322 65652
rect 41266 65606 41277 65640
rect 41311 65606 41322 65640
rect 41266 65572 41322 65606
rect 41266 65538 41277 65572
rect 41311 65538 41322 65572
rect 41266 65504 41322 65538
rect 41266 65470 41277 65504
rect 41311 65470 41322 65504
rect 41266 65436 41322 65470
rect 41266 65402 41277 65436
rect 41311 65402 41322 65436
rect 41266 65368 41322 65402
rect 41266 65334 41277 65368
rect 41311 65334 41322 65368
rect 41266 65322 41322 65334
rect 41352 65640 41408 65652
rect 41352 65606 41363 65640
rect 41397 65606 41408 65640
rect 41352 65572 41408 65606
rect 41352 65538 41363 65572
rect 41397 65538 41408 65572
rect 41352 65504 41408 65538
rect 41352 65470 41363 65504
rect 41397 65470 41408 65504
rect 41352 65436 41408 65470
rect 41352 65402 41363 65436
rect 41397 65402 41408 65436
rect 41352 65368 41408 65402
rect 41352 65334 41363 65368
rect 41397 65334 41408 65368
rect 41352 65322 41408 65334
rect 41438 65640 41494 65652
rect 41438 65606 41449 65640
rect 41483 65606 41494 65640
rect 41438 65572 41494 65606
rect 41438 65538 41449 65572
rect 41483 65538 41494 65572
rect 41438 65504 41494 65538
rect 41438 65470 41449 65504
rect 41483 65470 41494 65504
rect 41438 65436 41494 65470
rect 41438 65402 41449 65436
rect 41483 65402 41494 65436
rect 41438 65368 41494 65402
rect 41438 65334 41449 65368
rect 41483 65334 41494 65368
rect 41438 65322 41494 65334
rect 50466 65640 50522 65652
rect 50466 65606 50477 65640
rect 50511 65606 50522 65640
rect 50466 65572 50522 65606
rect 50466 65538 50477 65572
rect 50511 65538 50522 65572
rect 50466 65504 50522 65538
rect 50466 65470 50477 65504
rect 50511 65470 50522 65504
rect 50466 65436 50522 65470
rect 50466 65402 50477 65436
rect 50511 65402 50522 65436
rect 50466 65368 50522 65402
rect 50466 65334 50477 65368
rect 50511 65334 50522 65368
rect 50466 65322 50522 65334
rect 50552 65640 50608 65652
rect 50552 65606 50563 65640
rect 50597 65606 50608 65640
rect 50552 65572 50608 65606
rect 50552 65538 50563 65572
rect 50597 65538 50608 65572
rect 50552 65504 50608 65538
rect 50552 65470 50563 65504
rect 50597 65470 50608 65504
rect 50552 65436 50608 65470
rect 50552 65402 50563 65436
rect 50597 65402 50608 65436
rect 50552 65368 50608 65402
rect 50552 65334 50563 65368
rect 50597 65334 50608 65368
rect 50552 65322 50608 65334
rect 50638 65640 50694 65652
rect 50638 65606 50649 65640
rect 50683 65606 50694 65640
rect 50638 65572 50694 65606
rect 50638 65538 50649 65572
rect 50683 65538 50694 65572
rect 50638 65504 50694 65538
rect 50638 65470 50649 65504
rect 50683 65470 50694 65504
rect 50638 65436 50694 65470
rect 50638 65402 50649 65436
rect 50683 65402 50694 65436
rect 50638 65368 50694 65402
rect 50638 65334 50649 65368
rect 50683 65334 50694 65368
rect 50638 65322 50694 65334
rect 59666 65640 59722 65652
rect 59666 65606 59677 65640
rect 59711 65606 59722 65640
rect 59666 65572 59722 65606
rect 59666 65538 59677 65572
rect 59711 65538 59722 65572
rect 59666 65504 59722 65538
rect 59666 65470 59677 65504
rect 59711 65470 59722 65504
rect 59666 65436 59722 65470
rect 59666 65402 59677 65436
rect 59711 65402 59722 65436
rect 59666 65368 59722 65402
rect 59666 65334 59677 65368
rect 59711 65334 59722 65368
rect 59666 65322 59722 65334
rect 59752 65640 59808 65652
rect 59752 65606 59763 65640
rect 59797 65606 59808 65640
rect 59752 65572 59808 65606
rect 59752 65538 59763 65572
rect 59797 65538 59808 65572
rect 59752 65504 59808 65538
rect 59752 65470 59763 65504
rect 59797 65470 59808 65504
rect 59752 65436 59808 65470
rect 59752 65402 59763 65436
rect 59797 65402 59808 65436
rect 59752 65368 59808 65402
rect 59752 65334 59763 65368
rect 59797 65334 59808 65368
rect 59752 65322 59808 65334
rect 59838 65640 59894 65652
rect 59838 65606 59849 65640
rect 59883 65606 59894 65640
rect 59838 65572 59894 65606
rect 59838 65538 59849 65572
rect 59883 65538 59894 65572
rect 59838 65504 59894 65538
rect 59838 65470 59849 65504
rect 59883 65470 59894 65504
rect 59838 65436 59894 65470
rect 59838 65402 59849 65436
rect 59883 65402 59894 65436
rect 59838 65368 59894 65402
rect 59838 65334 59849 65368
rect 59883 65334 59894 65368
rect 59838 65322 59894 65334
rect 68866 65640 68922 65652
rect 68866 65606 68877 65640
rect 68911 65606 68922 65640
rect 68866 65572 68922 65606
rect 68866 65538 68877 65572
rect 68911 65538 68922 65572
rect 68866 65504 68922 65538
rect 68866 65470 68877 65504
rect 68911 65470 68922 65504
rect 68866 65436 68922 65470
rect 68866 65402 68877 65436
rect 68911 65402 68922 65436
rect 68866 65368 68922 65402
rect 68866 65334 68877 65368
rect 68911 65334 68922 65368
rect 68866 65322 68922 65334
rect 68952 65640 69008 65652
rect 68952 65606 68963 65640
rect 68997 65606 69008 65640
rect 68952 65572 69008 65606
rect 68952 65538 68963 65572
rect 68997 65538 69008 65572
rect 68952 65504 69008 65538
rect 68952 65470 68963 65504
rect 68997 65470 69008 65504
rect 68952 65436 69008 65470
rect 68952 65402 68963 65436
rect 68997 65402 69008 65436
rect 68952 65368 69008 65402
rect 68952 65334 68963 65368
rect 68997 65334 69008 65368
rect 68952 65322 69008 65334
rect 69038 65640 69094 65652
rect 69038 65606 69049 65640
rect 69083 65606 69094 65640
rect 69038 65572 69094 65606
rect 69038 65538 69049 65572
rect 69083 65538 69094 65572
rect 69038 65504 69094 65538
rect 69038 65470 69049 65504
rect 69083 65470 69094 65504
rect 69038 65436 69094 65470
rect 69038 65402 69049 65436
rect 69083 65402 69094 65436
rect 69038 65368 69094 65402
rect 69038 65334 69049 65368
rect 69083 65334 69094 65368
rect 69038 65322 69094 65334
rect -436 65014 -378 65026
rect -436 64738 -424 65014
rect -390 64738 -378 65014
rect -436 64726 -378 64738
rect -348 65014 -290 65026
rect -348 64738 -336 65014
rect -302 64738 -290 65014
rect -348 64726 -290 64738
rect 4466 55760 4522 55772
rect 4466 55726 4477 55760
rect 4511 55726 4522 55760
rect 4466 55692 4522 55726
rect 4466 55658 4477 55692
rect 4511 55658 4522 55692
rect 4466 55624 4522 55658
rect 4466 55590 4477 55624
rect 4511 55590 4522 55624
rect 4466 55556 4522 55590
rect 4466 55522 4477 55556
rect 4511 55522 4522 55556
rect 4466 55488 4522 55522
rect 4466 55454 4477 55488
rect 4511 55454 4522 55488
rect 4466 55442 4522 55454
rect 4552 55760 4608 55772
rect 4552 55726 4563 55760
rect 4597 55726 4608 55760
rect 4552 55692 4608 55726
rect 4552 55658 4563 55692
rect 4597 55658 4608 55692
rect 4552 55624 4608 55658
rect 4552 55590 4563 55624
rect 4597 55590 4608 55624
rect 4552 55556 4608 55590
rect 4552 55522 4563 55556
rect 4597 55522 4608 55556
rect 4552 55488 4608 55522
rect 4552 55454 4563 55488
rect 4597 55454 4608 55488
rect 4552 55442 4608 55454
rect 4638 55760 4694 55772
rect 4638 55726 4649 55760
rect 4683 55726 4694 55760
rect 4638 55692 4694 55726
rect 4638 55658 4649 55692
rect 4683 55658 4694 55692
rect 4638 55624 4694 55658
rect 4638 55590 4649 55624
rect 4683 55590 4694 55624
rect 4638 55556 4694 55590
rect 4638 55522 4649 55556
rect 4683 55522 4694 55556
rect 4638 55488 4694 55522
rect 4638 55454 4649 55488
rect 4683 55454 4694 55488
rect 4638 55442 4694 55454
rect 13666 55760 13722 55772
rect 13666 55726 13677 55760
rect 13711 55726 13722 55760
rect 13666 55692 13722 55726
rect 13666 55658 13677 55692
rect 13711 55658 13722 55692
rect 13666 55624 13722 55658
rect 13666 55590 13677 55624
rect 13711 55590 13722 55624
rect 13666 55556 13722 55590
rect 13666 55522 13677 55556
rect 13711 55522 13722 55556
rect 13666 55488 13722 55522
rect 13666 55454 13677 55488
rect 13711 55454 13722 55488
rect 13666 55442 13722 55454
rect 13752 55760 13808 55772
rect 13752 55726 13763 55760
rect 13797 55726 13808 55760
rect 13752 55692 13808 55726
rect 13752 55658 13763 55692
rect 13797 55658 13808 55692
rect 13752 55624 13808 55658
rect 13752 55590 13763 55624
rect 13797 55590 13808 55624
rect 13752 55556 13808 55590
rect 13752 55522 13763 55556
rect 13797 55522 13808 55556
rect 13752 55488 13808 55522
rect 13752 55454 13763 55488
rect 13797 55454 13808 55488
rect 13752 55442 13808 55454
rect 13838 55760 13894 55772
rect 13838 55726 13849 55760
rect 13883 55726 13894 55760
rect 13838 55692 13894 55726
rect 13838 55658 13849 55692
rect 13883 55658 13894 55692
rect 13838 55624 13894 55658
rect 13838 55590 13849 55624
rect 13883 55590 13894 55624
rect 13838 55556 13894 55590
rect 13838 55522 13849 55556
rect 13883 55522 13894 55556
rect 13838 55488 13894 55522
rect 13838 55454 13849 55488
rect 13883 55454 13894 55488
rect 13838 55442 13894 55454
rect 22866 55760 22922 55772
rect 22866 55726 22877 55760
rect 22911 55726 22922 55760
rect 22866 55692 22922 55726
rect 22866 55658 22877 55692
rect 22911 55658 22922 55692
rect 22866 55624 22922 55658
rect 22866 55590 22877 55624
rect 22911 55590 22922 55624
rect 22866 55556 22922 55590
rect 22866 55522 22877 55556
rect 22911 55522 22922 55556
rect 22866 55488 22922 55522
rect 22866 55454 22877 55488
rect 22911 55454 22922 55488
rect 22866 55442 22922 55454
rect 22952 55760 23008 55772
rect 22952 55726 22963 55760
rect 22997 55726 23008 55760
rect 22952 55692 23008 55726
rect 22952 55658 22963 55692
rect 22997 55658 23008 55692
rect 22952 55624 23008 55658
rect 22952 55590 22963 55624
rect 22997 55590 23008 55624
rect 22952 55556 23008 55590
rect 22952 55522 22963 55556
rect 22997 55522 23008 55556
rect 22952 55488 23008 55522
rect 22952 55454 22963 55488
rect 22997 55454 23008 55488
rect 22952 55442 23008 55454
rect 23038 55760 23094 55772
rect 23038 55726 23049 55760
rect 23083 55726 23094 55760
rect 23038 55692 23094 55726
rect 23038 55658 23049 55692
rect 23083 55658 23094 55692
rect 23038 55624 23094 55658
rect 23038 55590 23049 55624
rect 23083 55590 23094 55624
rect 23038 55556 23094 55590
rect 23038 55522 23049 55556
rect 23083 55522 23094 55556
rect 23038 55488 23094 55522
rect 23038 55454 23049 55488
rect 23083 55454 23094 55488
rect 23038 55442 23094 55454
rect 32066 55760 32122 55772
rect 32066 55726 32077 55760
rect 32111 55726 32122 55760
rect 32066 55692 32122 55726
rect 32066 55658 32077 55692
rect 32111 55658 32122 55692
rect 32066 55624 32122 55658
rect 32066 55590 32077 55624
rect 32111 55590 32122 55624
rect 32066 55556 32122 55590
rect 32066 55522 32077 55556
rect 32111 55522 32122 55556
rect 32066 55488 32122 55522
rect 32066 55454 32077 55488
rect 32111 55454 32122 55488
rect 32066 55442 32122 55454
rect 32152 55760 32208 55772
rect 32152 55726 32163 55760
rect 32197 55726 32208 55760
rect 32152 55692 32208 55726
rect 32152 55658 32163 55692
rect 32197 55658 32208 55692
rect 32152 55624 32208 55658
rect 32152 55590 32163 55624
rect 32197 55590 32208 55624
rect 32152 55556 32208 55590
rect 32152 55522 32163 55556
rect 32197 55522 32208 55556
rect 32152 55488 32208 55522
rect 32152 55454 32163 55488
rect 32197 55454 32208 55488
rect 32152 55442 32208 55454
rect 32238 55760 32294 55772
rect 32238 55726 32249 55760
rect 32283 55726 32294 55760
rect 32238 55692 32294 55726
rect 32238 55658 32249 55692
rect 32283 55658 32294 55692
rect 32238 55624 32294 55658
rect 32238 55590 32249 55624
rect 32283 55590 32294 55624
rect 32238 55556 32294 55590
rect 32238 55522 32249 55556
rect 32283 55522 32294 55556
rect 32238 55488 32294 55522
rect 32238 55454 32249 55488
rect 32283 55454 32294 55488
rect 32238 55442 32294 55454
rect 41266 55760 41322 55772
rect 41266 55726 41277 55760
rect 41311 55726 41322 55760
rect 41266 55692 41322 55726
rect 41266 55658 41277 55692
rect 41311 55658 41322 55692
rect 41266 55624 41322 55658
rect 41266 55590 41277 55624
rect 41311 55590 41322 55624
rect 41266 55556 41322 55590
rect 41266 55522 41277 55556
rect 41311 55522 41322 55556
rect 41266 55488 41322 55522
rect 41266 55454 41277 55488
rect 41311 55454 41322 55488
rect 41266 55442 41322 55454
rect 41352 55760 41408 55772
rect 41352 55726 41363 55760
rect 41397 55726 41408 55760
rect 41352 55692 41408 55726
rect 41352 55658 41363 55692
rect 41397 55658 41408 55692
rect 41352 55624 41408 55658
rect 41352 55590 41363 55624
rect 41397 55590 41408 55624
rect 41352 55556 41408 55590
rect 41352 55522 41363 55556
rect 41397 55522 41408 55556
rect 41352 55488 41408 55522
rect 41352 55454 41363 55488
rect 41397 55454 41408 55488
rect 41352 55442 41408 55454
rect 41438 55760 41494 55772
rect 41438 55726 41449 55760
rect 41483 55726 41494 55760
rect 41438 55692 41494 55726
rect 41438 55658 41449 55692
rect 41483 55658 41494 55692
rect 41438 55624 41494 55658
rect 41438 55590 41449 55624
rect 41483 55590 41494 55624
rect 41438 55556 41494 55590
rect 41438 55522 41449 55556
rect 41483 55522 41494 55556
rect 41438 55488 41494 55522
rect 41438 55454 41449 55488
rect 41483 55454 41494 55488
rect 41438 55442 41494 55454
rect 50466 55760 50522 55772
rect 50466 55726 50477 55760
rect 50511 55726 50522 55760
rect 50466 55692 50522 55726
rect 50466 55658 50477 55692
rect 50511 55658 50522 55692
rect 50466 55624 50522 55658
rect 50466 55590 50477 55624
rect 50511 55590 50522 55624
rect 50466 55556 50522 55590
rect 50466 55522 50477 55556
rect 50511 55522 50522 55556
rect 50466 55488 50522 55522
rect 50466 55454 50477 55488
rect 50511 55454 50522 55488
rect 50466 55442 50522 55454
rect 50552 55760 50608 55772
rect 50552 55726 50563 55760
rect 50597 55726 50608 55760
rect 50552 55692 50608 55726
rect 50552 55658 50563 55692
rect 50597 55658 50608 55692
rect 50552 55624 50608 55658
rect 50552 55590 50563 55624
rect 50597 55590 50608 55624
rect 50552 55556 50608 55590
rect 50552 55522 50563 55556
rect 50597 55522 50608 55556
rect 50552 55488 50608 55522
rect 50552 55454 50563 55488
rect 50597 55454 50608 55488
rect 50552 55442 50608 55454
rect 50638 55760 50694 55772
rect 50638 55726 50649 55760
rect 50683 55726 50694 55760
rect 50638 55692 50694 55726
rect 50638 55658 50649 55692
rect 50683 55658 50694 55692
rect 50638 55624 50694 55658
rect 50638 55590 50649 55624
rect 50683 55590 50694 55624
rect 50638 55556 50694 55590
rect 50638 55522 50649 55556
rect 50683 55522 50694 55556
rect 50638 55488 50694 55522
rect 50638 55454 50649 55488
rect 50683 55454 50694 55488
rect 50638 55442 50694 55454
rect 59666 55760 59722 55772
rect 59666 55726 59677 55760
rect 59711 55726 59722 55760
rect 59666 55692 59722 55726
rect 59666 55658 59677 55692
rect 59711 55658 59722 55692
rect 59666 55624 59722 55658
rect 59666 55590 59677 55624
rect 59711 55590 59722 55624
rect 59666 55556 59722 55590
rect 59666 55522 59677 55556
rect 59711 55522 59722 55556
rect 59666 55488 59722 55522
rect 59666 55454 59677 55488
rect 59711 55454 59722 55488
rect 59666 55442 59722 55454
rect 59752 55760 59808 55772
rect 59752 55726 59763 55760
rect 59797 55726 59808 55760
rect 59752 55692 59808 55726
rect 59752 55658 59763 55692
rect 59797 55658 59808 55692
rect 59752 55624 59808 55658
rect 59752 55590 59763 55624
rect 59797 55590 59808 55624
rect 59752 55556 59808 55590
rect 59752 55522 59763 55556
rect 59797 55522 59808 55556
rect 59752 55488 59808 55522
rect 59752 55454 59763 55488
rect 59797 55454 59808 55488
rect 59752 55442 59808 55454
rect 59838 55760 59894 55772
rect 59838 55726 59849 55760
rect 59883 55726 59894 55760
rect 59838 55692 59894 55726
rect 59838 55658 59849 55692
rect 59883 55658 59894 55692
rect 59838 55624 59894 55658
rect 59838 55590 59849 55624
rect 59883 55590 59894 55624
rect 59838 55556 59894 55590
rect 59838 55522 59849 55556
rect 59883 55522 59894 55556
rect 59838 55488 59894 55522
rect 59838 55454 59849 55488
rect 59883 55454 59894 55488
rect 59838 55442 59894 55454
rect 68866 55760 68922 55772
rect 68866 55726 68877 55760
rect 68911 55726 68922 55760
rect 68866 55692 68922 55726
rect 68866 55658 68877 55692
rect 68911 55658 68922 55692
rect 68866 55624 68922 55658
rect 68866 55590 68877 55624
rect 68911 55590 68922 55624
rect 68866 55556 68922 55590
rect 68866 55522 68877 55556
rect 68911 55522 68922 55556
rect 68866 55488 68922 55522
rect 68866 55454 68877 55488
rect 68911 55454 68922 55488
rect 68866 55442 68922 55454
rect 68952 55760 69008 55772
rect 68952 55726 68963 55760
rect 68997 55726 69008 55760
rect 68952 55692 69008 55726
rect 68952 55658 68963 55692
rect 68997 55658 69008 55692
rect 68952 55624 69008 55658
rect 68952 55590 68963 55624
rect 68997 55590 69008 55624
rect 68952 55556 69008 55590
rect 68952 55522 68963 55556
rect 68997 55522 69008 55556
rect 68952 55488 69008 55522
rect 68952 55454 68963 55488
rect 68997 55454 69008 55488
rect 68952 55442 69008 55454
rect 69038 55760 69094 55772
rect 69038 55726 69049 55760
rect 69083 55726 69094 55760
rect 69038 55692 69094 55726
rect 69038 55658 69049 55692
rect 69083 55658 69094 55692
rect 69038 55624 69094 55658
rect 69038 55590 69049 55624
rect 69083 55590 69094 55624
rect 69038 55556 69094 55590
rect 69038 55522 69049 55556
rect 69083 55522 69094 55556
rect 69038 55488 69094 55522
rect 69038 55454 69049 55488
rect 69083 55454 69094 55488
rect 69038 55442 69094 55454
rect 4466 45880 4522 45892
rect 4466 45846 4477 45880
rect 4511 45846 4522 45880
rect 4466 45812 4522 45846
rect 4466 45778 4477 45812
rect 4511 45778 4522 45812
rect 4466 45744 4522 45778
rect 4466 45710 4477 45744
rect 4511 45710 4522 45744
rect 4466 45676 4522 45710
rect 4466 45642 4477 45676
rect 4511 45642 4522 45676
rect 4466 45608 4522 45642
rect 4466 45574 4477 45608
rect 4511 45574 4522 45608
rect 4466 45562 4522 45574
rect 4552 45880 4608 45892
rect 4552 45846 4563 45880
rect 4597 45846 4608 45880
rect 4552 45812 4608 45846
rect 4552 45778 4563 45812
rect 4597 45778 4608 45812
rect 4552 45744 4608 45778
rect 4552 45710 4563 45744
rect 4597 45710 4608 45744
rect 4552 45676 4608 45710
rect 4552 45642 4563 45676
rect 4597 45642 4608 45676
rect 4552 45608 4608 45642
rect 4552 45574 4563 45608
rect 4597 45574 4608 45608
rect 4552 45562 4608 45574
rect 4638 45880 4694 45892
rect 4638 45846 4649 45880
rect 4683 45846 4694 45880
rect 4638 45812 4694 45846
rect 4638 45778 4649 45812
rect 4683 45778 4694 45812
rect 4638 45744 4694 45778
rect 4638 45710 4649 45744
rect 4683 45710 4694 45744
rect 4638 45676 4694 45710
rect 4638 45642 4649 45676
rect 4683 45642 4694 45676
rect 4638 45608 4694 45642
rect 4638 45574 4649 45608
rect 4683 45574 4694 45608
rect 4638 45562 4694 45574
rect 13666 45880 13722 45892
rect 13666 45846 13677 45880
rect 13711 45846 13722 45880
rect 13666 45812 13722 45846
rect 13666 45778 13677 45812
rect 13711 45778 13722 45812
rect 13666 45744 13722 45778
rect 13666 45710 13677 45744
rect 13711 45710 13722 45744
rect 13666 45676 13722 45710
rect 13666 45642 13677 45676
rect 13711 45642 13722 45676
rect 13666 45608 13722 45642
rect 13666 45574 13677 45608
rect 13711 45574 13722 45608
rect 13666 45562 13722 45574
rect 13752 45880 13808 45892
rect 13752 45846 13763 45880
rect 13797 45846 13808 45880
rect 13752 45812 13808 45846
rect 13752 45778 13763 45812
rect 13797 45778 13808 45812
rect 13752 45744 13808 45778
rect 13752 45710 13763 45744
rect 13797 45710 13808 45744
rect 13752 45676 13808 45710
rect 13752 45642 13763 45676
rect 13797 45642 13808 45676
rect 13752 45608 13808 45642
rect 13752 45574 13763 45608
rect 13797 45574 13808 45608
rect 13752 45562 13808 45574
rect 13838 45880 13894 45892
rect 13838 45846 13849 45880
rect 13883 45846 13894 45880
rect 13838 45812 13894 45846
rect 13838 45778 13849 45812
rect 13883 45778 13894 45812
rect 13838 45744 13894 45778
rect 13838 45710 13849 45744
rect 13883 45710 13894 45744
rect 13838 45676 13894 45710
rect 13838 45642 13849 45676
rect 13883 45642 13894 45676
rect 13838 45608 13894 45642
rect 13838 45574 13849 45608
rect 13883 45574 13894 45608
rect 13838 45562 13894 45574
rect 22866 45880 22922 45892
rect 22866 45846 22877 45880
rect 22911 45846 22922 45880
rect 22866 45812 22922 45846
rect 22866 45778 22877 45812
rect 22911 45778 22922 45812
rect 22866 45744 22922 45778
rect 22866 45710 22877 45744
rect 22911 45710 22922 45744
rect 22866 45676 22922 45710
rect 22866 45642 22877 45676
rect 22911 45642 22922 45676
rect 22866 45608 22922 45642
rect 22866 45574 22877 45608
rect 22911 45574 22922 45608
rect 22866 45562 22922 45574
rect 22952 45880 23008 45892
rect 22952 45846 22963 45880
rect 22997 45846 23008 45880
rect 22952 45812 23008 45846
rect 22952 45778 22963 45812
rect 22997 45778 23008 45812
rect 22952 45744 23008 45778
rect 22952 45710 22963 45744
rect 22997 45710 23008 45744
rect 22952 45676 23008 45710
rect 22952 45642 22963 45676
rect 22997 45642 23008 45676
rect 22952 45608 23008 45642
rect 22952 45574 22963 45608
rect 22997 45574 23008 45608
rect 22952 45562 23008 45574
rect 23038 45880 23094 45892
rect 23038 45846 23049 45880
rect 23083 45846 23094 45880
rect 23038 45812 23094 45846
rect 23038 45778 23049 45812
rect 23083 45778 23094 45812
rect 23038 45744 23094 45778
rect 23038 45710 23049 45744
rect 23083 45710 23094 45744
rect 23038 45676 23094 45710
rect 23038 45642 23049 45676
rect 23083 45642 23094 45676
rect 23038 45608 23094 45642
rect 23038 45574 23049 45608
rect 23083 45574 23094 45608
rect 23038 45562 23094 45574
rect 32066 45880 32122 45892
rect 32066 45846 32077 45880
rect 32111 45846 32122 45880
rect 32066 45812 32122 45846
rect 32066 45778 32077 45812
rect 32111 45778 32122 45812
rect 32066 45744 32122 45778
rect 32066 45710 32077 45744
rect 32111 45710 32122 45744
rect 32066 45676 32122 45710
rect 32066 45642 32077 45676
rect 32111 45642 32122 45676
rect 32066 45608 32122 45642
rect 32066 45574 32077 45608
rect 32111 45574 32122 45608
rect 32066 45562 32122 45574
rect 32152 45880 32208 45892
rect 32152 45846 32163 45880
rect 32197 45846 32208 45880
rect 32152 45812 32208 45846
rect 32152 45778 32163 45812
rect 32197 45778 32208 45812
rect 32152 45744 32208 45778
rect 32152 45710 32163 45744
rect 32197 45710 32208 45744
rect 32152 45676 32208 45710
rect 32152 45642 32163 45676
rect 32197 45642 32208 45676
rect 32152 45608 32208 45642
rect 32152 45574 32163 45608
rect 32197 45574 32208 45608
rect 32152 45562 32208 45574
rect 32238 45880 32294 45892
rect 32238 45846 32249 45880
rect 32283 45846 32294 45880
rect 32238 45812 32294 45846
rect 32238 45778 32249 45812
rect 32283 45778 32294 45812
rect 32238 45744 32294 45778
rect 32238 45710 32249 45744
rect 32283 45710 32294 45744
rect 32238 45676 32294 45710
rect 32238 45642 32249 45676
rect 32283 45642 32294 45676
rect 32238 45608 32294 45642
rect 32238 45574 32249 45608
rect 32283 45574 32294 45608
rect 32238 45562 32294 45574
rect 41266 45880 41322 45892
rect 41266 45846 41277 45880
rect 41311 45846 41322 45880
rect 41266 45812 41322 45846
rect 41266 45778 41277 45812
rect 41311 45778 41322 45812
rect 41266 45744 41322 45778
rect 41266 45710 41277 45744
rect 41311 45710 41322 45744
rect 41266 45676 41322 45710
rect 41266 45642 41277 45676
rect 41311 45642 41322 45676
rect 41266 45608 41322 45642
rect 41266 45574 41277 45608
rect 41311 45574 41322 45608
rect 41266 45562 41322 45574
rect 41352 45880 41408 45892
rect 41352 45846 41363 45880
rect 41397 45846 41408 45880
rect 41352 45812 41408 45846
rect 41352 45778 41363 45812
rect 41397 45778 41408 45812
rect 41352 45744 41408 45778
rect 41352 45710 41363 45744
rect 41397 45710 41408 45744
rect 41352 45676 41408 45710
rect 41352 45642 41363 45676
rect 41397 45642 41408 45676
rect 41352 45608 41408 45642
rect 41352 45574 41363 45608
rect 41397 45574 41408 45608
rect 41352 45562 41408 45574
rect 41438 45880 41494 45892
rect 41438 45846 41449 45880
rect 41483 45846 41494 45880
rect 41438 45812 41494 45846
rect 41438 45778 41449 45812
rect 41483 45778 41494 45812
rect 41438 45744 41494 45778
rect 41438 45710 41449 45744
rect 41483 45710 41494 45744
rect 41438 45676 41494 45710
rect 41438 45642 41449 45676
rect 41483 45642 41494 45676
rect 41438 45608 41494 45642
rect 41438 45574 41449 45608
rect 41483 45574 41494 45608
rect 41438 45562 41494 45574
rect 50466 45880 50522 45892
rect 50466 45846 50477 45880
rect 50511 45846 50522 45880
rect 50466 45812 50522 45846
rect 50466 45778 50477 45812
rect 50511 45778 50522 45812
rect 50466 45744 50522 45778
rect 50466 45710 50477 45744
rect 50511 45710 50522 45744
rect 50466 45676 50522 45710
rect 50466 45642 50477 45676
rect 50511 45642 50522 45676
rect 50466 45608 50522 45642
rect 50466 45574 50477 45608
rect 50511 45574 50522 45608
rect 50466 45562 50522 45574
rect 50552 45880 50608 45892
rect 50552 45846 50563 45880
rect 50597 45846 50608 45880
rect 50552 45812 50608 45846
rect 50552 45778 50563 45812
rect 50597 45778 50608 45812
rect 50552 45744 50608 45778
rect 50552 45710 50563 45744
rect 50597 45710 50608 45744
rect 50552 45676 50608 45710
rect 50552 45642 50563 45676
rect 50597 45642 50608 45676
rect 50552 45608 50608 45642
rect 50552 45574 50563 45608
rect 50597 45574 50608 45608
rect 50552 45562 50608 45574
rect 50638 45880 50694 45892
rect 50638 45846 50649 45880
rect 50683 45846 50694 45880
rect 50638 45812 50694 45846
rect 50638 45778 50649 45812
rect 50683 45778 50694 45812
rect 50638 45744 50694 45778
rect 50638 45710 50649 45744
rect 50683 45710 50694 45744
rect 50638 45676 50694 45710
rect 50638 45642 50649 45676
rect 50683 45642 50694 45676
rect 50638 45608 50694 45642
rect 50638 45574 50649 45608
rect 50683 45574 50694 45608
rect 50638 45562 50694 45574
rect 59666 45880 59722 45892
rect 59666 45846 59677 45880
rect 59711 45846 59722 45880
rect 59666 45812 59722 45846
rect 59666 45778 59677 45812
rect 59711 45778 59722 45812
rect 59666 45744 59722 45778
rect 59666 45710 59677 45744
rect 59711 45710 59722 45744
rect 59666 45676 59722 45710
rect 59666 45642 59677 45676
rect 59711 45642 59722 45676
rect 59666 45608 59722 45642
rect 59666 45574 59677 45608
rect 59711 45574 59722 45608
rect 59666 45562 59722 45574
rect 59752 45880 59808 45892
rect 59752 45846 59763 45880
rect 59797 45846 59808 45880
rect 59752 45812 59808 45846
rect 59752 45778 59763 45812
rect 59797 45778 59808 45812
rect 59752 45744 59808 45778
rect 59752 45710 59763 45744
rect 59797 45710 59808 45744
rect 59752 45676 59808 45710
rect 59752 45642 59763 45676
rect 59797 45642 59808 45676
rect 59752 45608 59808 45642
rect 59752 45574 59763 45608
rect 59797 45574 59808 45608
rect 59752 45562 59808 45574
rect 59838 45880 59894 45892
rect 59838 45846 59849 45880
rect 59883 45846 59894 45880
rect 59838 45812 59894 45846
rect 59838 45778 59849 45812
rect 59883 45778 59894 45812
rect 59838 45744 59894 45778
rect 59838 45710 59849 45744
rect 59883 45710 59894 45744
rect 59838 45676 59894 45710
rect 59838 45642 59849 45676
rect 59883 45642 59894 45676
rect 59838 45608 59894 45642
rect 59838 45574 59849 45608
rect 59883 45574 59894 45608
rect 59838 45562 59894 45574
rect 68866 45880 68922 45892
rect 68866 45846 68877 45880
rect 68911 45846 68922 45880
rect 68866 45812 68922 45846
rect 68866 45778 68877 45812
rect 68911 45778 68922 45812
rect 68866 45744 68922 45778
rect 68866 45710 68877 45744
rect 68911 45710 68922 45744
rect 68866 45676 68922 45710
rect 68866 45642 68877 45676
rect 68911 45642 68922 45676
rect 68866 45608 68922 45642
rect 68866 45574 68877 45608
rect 68911 45574 68922 45608
rect 68866 45562 68922 45574
rect 68952 45880 69008 45892
rect 68952 45846 68963 45880
rect 68997 45846 69008 45880
rect 68952 45812 69008 45846
rect 68952 45778 68963 45812
rect 68997 45778 69008 45812
rect 68952 45744 69008 45778
rect 68952 45710 68963 45744
rect 68997 45710 69008 45744
rect 68952 45676 69008 45710
rect 68952 45642 68963 45676
rect 68997 45642 69008 45676
rect 68952 45608 69008 45642
rect 68952 45574 68963 45608
rect 68997 45574 69008 45608
rect 68952 45562 69008 45574
rect 69038 45880 69094 45892
rect 69038 45846 69049 45880
rect 69083 45846 69094 45880
rect 69038 45812 69094 45846
rect 69038 45778 69049 45812
rect 69083 45778 69094 45812
rect 69038 45744 69094 45778
rect 69038 45710 69049 45744
rect 69083 45710 69094 45744
rect 69038 45676 69094 45710
rect 69038 45642 69049 45676
rect 69083 45642 69094 45676
rect 69038 45608 69094 45642
rect 69038 45574 69049 45608
rect 69083 45574 69094 45608
rect 69038 45562 69094 45574
rect -436 45254 -378 45266
rect -436 44978 -424 45254
rect -390 44978 -378 45254
rect -436 44966 -378 44978
rect -348 45254 -290 45266
rect -348 44978 -336 45254
rect -302 44978 -290 45254
rect -348 44966 -290 44978
rect 4466 36000 4522 36012
rect 4466 35966 4477 36000
rect 4511 35966 4522 36000
rect 4466 35932 4522 35966
rect 4466 35898 4477 35932
rect 4511 35898 4522 35932
rect 4466 35864 4522 35898
rect 4466 35830 4477 35864
rect 4511 35830 4522 35864
rect 4466 35796 4522 35830
rect 4466 35762 4477 35796
rect 4511 35762 4522 35796
rect 4466 35728 4522 35762
rect 4466 35694 4477 35728
rect 4511 35694 4522 35728
rect 4466 35682 4522 35694
rect 4552 36000 4608 36012
rect 4552 35966 4563 36000
rect 4597 35966 4608 36000
rect 4552 35932 4608 35966
rect 4552 35898 4563 35932
rect 4597 35898 4608 35932
rect 4552 35864 4608 35898
rect 4552 35830 4563 35864
rect 4597 35830 4608 35864
rect 4552 35796 4608 35830
rect 4552 35762 4563 35796
rect 4597 35762 4608 35796
rect 4552 35728 4608 35762
rect 4552 35694 4563 35728
rect 4597 35694 4608 35728
rect 4552 35682 4608 35694
rect 4638 36000 4694 36012
rect 4638 35966 4649 36000
rect 4683 35966 4694 36000
rect 4638 35932 4694 35966
rect 4638 35898 4649 35932
rect 4683 35898 4694 35932
rect 4638 35864 4694 35898
rect 4638 35830 4649 35864
rect 4683 35830 4694 35864
rect 4638 35796 4694 35830
rect 4638 35762 4649 35796
rect 4683 35762 4694 35796
rect 4638 35728 4694 35762
rect 4638 35694 4649 35728
rect 4683 35694 4694 35728
rect 4638 35682 4694 35694
rect 13666 36000 13722 36012
rect 13666 35966 13677 36000
rect 13711 35966 13722 36000
rect 13666 35932 13722 35966
rect 13666 35898 13677 35932
rect 13711 35898 13722 35932
rect 13666 35864 13722 35898
rect 13666 35830 13677 35864
rect 13711 35830 13722 35864
rect 13666 35796 13722 35830
rect 13666 35762 13677 35796
rect 13711 35762 13722 35796
rect 13666 35728 13722 35762
rect 13666 35694 13677 35728
rect 13711 35694 13722 35728
rect 13666 35682 13722 35694
rect 13752 36000 13808 36012
rect 13752 35966 13763 36000
rect 13797 35966 13808 36000
rect 13752 35932 13808 35966
rect 13752 35898 13763 35932
rect 13797 35898 13808 35932
rect 13752 35864 13808 35898
rect 13752 35830 13763 35864
rect 13797 35830 13808 35864
rect 13752 35796 13808 35830
rect 13752 35762 13763 35796
rect 13797 35762 13808 35796
rect 13752 35728 13808 35762
rect 13752 35694 13763 35728
rect 13797 35694 13808 35728
rect 13752 35682 13808 35694
rect 13838 36000 13894 36012
rect 13838 35966 13849 36000
rect 13883 35966 13894 36000
rect 13838 35932 13894 35966
rect 13838 35898 13849 35932
rect 13883 35898 13894 35932
rect 13838 35864 13894 35898
rect 13838 35830 13849 35864
rect 13883 35830 13894 35864
rect 13838 35796 13894 35830
rect 13838 35762 13849 35796
rect 13883 35762 13894 35796
rect 13838 35728 13894 35762
rect 13838 35694 13849 35728
rect 13883 35694 13894 35728
rect 13838 35682 13894 35694
rect 22866 36000 22922 36012
rect 22866 35966 22877 36000
rect 22911 35966 22922 36000
rect 22866 35932 22922 35966
rect 22866 35898 22877 35932
rect 22911 35898 22922 35932
rect 22866 35864 22922 35898
rect 22866 35830 22877 35864
rect 22911 35830 22922 35864
rect 22866 35796 22922 35830
rect 22866 35762 22877 35796
rect 22911 35762 22922 35796
rect 22866 35728 22922 35762
rect 22866 35694 22877 35728
rect 22911 35694 22922 35728
rect 22866 35682 22922 35694
rect 22952 36000 23008 36012
rect 22952 35966 22963 36000
rect 22997 35966 23008 36000
rect 22952 35932 23008 35966
rect 22952 35898 22963 35932
rect 22997 35898 23008 35932
rect 22952 35864 23008 35898
rect 22952 35830 22963 35864
rect 22997 35830 23008 35864
rect 22952 35796 23008 35830
rect 22952 35762 22963 35796
rect 22997 35762 23008 35796
rect 22952 35728 23008 35762
rect 22952 35694 22963 35728
rect 22997 35694 23008 35728
rect 22952 35682 23008 35694
rect 23038 36000 23094 36012
rect 23038 35966 23049 36000
rect 23083 35966 23094 36000
rect 23038 35932 23094 35966
rect 23038 35898 23049 35932
rect 23083 35898 23094 35932
rect 23038 35864 23094 35898
rect 23038 35830 23049 35864
rect 23083 35830 23094 35864
rect 23038 35796 23094 35830
rect 23038 35762 23049 35796
rect 23083 35762 23094 35796
rect 23038 35728 23094 35762
rect 23038 35694 23049 35728
rect 23083 35694 23094 35728
rect 23038 35682 23094 35694
rect 32066 36000 32122 36012
rect 32066 35966 32077 36000
rect 32111 35966 32122 36000
rect 32066 35932 32122 35966
rect 32066 35898 32077 35932
rect 32111 35898 32122 35932
rect 32066 35864 32122 35898
rect 32066 35830 32077 35864
rect 32111 35830 32122 35864
rect 32066 35796 32122 35830
rect 32066 35762 32077 35796
rect 32111 35762 32122 35796
rect 32066 35728 32122 35762
rect 32066 35694 32077 35728
rect 32111 35694 32122 35728
rect 32066 35682 32122 35694
rect 32152 36000 32208 36012
rect 32152 35966 32163 36000
rect 32197 35966 32208 36000
rect 32152 35932 32208 35966
rect 32152 35898 32163 35932
rect 32197 35898 32208 35932
rect 32152 35864 32208 35898
rect 32152 35830 32163 35864
rect 32197 35830 32208 35864
rect 32152 35796 32208 35830
rect 32152 35762 32163 35796
rect 32197 35762 32208 35796
rect 32152 35728 32208 35762
rect 32152 35694 32163 35728
rect 32197 35694 32208 35728
rect 32152 35682 32208 35694
rect 32238 36000 32294 36012
rect 32238 35966 32249 36000
rect 32283 35966 32294 36000
rect 32238 35932 32294 35966
rect 32238 35898 32249 35932
rect 32283 35898 32294 35932
rect 32238 35864 32294 35898
rect 32238 35830 32249 35864
rect 32283 35830 32294 35864
rect 32238 35796 32294 35830
rect 32238 35762 32249 35796
rect 32283 35762 32294 35796
rect 32238 35728 32294 35762
rect 32238 35694 32249 35728
rect 32283 35694 32294 35728
rect 32238 35682 32294 35694
rect 41266 36000 41322 36012
rect 41266 35966 41277 36000
rect 41311 35966 41322 36000
rect 41266 35932 41322 35966
rect 41266 35898 41277 35932
rect 41311 35898 41322 35932
rect 41266 35864 41322 35898
rect 41266 35830 41277 35864
rect 41311 35830 41322 35864
rect 41266 35796 41322 35830
rect 41266 35762 41277 35796
rect 41311 35762 41322 35796
rect 41266 35728 41322 35762
rect 41266 35694 41277 35728
rect 41311 35694 41322 35728
rect 41266 35682 41322 35694
rect 41352 36000 41408 36012
rect 41352 35966 41363 36000
rect 41397 35966 41408 36000
rect 41352 35932 41408 35966
rect 41352 35898 41363 35932
rect 41397 35898 41408 35932
rect 41352 35864 41408 35898
rect 41352 35830 41363 35864
rect 41397 35830 41408 35864
rect 41352 35796 41408 35830
rect 41352 35762 41363 35796
rect 41397 35762 41408 35796
rect 41352 35728 41408 35762
rect 41352 35694 41363 35728
rect 41397 35694 41408 35728
rect 41352 35682 41408 35694
rect 41438 36000 41494 36012
rect 41438 35966 41449 36000
rect 41483 35966 41494 36000
rect 41438 35932 41494 35966
rect 41438 35898 41449 35932
rect 41483 35898 41494 35932
rect 41438 35864 41494 35898
rect 41438 35830 41449 35864
rect 41483 35830 41494 35864
rect 41438 35796 41494 35830
rect 41438 35762 41449 35796
rect 41483 35762 41494 35796
rect 41438 35728 41494 35762
rect 41438 35694 41449 35728
rect 41483 35694 41494 35728
rect 41438 35682 41494 35694
rect 50466 36000 50522 36012
rect 50466 35966 50477 36000
rect 50511 35966 50522 36000
rect 50466 35932 50522 35966
rect 50466 35898 50477 35932
rect 50511 35898 50522 35932
rect 50466 35864 50522 35898
rect 50466 35830 50477 35864
rect 50511 35830 50522 35864
rect 50466 35796 50522 35830
rect 50466 35762 50477 35796
rect 50511 35762 50522 35796
rect 50466 35728 50522 35762
rect 50466 35694 50477 35728
rect 50511 35694 50522 35728
rect 50466 35682 50522 35694
rect 50552 36000 50608 36012
rect 50552 35966 50563 36000
rect 50597 35966 50608 36000
rect 50552 35932 50608 35966
rect 50552 35898 50563 35932
rect 50597 35898 50608 35932
rect 50552 35864 50608 35898
rect 50552 35830 50563 35864
rect 50597 35830 50608 35864
rect 50552 35796 50608 35830
rect 50552 35762 50563 35796
rect 50597 35762 50608 35796
rect 50552 35728 50608 35762
rect 50552 35694 50563 35728
rect 50597 35694 50608 35728
rect 50552 35682 50608 35694
rect 50638 36000 50694 36012
rect 50638 35966 50649 36000
rect 50683 35966 50694 36000
rect 50638 35932 50694 35966
rect 50638 35898 50649 35932
rect 50683 35898 50694 35932
rect 50638 35864 50694 35898
rect 50638 35830 50649 35864
rect 50683 35830 50694 35864
rect 50638 35796 50694 35830
rect 50638 35762 50649 35796
rect 50683 35762 50694 35796
rect 50638 35728 50694 35762
rect 50638 35694 50649 35728
rect 50683 35694 50694 35728
rect 50638 35682 50694 35694
rect 59666 36000 59722 36012
rect 59666 35966 59677 36000
rect 59711 35966 59722 36000
rect 59666 35932 59722 35966
rect 59666 35898 59677 35932
rect 59711 35898 59722 35932
rect 59666 35864 59722 35898
rect 59666 35830 59677 35864
rect 59711 35830 59722 35864
rect 59666 35796 59722 35830
rect 59666 35762 59677 35796
rect 59711 35762 59722 35796
rect 59666 35728 59722 35762
rect 59666 35694 59677 35728
rect 59711 35694 59722 35728
rect 59666 35682 59722 35694
rect 59752 36000 59808 36012
rect 59752 35966 59763 36000
rect 59797 35966 59808 36000
rect 59752 35932 59808 35966
rect 59752 35898 59763 35932
rect 59797 35898 59808 35932
rect 59752 35864 59808 35898
rect 59752 35830 59763 35864
rect 59797 35830 59808 35864
rect 59752 35796 59808 35830
rect 59752 35762 59763 35796
rect 59797 35762 59808 35796
rect 59752 35728 59808 35762
rect 59752 35694 59763 35728
rect 59797 35694 59808 35728
rect 59752 35682 59808 35694
rect 59838 36000 59894 36012
rect 59838 35966 59849 36000
rect 59883 35966 59894 36000
rect 59838 35932 59894 35966
rect 59838 35898 59849 35932
rect 59883 35898 59894 35932
rect 59838 35864 59894 35898
rect 59838 35830 59849 35864
rect 59883 35830 59894 35864
rect 59838 35796 59894 35830
rect 59838 35762 59849 35796
rect 59883 35762 59894 35796
rect 59838 35728 59894 35762
rect 59838 35694 59849 35728
rect 59883 35694 59894 35728
rect 59838 35682 59894 35694
rect 68866 36000 68922 36012
rect 68866 35966 68877 36000
rect 68911 35966 68922 36000
rect 68866 35932 68922 35966
rect 68866 35898 68877 35932
rect 68911 35898 68922 35932
rect 68866 35864 68922 35898
rect 68866 35830 68877 35864
rect 68911 35830 68922 35864
rect 68866 35796 68922 35830
rect 68866 35762 68877 35796
rect 68911 35762 68922 35796
rect 68866 35728 68922 35762
rect 68866 35694 68877 35728
rect 68911 35694 68922 35728
rect 68866 35682 68922 35694
rect 68952 36000 69008 36012
rect 68952 35966 68963 36000
rect 68997 35966 69008 36000
rect 68952 35932 69008 35966
rect 68952 35898 68963 35932
rect 68997 35898 69008 35932
rect 68952 35864 69008 35898
rect 68952 35830 68963 35864
rect 68997 35830 69008 35864
rect 68952 35796 69008 35830
rect 68952 35762 68963 35796
rect 68997 35762 69008 35796
rect 68952 35728 69008 35762
rect 68952 35694 68963 35728
rect 68997 35694 69008 35728
rect 68952 35682 69008 35694
rect 69038 36000 69094 36012
rect 69038 35966 69049 36000
rect 69083 35966 69094 36000
rect 69038 35932 69094 35966
rect 69038 35898 69049 35932
rect 69083 35898 69094 35932
rect 69038 35864 69094 35898
rect 69038 35830 69049 35864
rect 69083 35830 69094 35864
rect 69038 35796 69094 35830
rect 69038 35762 69049 35796
rect 69083 35762 69094 35796
rect 69038 35728 69094 35762
rect 69038 35694 69049 35728
rect 69083 35694 69094 35728
rect 69038 35682 69094 35694
rect 4466 26120 4522 26132
rect 4466 26086 4477 26120
rect 4511 26086 4522 26120
rect 4466 26052 4522 26086
rect 4466 26018 4477 26052
rect 4511 26018 4522 26052
rect 4466 25984 4522 26018
rect 4466 25950 4477 25984
rect 4511 25950 4522 25984
rect 4466 25916 4522 25950
rect 4466 25882 4477 25916
rect 4511 25882 4522 25916
rect 4466 25848 4522 25882
rect 4466 25814 4477 25848
rect 4511 25814 4522 25848
rect 4466 25802 4522 25814
rect 4552 26120 4608 26132
rect 4552 26086 4563 26120
rect 4597 26086 4608 26120
rect 4552 26052 4608 26086
rect 4552 26018 4563 26052
rect 4597 26018 4608 26052
rect 4552 25984 4608 26018
rect 4552 25950 4563 25984
rect 4597 25950 4608 25984
rect 4552 25916 4608 25950
rect 4552 25882 4563 25916
rect 4597 25882 4608 25916
rect 4552 25848 4608 25882
rect 4552 25814 4563 25848
rect 4597 25814 4608 25848
rect 4552 25802 4608 25814
rect 4638 26120 4694 26132
rect 4638 26086 4649 26120
rect 4683 26086 4694 26120
rect 4638 26052 4694 26086
rect 4638 26018 4649 26052
rect 4683 26018 4694 26052
rect 4638 25984 4694 26018
rect 4638 25950 4649 25984
rect 4683 25950 4694 25984
rect 4638 25916 4694 25950
rect 4638 25882 4649 25916
rect 4683 25882 4694 25916
rect 4638 25848 4694 25882
rect 4638 25814 4649 25848
rect 4683 25814 4694 25848
rect 4638 25802 4694 25814
rect 13666 26120 13722 26132
rect 13666 26086 13677 26120
rect 13711 26086 13722 26120
rect 13666 26052 13722 26086
rect 13666 26018 13677 26052
rect 13711 26018 13722 26052
rect 13666 25984 13722 26018
rect 13666 25950 13677 25984
rect 13711 25950 13722 25984
rect 13666 25916 13722 25950
rect 13666 25882 13677 25916
rect 13711 25882 13722 25916
rect 13666 25848 13722 25882
rect 13666 25814 13677 25848
rect 13711 25814 13722 25848
rect 13666 25802 13722 25814
rect 13752 26120 13808 26132
rect 13752 26086 13763 26120
rect 13797 26086 13808 26120
rect 13752 26052 13808 26086
rect 13752 26018 13763 26052
rect 13797 26018 13808 26052
rect 13752 25984 13808 26018
rect 13752 25950 13763 25984
rect 13797 25950 13808 25984
rect 13752 25916 13808 25950
rect 13752 25882 13763 25916
rect 13797 25882 13808 25916
rect 13752 25848 13808 25882
rect 13752 25814 13763 25848
rect 13797 25814 13808 25848
rect 13752 25802 13808 25814
rect 13838 26120 13894 26132
rect 13838 26086 13849 26120
rect 13883 26086 13894 26120
rect 13838 26052 13894 26086
rect 13838 26018 13849 26052
rect 13883 26018 13894 26052
rect 13838 25984 13894 26018
rect 13838 25950 13849 25984
rect 13883 25950 13894 25984
rect 13838 25916 13894 25950
rect 13838 25882 13849 25916
rect 13883 25882 13894 25916
rect 13838 25848 13894 25882
rect 13838 25814 13849 25848
rect 13883 25814 13894 25848
rect 13838 25802 13894 25814
rect 22866 26120 22922 26132
rect 22866 26086 22877 26120
rect 22911 26086 22922 26120
rect 22866 26052 22922 26086
rect 22866 26018 22877 26052
rect 22911 26018 22922 26052
rect 22866 25984 22922 26018
rect 22866 25950 22877 25984
rect 22911 25950 22922 25984
rect 22866 25916 22922 25950
rect 22866 25882 22877 25916
rect 22911 25882 22922 25916
rect 22866 25848 22922 25882
rect 22866 25814 22877 25848
rect 22911 25814 22922 25848
rect 22866 25802 22922 25814
rect 22952 26120 23008 26132
rect 22952 26086 22963 26120
rect 22997 26086 23008 26120
rect 22952 26052 23008 26086
rect 22952 26018 22963 26052
rect 22997 26018 23008 26052
rect 22952 25984 23008 26018
rect 22952 25950 22963 25984
rect 22997 25950 23008 25984
rect 22952 25916 23008 25950
rect 22952 25882 22963 25916
rect 22997 25882 23008 25916
rect 22952 25848 23008 25882
rect 22952 25814 22963 25848
rect 22997 25814 23008 25848
rect 22952 25802 23008 25814
rect 23038 26120 23094 26132
rect 23038 26086 23049 26120
rect 23083 26086 23094 26120
rect 23038 26052 23094 26086
rect 23038 26018 23049 26052
rect 23083 26018 23094 26052
rect 23038 25984 23094 26018
rect 23038 25950 23049 25984
rect 23083 25950 23094 25984
rect 23038 25916 23094 25950
rect 23038 25882 23049 25916
rect 23083 25882 23094 25916
rect 23038 25848 23094 25882
rect 23038 25814 23049 25848
rect 23083 25814 23094 25848
rect 23038 25802 23094 25814
rect 32066 26120 32122 26132
rect 32066 26086 32077 26120
rect 32111 26086 32122 26120
rect 32066 26052 32122 26086
rect 32066 26018 32077 26052
rect 32111 26018 32122 26052
rect 32066 25984 32122 26018
rect 32066 25950 32077 25984
rect 32111 25950 32122 25984
rect 32066 25916 32122 25950
rect 32066 25882 32077 25916
rect 32111 25882 32122 25916
rect 32066 25848 32122 25882
rect 32066 25814 32077 25848
rect 32111 25814 32122 25848
rect 32066 25802 32122 25814
rect 32152 26120 32208 26132
rect 32152 26086 32163 26120
rect 32197 26086 32208 26120
rect 32152 26052 32208 26086
rect 32152 26018 32163 26052
rect 32197 26018 32208 26052
rect 32152 25984 32208 26018
rect 32152 25950 32163 25984
rect 32197 25950 32208 25984
rect 32152 25916 32208 25950
rect 32152 25882 32163 25916
rect 32197 25882 32208 25916
rect 32152 25848 32208 25882
rect 32152 25814 32163 25848
rect 32197 25814 32208 25848
rect 32152 25802 32208 25814
rect 32238 26120 32294 26132
rect 32238 26086 32249 26120
rect 32283 26086 32294 26120
rect 32238 26052 32294 26086
rect 32238 26018 32249 26052
rect 32283 26018 32294 26052
rect 32238 25984 32294 26018
rect 32238 25950 32249 25984
rect 32283 25950 32294 25984
rect 32238 25916 32294 25950
rect 32238 25882 32249 25916
rect 32283 25882 32294 25916
rect 32238 25848 32294 25882
rect 32238 25814 32249 25848
rect 32283 25814 32294 25848
rect 32238 25802 32294 25814
rect 41266 26120 41322 26132
rect 41266 26086 41277 26120
rect 41311 26086 41322 26120
rect 41266 26052 41322 26086
rect 41266 26018 41277 26052
rect 41311 26018 41322 26052
rect 41266 25984 41322 26018
rect 41266 25950 41277 25984
rect 41311 25950 41322 25984
rect 41266 25916 41322 25950
rect 41266 25882 41277 25916
rect 41311 25882 41322 25916
rect 41266 25848 41322 25882
rect 41266 25814 41277 25848
rect 41311 25814 41322 25848
rect 41266 25802 41322 25814
rect 41352 26120 41408 26132
rect 41352 26086 41363 26120
rect 41397 26086 41408 26120
rect 41352 26052 41408 26086
rect 41352 26018 41363 26052
rect 41397 26018 41408 26052
rect 41352 25984 41408 26018
rect 41352 25950 41363 25984
rect 41397 25950 41408 25984
rect 41352 25916 41408 25950
rect 41352 25882 41363 25916
rect 41397 25882 41408 25916
rect 41352 25848 41408 25882
rect 41352 25814 41363 25848
rect 41397 25814 41408 25848
rect 41352 25802 41408 25814
rect 41438 26120 41494 26132
rect 41438 26086 41449 26120
rect 41483 26086 41494 26120
rect 41438 26052 41494 26086
rect 41438 26018 41449 26052
rect 41483 26018 41494 26052
rect 41438 25984 41494 26018
rect 41438 25950 41449 25984
rect 41483 25950 41494 25984
rect 41438 25916 41494 25950
rect 41438 25882 41449 25916
rect 41483 25882 41494 25916
rect 41438 25848 41494 25882
rect 41438 25814 41449 25848
rect 41483 25814 41494 25848
rect 41438 25802 41494 25814
rect 50466 26120 50522 26132
rect 50466 26086 50477 26120
rect 50511 26086 50522 26120
rect 50466 26052 50522 26086
rect 50466 26018 50477 26052
rect 50511 26018 50522 26052
rect 50466 25984 50522 26018
rect 50466 25950 50477 25984
rect 50511 25950 50522 25984
rect 50466 25916 50522 25950
rect 50466 25882 50477 25916
rect 50511 25882 50522 25916
rect 50466 25848 50522 25882
rect 50466 25814 50477 25848
rect 50511 25814 50522 25848
rect 50466 25802 50522 25814
rect 50552 26120 50608 26132
rect 50552 26086 50563 26120
rect 50597 26086 50608 26120
rect 50552 26052 50608 26086
rect 50552 26018 50563 26052
rect 50597 26018 50608 26052
rect 50552 25984 50608 26018
rect 50552 25950 50563 25984
rect 50597 25950 50608 25984
rect 50552 25916 50608 25950
rect 50552 25882 50563 25916
rect 50597 25882 50608 25916
rect 50552 25848 50608 25882
rect 50552 25814 50563 25848
rect 50597 25814 50608 25848
rect 50552 25802 50608 25814
rect 50638 26120 50694 26132
rect 50638 26086 50649 26120
rect 50683 26086 50694 26120
rect 50638 26052 50694 26086
rect 50638 26018 50649 26052
rect 50683 26018 50694 26052
rect 50638 25984 50694 26018
rect 50638 25950 50649 25984
rect 50683 25950 50694 25984
rect 50638 25916 50694 25950
rect 50638 25882 50649 25916
rect 50683 25882 50694 25916
rect 50638 25848 50694 25882
rect 50638 25814 50649 25848
rect 50683 25814 50694 25848
rect 50638 25802 50694 25814
rect 59666 26120 59722 26132
rect 59666 26086 59677 26120
rect 59711 26086 59722 26120
rect 59666 26052 59722 26086
rect 59666 26018 59677 26052
rect 59711 26018 59722 26052
rect 59666 25984 59722 26018
rect 59666 25950 59677 25984
rect 59711 25950 59722 25984
rect 59666 25916 59722 25950
rect 59666 25882 59677 25916
rect 59711 25882 59722 25916
rect 59666 25848 59722 25882
rect 59666 25814 59677 25848
rect 59711 25814 59722 25848
rect 59666 25802 59722 25814
rect 59752 26120 59808 26132
rect 59752 26086 59763 26120
rect 59797 26086 59808 26120
rect 59752 26052 59808 26086
rect 59752 26018 59763 26052
rect 59797 26018 59808 26052
rect 59752 25984 59808 26018
rect 59752 25950 59763 25984
rect 59797 25950 59808 25984
rect 59752 25916 59808 25950
rect 59752 25882 59763 25916
rect 59797 25882 59808 25916
rect 59752 25848 59808 25882
rect 59752 25814 59763 25848
rect 59797 25814 59808 25848
rect 59752 25802 59808 25814
rect 59838 26120 59894 26132
rect 59838 26086 59849 26120
rect 59883 26086 59894 26120
rect 59838 26052 59894 26086
rect 59838 26018 59849 26052
rect 59883 26018 59894 26052
rect 59838 25984 59894 26018
rect 59838 25950 59849 25984
rect 59883 25950 59894 25984
rect 59838 25916 59894 25950
rect 59838 25882 59849 25916
rect 59883 25882 59894 25916
rect 59838 25848 59894 25882
rect 59838 25814 59849 25848
rect 59883 25814 59894 25848
rect 59838 25802 59894 25814
rect 68866 26120 68922 26132
rect 68866 26086 68877 26120
rect 68911 26086 68922 26120
rect 68866 26052 68922 26086
rect 68866 26018 68877 26052
rect 68911 26018 68922 26052
rect 68866 25984 68922 26018
rect 68866 25950 68877 25984
rect 68911 25950 68922 25984
rect 68866 25916 68922 25950
rect 68866 25882 68877 25916
rect 68911 25882 68922 25916
rect 68866 25848 68922 25882
rect 68866 25814 68877 25848
rect 68911 25814 68922 25848
rect 68866 25802 68922 25814
rect 68952 26120 69008 26132
rect 68952 26086 68963 26120
rect 68997 26086 69008 26120
rect 68952 26052 69008 26086
rect 68952 26018 68963 26052
rect 68997 26018 69008 26052
rect 68952 25984 69008 26018
rect 68952 25950 68963 25984
rect 68997 25950 69008 25984
rect 68952 25916 69008 25950
rect 68952 25882 68963 25916
rect 68997 25882 69008 25916
rect 68952 25848 69008 25882
rect 68952 25814 68963 25848
rect 68997 25814 69008 25848
rect 68952 25802 69008 25814
rect 69038 26120 69094 26132
rect 69038 26086 69049 26120
rect 69083 26086 69094 26120
rect 69038 26052 69094 26086
rect 69038 26018 69049 26052
rect 69083 26018 69094 26052
rect 69038 25984 69094 26018
rect 69038 25950 69049 25984
rect 69083 25950 69094 25984
rect 69038 25916 69094 25950
rect 69038 25882 69049 25916
rect 69083 25882 69094 25916
rect 69038 25848 69094 25882
rect 69038 25814 69049 25848
rect 69083 25814 69094 25848
rect 69038 25802 69094 25814
rect 4466 16240 4522 16252
rect 4466 16206 4477 16240
rect 4511 16206 4522 16240
rect 4466 16172 4522 16206
rect 4466 16138 4477 16172
rect 4511 16138 4522 16172
rect 4466 16104 4522 16138
rect 4466 16070 4477 16104
rect 4511 16070 4522 16104
rect 4466 16036 4522 16070
rect 4466 16002 4477 16036
rect 4511 16002 4522 16036
rect 4466 15968 4522 16002
rect 4466 15934 4477 15968
rect 4511 15934 4522 15968
rect 4466 15922 4522 15934
rect 4552 16240 4608 16252
rect 4552 16206 4563 16240
rect 4597 16206 4608 16240
rect 4552 16172 4608 16206
rect 4552 16138 4563 16172
rect 4597 16138 4608 16172
rect 4552 16104 4608 16138
rect 4552 16070 4563 16104
rect 4597 16070 4608 16104
rect 4552 16036 4608 16070
rect 4552 16002 4563 16036
rect 4597 16002 4608 16036
rect 4552 15968 4608 16002
rect 4552 15934 4563 15968
rect 4597 15934 4608 15968
rect 4552 15922 4608 15934
rect 4638 16240 4694 16252
rect 4638 16206 4649 16240
rect 4683 16206 4694 16240
rect 4638 16172 4694 16206
rect 4638 16138 4649 16172
rect 4683 16138 4694 16172
rect 4638 16104 4694 16138
rect 4638 16070 4649 16104
rect 4683 16070 4694 16104
rect 4638 16036 4694 16070
rect 4638 16002 4649 16036
rect 4683 16002 4694 16036
rect 4638 15968 4694 16002
rect 4638 15934 4649 15968
rect 4683 15934 4694 15968
rect 4638 15922 4694 15934
rect 13666 16240 13722 16252
rect 13666 16206 13677 16240
rect 13711 16206 13722 16240
rect 13666 16172 13722 16206
rect 13666 16138 13677 16172
rect 13711 16138 13722 16172
rect 13666 16104 13722 16138
rect 13666 16070 13677 16104
rect 13711 16070 13722 16104
rect 13666 16036 13722 16070
rect 13666 16002 13677 16036
rect 13711 16002 13722 16036
rect 13666 15968 13722 16002
rect 13666 15934 13677 15968
rect 13711 15934 13722 15968
rect 13666 15922 13722 15934
rect 13752 16240 13808 16252
rect 13752 16206 13763 16240
rect 13797 16206 13808 16240
rect 13752 16172 13808 16206
rect 13752 16138 13763 16172
rect 13797 16138 13808 16172
rect 13752 16104 13808 16138
rect 13752 16070 13763 16104
rect 13797 16070 13808 16104
rect 13752 16036 13808 16070
rect 13752 16002 13763 16036
rect 13797 16002 13808 16036
rect 13752 15968 13808 16002
rect 13752 15934 13763 15968
rect 13797 15934 13808 15968
rect 13752 15922 13808 15934
rect 13838 16240 13894 16252
rect 13838 16206 13849 16240
rect 13883 16206 13894 16240
rect 13838 16172 13894 16206
rect 13838 16138 13849 16172
rect 13883 16138 13894 16172
rect 13838 16104 13894 16138
rect 13838 16070 13849 16104
rect 13883 16070 13894 16104
rect 13838 16036 13894 16070
rect 13838 16002 13849 16036
rect 13883 16002 13894 16036
rect 13838 15968 13894 16002
rect 13838 15934 13849 15968
rect 13883 15934 13894 15968
rect 13838 15922 13894 15934
rect 22866 16240 22922 16252
rect 22866 16206 22877 16240
rect 22911 16206 22922 16240
rect 22866 16172 22922 16206
rect 22866 16138 22877 16172
rect 22911 16138 22922 16172
rect 22866 16104 22922 16138
rect 22866 16070 22877 16104
rect 22911 16070 22922 16104
rect 22866 16036 22922 16070
rect 22866 16002 22877 16036
rect 22911 16002 22922 16036
rect 22866 15968 22922 16002
rect 22866 15934 22877 15968
rect 22911 15934 22922 15968
rect 22866 15922 22922 15934
rect 22952 16240 23008 16252
rect 22952 16206 22963 16240
rect 22997 16206 23008 16240
rect 22952 16172 23008 16206
rect 22952 16138 22963 16172
rect 22997 16138 23008 16172
rect 22952 16104 23008 16138
rect 22952 16070 22963 16104
rect 22997 16070 23008 16104
rect 22952 16036 23008 16070
rect 22952 16002 22963 16036
rect 22997 16002 23008 16036
rect 22952 15968 23008 16002
rect 22952 15934 22963 15968
rect 22997 15934 23008 15968
rect 22952 15922 23008 15934
rect 23038 16240 23094 16252
rect 23038 16206 23049 16240
rect 23083 16206 23094 16240
rect 23038 16172 23094 16206
rect 23038 16138 23049 16172
rect 23083 16138 23094 16172
rect 23038 16104 23094 16138
rect 23038 16070 23049 16104
rect 23083 16070 23094 16104
rect 23038 16036 23094 16070
rect 23038 16002 23049 16036
rect 23083 16002 23094 16036
rect 23038 15968 23094 16002
rect 23038 15934 23049 15968
rect 23083 15934 23094 15968
rect 23038 15922 23094 15934
rect 32066 16240 32122 16252
rect 32066 16206 32077 16240
rect 32111 16206 32122 16240
rect 32066 16172 32122 16206
rect 32066 16138 32077 16172
rect 32111 16138 32122 16172
rect 32066 16104 32122 16138
rect 32066 16070 32077 16104
rect 32111 16070 32122 16104
rect 32066 16036 32122 16070
rect 32066 16002 32077 16036
rect 32111 16002 32122 16036
rect 32066 15968 32122 16002
rect 32066 15934 32077 15968
rect 32111 15934 32122 15968
rect 32066 15922 32122 15934
rect 32152 16240 32208 16252
rect 32152 16206 32163 16240
rect 32197 16206 32208 16240
rect 32152 16172 32208 16206
rect 32152 16138 32163 16172
rect 32197 16138 32208 16172
rect 32152 16104 32208 16138
rect 32152 16070 32163 16104
rect 32197 16070 32208 16104
rect 32152 16036 32208 16070
rect 32152 16002 32163 16036
rect 32197 16002 32208 16036
rect 32152 15968 32208 16002
rect 32152 15934 32163 15968
rect 32197 15934 32208 15968
rect 32152 15922 32208 15934
rect 32238 16240 32294 16252
rect 32238 16206 32249 16240
rect 32283 16206 32294 16240
rect 32238 16172 32294 16206
rect 32238 16138 32249 16172
rect 32283 16138 32294 16172
rect 32238 16104 32294 16138
rect 32238 16070 32249 16104
rect 32283 16070 32294 16104
rect 32238 16036 32294 16070
rect 32238 16002 32249 16036
rect 32283 16002 32294 16036
rect 32238 15968 32294 16002
rect 32238 15934 32249 15968
rect 32283 15934 32294 15968
rect 32238 15922 32294 15934
rect 41266 16240 41322 16252
rect 41266 16206 41277 16240
rect 41311 16206 41322 16240
rect 41266 16172 41322 16206
rect 41266 16138 41277 16172
rect 41311 16138 41322 16172
rect 41266 16104 41322 16138
rect 41266 16070 41277 16104
rect 41311 16070 41322 16104
rect 41266 16036 41322 16070
rect 41266 16002 41277 16036
rect 41311 16002 41322 16036
rect 41266 15968 41322 16002
rect 41266 15934 41277 15968
rect 41311 15934 41322 15968
rect 41266 15922 41322 15934
rect 41352 16240 41408 16252
rect 41352 16206 41363 16240
rect 41397 16206 41408 16240
rect 41352 16172 41408 16206
rect 41352 16138 41363 16172
rect 41397 16138 41408 16172
rect 41352 16104 41408 16138
rect 41352 16070 41363 16104
rect 41397 16070 41408 16104
rect 41352 16036 41408 16070
rect 41352 16002 41363 16036
rect 41397 16002 41408 16036
rect 41352 15968 41408 16002
rect 41352 15934 41363 15968
rect 41397 15934 41408 15968
rect 41352 15922 41408 15934
rect 41438 16240 41494 16252
rect 41438 16206 41449 16240
rect 41483 16206 41494 16240
rect 41438 16172 41494 16206
rect 41438 16138 41449 16172
rect 41483 16138 41494 16172
rect 41438 16104 41494 16138
rect 41438 16070 41449 16104
rect 41483 16070 41494 16104
rect 41438 16036 41494 16070
rect 41438 16002 41449 16036
rect 41483 16002 41494 16036
rect 41438 15968 41494 16002
rect 41438 15934 41449 15968
rect 41483 15934 41494 15968
rect 41438 15922 41494 15934
rect 50466 16240 50522 16252
rect 50466 16206 50477 16240
rect 50511 16206 50522 16240
rect 50466 16172 50522 16206
rect 50466 16138 50477 16172
rect 50511 16138 50522 16172
rect 50466 16104 50522 16138
rect 50466 16070 50477 16104
rect 50511 16070 50522 16104
rect 50466 16036 50522 16070
rect 50466 16002 50477 16036
rect 50511 16002 50522 16036
rect 50466 15968 50522 16002
rect 50466 15934 50477 15968
rect 50511 15934 50522 15968
rect 50466 15922 50522 15934
rect 50552 16240 50608 16252
rect 50552 16206 50563 16240
rect 50597 16206 50608 16240
rect 50552 16172 50608 16206
rect 50552 16138 50563 16172
rect 50597 16138 50608 16172
rect 50552 16104 50608 16138
rect 50552 16070 50563 16104
rect 50597 16070 50608 16104
rect 50552 16036 50608 16070
rect 50552 16002 50563 16036
rect 50597 16002 50608 16036
rect 50552 15968 50608 16002
rect 50552 15934 50563 15968
rect 50597 15934 50608 15968
rect 50552 15922 50608 15934
rect 50638 16240 50694 16252
rect 50638 16206 50649 16240
rect 50683 16206 50694 16240
rect 50638 16172 50694 16206
rect 50638 16138 50649 16172
rect 50683 16138 50694 16172
rect 50638 16104 50694 16138
rect 50638 16070 50649 16104
rect 50683 16070 50694 16104
rect 50638 16036 50694 16070
rect 50638 16002 50649 16036
rect 50683 16002 50694 16036
rect 50638 15968 50694 16002
rect 50638 15934 50649 15968
rect 50683 15934 50694 15968
rect 50638 15922 50694 15934
rect 59666 16240 59722 16252
rect 59666 16206 59677 16240
rect 59711 16206 59722 16240
rect 59666 16172 59722 16206
rect 59666 16138 59677 16172
rect 59711 16138 59722 16172
rect 59666 16104 59722 16138
rect 59666 16070 59677 16104
rect 59711 16070 59722 16104
rect 59666 16036 59722 16070
rect 59666 16002 59677 16036
rect 59711 16002 59722 16036
rect 59666 15968 59722 16002
rect 59666 15934 59677 15968
rect 59711 15934 59722 15968
rect 59666 15922 59722 15934
rect 59752 16240 59808 16252
rect 59752 16206 59763 16240
rect 59797 16206 59808 16240
rect 59752 16172 59808 16206
rect 59752 16138 59763 16172
rect 59797 16138 59808 16172
rect 59752 16104 59808 16138
rect 59752 16070 59763 16104
rect 59797 16070 59808 16104
rect 59752 16036 59808 16070
rect 59752 16002 59763 16036
rect 59797 16002 59808 16036
rect 59752 15968 59808 16002
rect 59752 15934 59763 15968
rect 59797 15934 59808 15968
rect 59752 15922 59808 15934
rect 59838 16240 59894 16252
rect 59838 16206 59849 16240
rect 59883 16206 59894 16240
rect 59838 16172 59894 16206
rect 59838 16138 59849 16172
rect 59883 16138 59894 16172
rect 59838 16104 59894 16138
rect 59838 16070 59849 16104
rect 59883 16070 59894 16104
rect 59838 16036 59894 16070
rect 59838 16002 59849 16036
rect 59883 16002 59894 16036
rect 59838 15968 59894 16002
rect 59838 15934 59849 15968
rect 59883 15934 59894 15968
rect 59838 15922 59894 15934
rect 68866 16240 68922 16252
rect 68866 16206 68877 16240
rect 68911 16206 68922 16240
rect 68866 16172 68922 16206
rect 68866 16138 68877 16172
rect 68911 16138 68922 16172
rect 68866 16104 68922 16138
rect 68866 16070 68877 16104
rect 68911 16070 68922 16104
rect 68866 16036 68922 16070
rect 68866 16002 68877 16036
rect 68911 16002 68922 16036
rect 68866 15968 68922 16002
rect 68866 15934 68877 15968
rect 68911 15934 68922 15968
rect 68866 15922 68922 15934
rect 68952 16240 69008 16252
rect 68952 16206 68963 16240
rect 68997 16206 69008 16240
rect 68952 16172 69008 16206
rect 68952 16138 68963 16172
rect 68997 16138 69008 16172
rect 68952 16104 69008 16138
rect 68952 16070 68963 16104
rect 68997 16070 69008 16104
rect 68952 16036 69008 16070
rect 68952 16002 68963 16036
rect 68997 16002 69008 16036
rect 68952 15968 69008 16002
rect 68952 15934 68963 15968
rect 68997 15934 69008 15968
rect 68952 15922 69008 15934
rect 69038 16240 69094 16252
rect 69038 16206 69049 16240
rect 69083 16206 69094 16240
rect 69038 16172 69094 16206
rect 69038 16138 69049 16172
rect 69083 16138 69094 16172
rect 69038 16104 69094 16138
rect 69038 16070 69049 16104
rect 69083 16070 69094 16104
rect 69038 16036 69094 16070
rect 69038 16002 69049 16036
rect 69083 16002 69094 16036
rect 69038 15968 69094 16002
rect 69038 15934 69049 15968
rect 69083 15934 69094 15968
rect 69038 15922 69094 15934
rect 4466 6360 4522 6372
rect 4466 6326 4477 6360
rect 4511 6326 4522 6360
rect 4466 6292 4522 6326
rect 4466 6258 4477 6292
rect 4511 6258 4522 6292
rect 4466 6224 4522 6258
rect 4466 6190 4477 6224
rect 4511 6190 4522 6224
rect 4466 6156 4522 6190
rect 4466 6122 4477 6156
rect 4511 6122 4522 6156
rect 4466 6088 4522 6122
rect 4466 6054 4477 6088
rect 4511 6054 4522 6088
rect 4466 6042 4522 6054
rect 4552 6360 4608 6372
rect 4552 6326 4563 6360
rect 4597 6326 4608 6360
rect 4552 6292 4608 6326
rect 4552 6258 4563 6292
rect 4597 6258 4608 6292
rect 4552 6224 4608 6258
rect 4552 6190 4563 6224
rect 4597 6190 4608 6224
rect 4552 6156 4608 6190
rect 4552 6122 4563 6156
rect 4597 6122 4608 6156
rect 4552 6088 4608 6122
rect 4552 6054 4563 6088
rect 4597 6054 4608 6088
rect 4552 6042 4608 6054
rect 4638 6360 4694 6372
rect 4638 6326 4649 6360
rect 4683 6326 4694 6360
rect 4638 6292 4694 6326
rect 4638 6258 4649 6292
rect 4683 6258 4694 6292
rect 4638 6224 4694 6258
rect 4638 6190 4649 6224
rect 4683 6190 4694 6224
rect 4638 6156 4694 6190
rect 4638 6122 4649 6156
rect 4683 6122 4694 6156
rect 4638 6088 4694 6122
rect 4638 6054 4649 6088
rect 4683 6054 4694 6088
rect 4638 6042 4694 6054
rect 13666 6360 13722 6372
rect 13666 6326 13677 6360
rect 13711 6326 13722 6360
rect 13666 6292 13722 6326
rect 13666 6258 13677 6292
rect 13711 6258 13722 6292
rect 13666 6224 13722 6258
rect 13666 6190 13677 6224
rect 13711 6190 13722 6224
rect 13666 6156 13722 6190
rect 13666 6122 13677 6156
rect 13711 6122 13722 6156
rect 13666 6088 13722 6122
rect 13666 6054 13677 6088
rect 13711 6054 13722 6088
rect 13666 6042 13722 6054
rect 13752 6360 13808 6372
rect 13752 6326 13763 6360
rect 13797 6326 13808 6360
rect 13752 6292 13808 6326
rect 13752 6258 13763 6292
rect 13797 6258 13808 6292
rect 13752 6224 13808 6258
rect 13752 6190 13763 6224
rect 13797 6190 13808 6224
rect 13752 6156 13808 6190
rect 13752 6122 13763 6156
rect 13797 6122 13808 6156
rect 13752 6088 13808 6122
rect 13752 6054 13763 6088
rect 13797 6054 13808 6088
rect 13752 6042 13808 6054
rect 13838 6360 13894 6372
rect 13838 6326 13849 6360
rect 13883 6326 13894 6360
rect 13838 6292 13894 6326
rect 13838 6258 13849 6292
rect 13883 6258 13894 6292
rect 13838 6224 13894 6258
rect 13838 6190 13849 6224
rect 13883 6190 13894 6224
rect 13838 6156 13894 6190
rect 13838 6122 13849 6156
rect 13883 6122 13894 6156
rect 13838 6088 13894 6122
rect 13838 6054 13849 6088
rect 13883 6054 13894 6088
rect 13838 6042 13894 6054
rect 22866 6360 22922 6372
rect 22866 6326 22877 6360
rect 22911 6326 22922 6360
rect 22866 6292 22922 6326
rect 22866 6258 22877 6292
rect 22911 6258 22922 6292
rect 22866 6224 22922 6258
rect 22866 6190 22877 6224
rect 22911 6190 22922 6224
rect 22866 6156 22922 6190
rect 22866 6122 22877 6156
rect 22911 6122 22922 6156
rect 22866 6088 22922 6122
rect 22866 6054 22877 6088
rect 22911 6054 22922 6088
rect 22866 6042 22922 6054
rect 22952 6360 23008 6372
rect 22952 6326 22963 6360
rect 22997 6326 23008 6360
rect 22952 6292 23008 6326
rect 22952 6258 22963 6292
rect 22997 6258 23008 6292
rect 22952 6224 23008 6258
rect 22952 6190 22963 6224
rect 22997 6190 23008 6224
rect 22952 6156 23008 6190
rect 22952 6122 22963 6156
rect 22997 6122 23008 6156
rect 22952 6088 23008 6122
rect 22952 6054 22963 6088
rect 22997 6054 23008 6088
rect 22952 6042 23008 6054
rect 23038 6360 23094 6372
rect 23038 6326 23049 6360
rect 23083 6326 23094 6360
rect 23038 6292 23094 6326
rect 23038 6258 23049 6292
rect 23083 6258 23094 6292
rect 23038 6224 23094 6258
rect 23038 6190 23049 6224
rect 23083 6190 23094 6224
rect 23038 6156 23094 6190
rect 23038 6122 23049 6156
rect 23083 6122 23094 6156
rect 23038 6088 23094 6122
rect 23038 6054 23049 6088
rect 23083 6054 23094 6088
rect 23038 6042 23094 6054
rect 32066 6360 32122 6372
rect 32066 6326 32077 6360
rect 32111 6326 32122 6360
rect 32066 6292 32122 6326
rect 32066 6258 32077 6292
rect 32111 6258 32122 6292
rect 32066 6224 32122 6258
rect 32066 6190 32077 6224
rect 32111 6190 32122 6224
rect 32066 6156 32122 6190
rect 32066 6122 32077 6156
rect 32111 6122 32122 6156
rect 32066 6088 32122 6122
rect 32066 6054 32077 6088
rect 32111 6054 32122 6088
rect 32066 6042 32122 6054
rect 32152 6360 32208 6372
rect 32152 6326 32163 6360
rect 32197 6326 32208 6360
rect 32152 6292 32208 6326
rect 32152 6258 32163 6292
rect 32197 6258 32208 6292
rect 32152 6224 32208 6258
rect 32152 6190 32163 6224
rect 32197 6190 32208 6224
rect 32152 6156 32208 6190
rect 32152 6122 32163 6156
rect 32197 6122 32208 6156
rect 32152 6088 32208 6122
rect 32152 6054 32163 6088
rect 32197 6054 32208 6088
rect 32152 6042 32208 6054
rect 32238 6360 32294 6372
rect 32238 6326 32249 6360
rect 32283 6326 32294 6360
rect 32238 6292 32294 6326
rect 32238 6258 32249 6292
rect 32283 6258 32294 6292
rect 32238 6224 32294 6258
rect 32238 6190 32249 6224
rect 32283 6190 32294 6224
rect 32238 6156 32294 6190
rect 32238 6122 32249 6156
rect 32283 6122 32294 6156
rect 32238 6088 32294 6122
rect 32238 6054 32249 6088
rect 32283 6054 32294 6088
rect 32238 6042 32294 6054
rect 41266 6360 41322 6372
rect 41266 6326 41277 6360
rect 41311 6326 41322 6360
rect 41266 6292 41322 6326
rect 41266 6258 41277 6292
rect 41311 6258 41322 6292
rect 41266 6224 41322 6258
rect 41266 6190 41277 6224
rect 41311 6190 41322 6224
rect 41266 6156 41322 6190
rect 41266 6122 41277 6156
rect 41311 6122 41322 6156
rect 41266 6088 41322 6122
rect 41266 6054 41277 6088
rect 41311 6054 41322 6088
rect 41266 6042 41322 6054
rect 41352 6360 41408 6372
rect 41352 6326 41363 6360
rect 41397 6326 41408 6360
rect 41352 6292 41408 6326
rect 41352 6258 41363 6292
rect 41397 6258 41408 6292
rect 41352 6224 41408 6258
rect 41352 6190 41363 6224
rect 41397 6190 41408 6224
rect 41352 6156 41408 6190
rect 41352 6122 41363 6156
rect 41397 6122 41408 6156
rect 41352 6088 41408 6122
rect 41352 6054 41363 6088
rect 41397 6054 41408 6088
rect 41352 6042 41408 6054
rect 41438 6360 41494 6372
rect 41438 6326 41449 6360
rect 41483 6326 41494 6360
rect 41438 6292 41494 6326
rect 41438 6258 41449 6292
rect 41483 6258 41494 6292
rect 41438 6224 41494 6258
rect 41438 6190 41449 6224
rect 41483 6190 41494 6224
rect 41438 6156 41494 6190
rect 41438 6122 41449 6156
rect 41483 6122 41494 6156
rect 41438 6088 41494 6122
rect 41438 6054 41449 6088
rect 41483 6054 41494 6088
rect 41438 6042 41494 6054
rect 50466 6360 50522 6372
rect 50466 6326 50477 6360
rect 50511 6326 50522 6360
rect 50466 6292 50522 6326
rect 50466 6258 50477 6292
rect 50511 6258 50522 6292
rect 50466 6224 50522 6258
rect 50466 6190 50477 6224
rect 50511 6190 50522 6224
rect 50466 6156 50522 6190
rect 50466 6122 50477 6156
rect 50511 6122 50522 6156
rect 50466 6088 50522 6122
rect 50466 6054 50477 6088
rect 50511 6054 50522 6088
rect 50466 6042 50522 6054
rect 50552 6360 50608 6372
rect 50552 6326 50563 6360
rect 50597 6326 50608 6360
rect 50552 6292 50608 6326
rect 50552 6258 50563 6292
rect 50597 6258 50608 6292
rect 50552 6224 50608 6258
rect 50552 6190 50563 6224
rect 50597 6190 50608 6224
rect 50552 6156 50608 6190
rect 50552 6122 50563 6156
rect 50597 6122 50608 6156
rect 50552 6088 50608 6122
rect 50552 6054 50563 6088
rect 50597 6054 50608 6088
rect 50552 6042 50608 6054
rect 50638 6360 50694 6372
rect 50638 6326 50649 6360
rect 50683 6326 50694 6360
rect 50638 6292 50694 6326
rect 50638 6258 50649 6292
rect 50683 6258 50694 6292
rect 50638 6224 50694 6258
rect 50638 6190 50649 6224
rect 50683 6190 50694 6224
rect 50638 6156 50694 6190
rect 50638 6122 50649 6156
rect 50683 6122 50694 6156
rect 50638 6088 50694 6122
rect 50638 6054 50649 6088
rect 50683 6054 50694 6088
rect 50638 6042 50694 6054
rect 59666 6360 59722 6372
rect 59666 6326 59677 6360
rect 59711 6326 59722 6360
rect 59666 6292 59722 6326
rect 59666 6258 59677 6292
rect 59711 6258 59722 6292
rect 59666 6224 59722 6258
rect 59666 6190 59677 6224
rect 59711 6190 59722 6224
rect 59666 6156 59722 6190
rect 59666 6122 59677 6156
rect 59711 6122 59722 6156
rect 59666 6088 59722 6122
rect 59666 6054 59677 6088
rect 59711 6054 59722 6088
rect 59666 6042 59722 6054
rect 59752 6360 59808 6372
rect 59752 6326 59763 6360
rect 59797 6326 59808 6360
rect 59752 6292 59808 6326
rect 59752 6258 59763 6292
rect 59797 6258 59808 6292
rect 59752 6224 59808 6258
rect 59752 6190 59763 6224
rect 59797 6190 59808 6224
rect 59752 6156 59808 6190
rect 59752 6122 59763 6156
rect 59797 6122 59808 6156
rect 59752 6088 59808 6122
rect 59752 6054 59763 6088
rect 59797 6054 59808 6088
rect 59752 6042 59808 6054
rect 59838 6360 59894 6372
rect 59838 6326 59849 6360
rect 59883 6326 59894 6360
rect 59838 6292 59894 6326
rect 59838 6258 59849 6292
rect 59883 6258 59894 6292
rect 59838 6224 59894 6258
rect 59838 6190 59849 6224
rect 59883 6190 59894 6224
rect 59838 6156 59894 6190
rect 59838 6122 59849 6156
rect 59883 6122 59894 6156
rect 59838 6088 59894 6122
rect 59838 6054 59849 6088
rect 59883 6054 59894 6088
rect 59838 6042 59894 6054
rect 68866 6360 68922 6372
rect 68866 6326 68877 6360
rect 68911 6326 68922 6360
rect 68866 6292 68922 6326
rect 68866 6258 68877 6292
rect 68911 6258 68922 6292
rect 68866 6224 68922 6258
rect 68866 6190 68877 6224
rect 68911 6190 68922 6224
rect 68866 6156 68922 6190
rect 68866 6122 68877 6156
rect 68911 6122 68922 6156
rect 68866 6088 68922 6122
rect 68866 6054 68877 6088
rect 68911 6054 68922 6088
rect 68866 6042 68922 6054
rect 68952 6360 69008 6372
rect 68952 6326 68963 6360
rect 68997 6326 69008 6360
rect 68952 6292 69008 6326
rect 68952 6258 68963 6292
rect 68997 6258 69008 6292
rect 68952 6224 69008 6258
rect 68952 6190 68963 6224
rect 68997 6190 69008 6224
rect 68952 6156 69008 6190
rect 68952 6122 68963 6156
rect 68997 6122 69008 6156
rect 68952 6088 69008 6122
rect 68952 6054 68963 6088
rect 68997 6054 69008 6088
rect 68952 6042 69008 6054
rect 69038 6360 69094 6372
rect 69038 6326 69049 6360
rect 69083 6326 69094 6360
rect 69038 6292 69094 6326
rect 69038 6258 69049 6292
rect 69083 6258 69094 6292
rect 69038 6224 69094 6258
rect 69038 6190 69049 6224
rect 69083 6190 69094 6224
rect 69038 6156 69094 6190
rect 69038 6122 69049 6156
rect 69083 6122 69094 6156
rect 69038 6088 69094 6122
rect 69038 6054 69049 6088
rect 69083 6054 69094 6088
rect 69038 6042 69094 6054
rect -436 5734 -378 5746
rect -436 5458 -424 5734
rect -390 5458 -378 5734
rect -436 5446 -378 5458
rect -348 5734 -290 5746
rect -348 5458 -336 5734
rect -302 5458 -290 5734
rect -348 5446 -290 5458
<< pdiff >>
rect -436 95384 -378 95396
rect -436 94808 -424 95384
rect -390 94808 -378 95384
rect -436 94796 -378 94808
rect -348 95384 -290 95396
rect -348 94808 -336 95384
rect -302 94808 -290 95384
rect -348 94796 -290 94808
rect -436 85504 -378 85516
rect -436 84928 -424 85504
rect -390 84928 -378 85504
rect -436 84916 -378 84928
rect -348 85504 -290 85516
rect -348 84928 -336 85504
rect -302 84928 -290 85504
rect -348 84916 -290 84928
rect -436 75624 -378 75636
rect -436 75048 -424 75624
rect -390 75048 -378 75624
rect -436 75036 -378 75048
rect -348 75624 -290 75636
rect -348 75048 -336 75624
rect -302 75048 -290 75624
rect -348 75036 -290 75048
rect -436 65744 -378 65756
rect -436 65168 -424 65744
rect -390 65168 -378 65744
rect -436 65156 -378 65168
rect -348 65744 -290 65756
rect -348 65168 -336 65744
rect -302 65168 -290 65744
rect -348 65156 -290 65168
rect -436 45984 -378 45996
rect -436 45408 -424 45984
rect -390 45408 -378 45984
rect -436 45396 -378 45408
rect -348 45984 -290 45996
rect -348 45408 -336 45984
rect -302 45408 -290 45984
rect -348 45396 -290 45408
rect -436 6464 -378 6476
rect -436 5888 -424 6464
rect -390 5888 -378 6464
rect -436 5876 -378 5888
rect -348 6464 -290 6476
rect -348 5888 -336 6464
rect -302 5888 -290 6464
rect -348 5876 -290 5888
<< ndiffc >>
rect 4477 95246 4511 95280
rect 4477 95178 4511 95212
rect 4477 95110 4511 95144
rect 4477 95042 4511 95076
rect 4477 94974 4511 95008
rect 4563 95246 4597 95280
rect 4563 95178 4597 95212
rect 4563 95110 4597 95144
rect 4563 95042 4597 95076
rect 4563 94974 4597 95008
rect 4649 95246 4683 95280
rect 4649 95178 4683 95212
rect 4649 95110 4683 95144
rect 4649 95042 4683 95076
rect 4649 94974 4683 95008
rect -424 94378 -390 94654
rect -336 94378 -302 94654
rect 4477 85366 4511 85400
rect 4477 85298 4511 85332
rect 4477 85230 4511 85264
rect 4477 85162 4511 85196
rect 4477 85094 4511 85128
rect 4563 85366 4597 85400
rect 4563 85298 4597 85332
rect 4563 85230 4597 85264
rect 4563 85162 4597 85196
rect 4563 85094 4597 85128
rect 4649 85366 4683 85400
rect 4649 85298 4683 85332
rect 4649 85230 4683 85264
rect 4649 85162 4683 85196
rect 4649 85094 4683 85128
rect 13677 85366 13711 85400
rect 13677 85298 13711 85332
rect 13677 85230 13711 85264
rect 13677 85162 13711 85196
rect 13677 85094 13711 85128
rect 13763 85366 13797 85400
rect 13763 85298 13797 85332
rect 13763 85230 13797 85264
rect 13763 85162 13797 85196
rect 13763 85094 13797 85128
rect 13849 85366 13883 85400
rect 13849 85298 13883 85332
rect 13849 85230 13883 85264
rect 13849 85162 13883 85196
rect 13849 85094 13883 85128
rect -424 84498 -390 84774
rect -336 84498 -302 84774
rect 4477 75486 4511 75520
rect 4477 75418 4511 75452
rect 4477 75350 4511 75384
rect 4477 75282 4511 75316
rect 4477 75214 4511 75248
rect 4563 75486 4597 75520
rect 4563 75418 4597 75452
rect 4563 75350 4597 75384
rect 4563 75282 4597 75316
rect 4563 75214 4597 75248
rect 4649 75486 4683 75520
rect 4649 75418 4683 75452
rect 4649 75350 4683 75384
rect 4649 75282 4683 75316
rect 4649 75214 4683 75248
rect 13677 75486 13711 75520
rect 13677 75418 13711 75452
rect 13677 75350 13711 75384
rect 13677 75282 13711 75316
rect 13677 75214 13711 75248
rect 13763 75486 13797 75520
rect 13763 75418 13797 75452
rect 13763 75350 13797 75384
rect 13763 75282 13797 75316
rect 13763 75214 13797 75248
rect 13849 75486 13883 75520
rect 13849 75418 13883 75452
rect 13849 75350 13883 75384
rect 13849 75282 13883 75316
rect 13849 75214 13883 75248
rect 22877 75486 22911 75520
rect 22877 75418 22911 75452
rect 22877 75350 22911 75384
rect 22877 75282 22911 75316
rect 22877 75214 22911 75248
rect 22963 75486 22997 75520
rect 22963 75418 22997 75452
rect 22963 75350 22997 75384
rect 22963 75282 22997 75316
rect 22963 75214 22997 75248
rect 23049 75486 23083 75520
rect 23049 75418 23083 75452
rect 23049 75350 23083 75384
rect 23049 75282 23083 75316
rect 23049 75214 23083 75248
rect 32077 75486 32111 75520
rect 32077 75418 32111 75452
rect 32077 75350 32111 75384
rect 32077 75282 32111 75316
rect 32077 75214 32111 75248
rect 32163 75486 32197 75520
rect 32163 75418 32197 75452
rect 32163 75350 32197 75384
rect 32163 75282 32197 75316
rect 32163 75214 32197 75248
rect 32249 75486 32283 75520
rect 32249 75418 32283 75452
rect 32249 75350 32283 75384
rect 32249 75282 32283 75316
rect 32249 75214 32283 75248
rect -424 74618 -390 74894
rect -336 74618 -302 74894
rect 4477 65606 4511 65640
rect 4477 65538 4511 65572
rect 4477 65470 4511 65504
rect 4477 65402 4511 65436
rect 4477 65334 4511 65368
rect 4563 65606 4597 65640
rect 4563 65538 4597 65572
rect 4563 65470 4597 65504
rect 4563 65402 4597 65436
rect 4563 65334 4597 65368
rect 4649 65606 4683 65640
rect 4649 65538 4683 65572
rect 4649 65470 4683 65504
rect 4649 65402 4683 65436
rect 4649 65334 4683 65368
rect 13677 65606 13711 65640
rect 13677 65538 13711 65572
rect 13677 65470 13711 65504
rect 13677 65402 13711 65436
rect 13677 65334 13711 65368
rect 13763 65606 13797 65640
rect 13763 65538 13797 65572
rect 13763 65470 13797 65504
rect 13763 65402 13797 65436
rect 13763 65334 13797 65368
rect 13849 65606 13883 65640
rect 13849 65538 13883 65572
rect 13849 65470 13883 65504
rect 13849 65402 13883 65436
rect 13849 65334 13883 65368
rect 22877 65606 22911 65640
rect 22877 65538 22911 65572
rect 22877 65470 22911 65504
rect 22877 65402 22911 65436
rect 22877 65334 22911 65368
rect 22963 65606 22997 65640
rect 22963 65538 22997 65572
rect 22963 65470 22997 65504
rect 22963 65402 22997 65436
rect 22963 65334 22997 65368
rect 23049 65606 23083 65640
rect 23049 65538 23083 65572
rect 23049 65470 23083 65504
rect 23049 65402 23083 65436
rect 23049 65334 23083 65368
rect 32077 65606 32111 65640
rect 32077 65538 32111 65572
rect 32077 65470 32111 65504
rect 32077 65402 32111 65436
rect 32077 65334 32111 65368
rect 32163 65606 32197 65640
rect 32163 65538 32197 65572
rect 32163 65470 32197 65504
rect 32163 65402 32197 65436
rect 32163 65334 32197 65368
rect 32249 65606 32283 65640
rect 32249 65538 32283 65572
rect 32249 65470 32283 65504
rect 32249 65402 32283 65436
rect 32249 65334 32283 65368
rect 41277 65606 41311 65640
rect 41277 65538 41311 65572
rect 41277 65470 41311 65504
rect 41277 65402 41311 65436
rect 41277 65334 41311 65368
rect 41363 65606 41397 65640
rect 41363 65538 41397 65572
rect 41363 65470 41397 65504
rect 41363 65402 41397 65436
rect 41363 65334 41397 65368
rect 41449 65606 41483 65640
rect 41449 65538 41483 65572
rect 41449 65470 41483 65504
rect 41449 65402 41483 65436
rect 41449 65334 41483 65368
rect 50477 65606 50511 65640
rect 50477 65538 50511 65572
rect 50477 65470 50511 65504
rect 50477 65402 50511 65436
rect 50477 65334 50511 65368
rect 50563 65606 50597 65640
rect 50563 65538 50597 65572
rect 50563 65470 50597 65504
rect 50563 65402 50597 65436
rect 50563 65334 50597 65368
rect 50649 65606 50683 65640
rect 50649 65538 50683 65572
rect 50649 65470 50683 65504
rect 50649 65402 50683 65436
rect 50649 65334 50683 65368
rect 59677 65606 59711 65640
rect 59677 65538 59711 65572
rect 59677 65470 59711 65504
rect 59677 65402 59711 65436
rect 59677 65334 59711 65368
rect 59763 65606 59797 65640
rect 59763 65538 59797 65572
rect 59763 65470 59797 65504
rect 59763 65402 59797 65436
rect 59763 65334 59797 65368
rect 59849 65606 59883 65640
rect 59849 65538 59883 65572
rect 59849 65470 59883 65504
rect 59849 65402 59883 65436
rect 59849 65334 59883 65368
rect 68877 65606 68911 65640
rect 68877 65538 68911 65572
rect 68877 65470 68911 65504
rect 68877 65402 68911 65436
rect 68877 65334 68911 65368
rect 68963 65606 68997 65640
rect 68963 65538 68997 65572
rect 68963 65470 68997 65504
rect 68963 65402 68997 65436
rect 68963 65334 68997 65368
rect 69049 65606 69083 65640
rect 69049 65538 69083 65572
rect 69049 65470 69083 65504
rect 69049 65402 69083 65436
rect 69049 65334 69083 65368
rect -424 64738 -390 65014
rect -336 64738 -302 65014
rect 4477 55726 4511 55760
rect 4477 55658 4511 55692
rect 4477 55590 4511 55624
rect 4477 55522 4511 55556
rect 4477 55454 4511 55488
rect 4563 55726 4597 55760
rect 4563 55658 4597 55692
rect 4563 55590 4597 55624
rect 4563 55522 4597 55556
rect 4563 55454 4597 55488
rect 4649 55726 4683 55760
rect 4649 55658 4683 55692
rect 4649 55590 4683 55624
rect 4649 55522 4683 55556
rect 4649 55454 4683 55488
rect 13677 55726 13711 55760
rect 13677 55658 13711 55692
rect 13677 55590 13711 55624
rect 13677 55522 13711 55556
rect 13677 55454 13711 55488
rect 13763 55726 13797 55760
rect 13763 55658 13797 55692
rect 13763 55590 13797 55624
rect 13763 55522 13797 55556
rect 13763 55454 13797 55488
rect 13849 55726 13883 55760
rect 13849 55658 13883 55692
rect 13849 55590 13883 55624
rect 13849 55522 13883 55556
rect 13849 55454 13883 55488
rect 22877 55726 22911 55760
rect 22877 55658 22911 55692
rect 22877 55590 22911 55624
rect 22877 55522 22911 55556
rect 22877 55454 22911 55488
rect 22963 55726 22997 55760
rect 22963 55658 22997 55692
rect 22963 55590 22997 55624
rect 22963 55522 22997 55556
rect 22963 55454 22997 55488
rect 23049 55726 23083 55760
rect 23049 55658 23083 55692
rect 23049 55590 23083 55624
rect 23049 55522 23083 55556
rect 23049 55454 23083 55488
rect 32077 55726 32111 55760
rect 32077 55658 32111 55692
rect 32077 55590 32111 55624
rect 32077 55522 32111 55556
rect 32077 55454 32111 55488
rect 32163 55726 32197 55760
rect 32163 55658 32197 55692
rect 32163 55590 32197 55624
rect 32163 55522 32197 55556
rect 32163 55454 32197 55488
rect 32249 55726 32283 55760
rect 32249 55658 32283 55692
rect 32249 55590 32283 55624
rect 32249 55522 32283 55556
rect 32249 55454 32283 55488
rect 41277 55726 41311 55760
rect 41277 55658 41311 55692
rect 41277 55590 41311 55624
rect 41277 55522 41311 55556
rect 41277 55454 41311 55488
rect 41363 55726 41397 55760
rect 41363 55658 41397 55692
rect 41363 55590 41397 55624
rect 41363 55522 41397 55556
rect 41363 55454 41397 55488
rect 41449 55726 41483 55760
rect 41449 55658 41483 55692
rect 41449 55590 41483 55624
rect 41449 55522 41483 55556
rect 41449 55454 41483 55488
rect 50477 55726 50511 55760
rect 50477 55658 50511 55692
rect 50477 55590 50511 55624
rect 50477 55522 50511 55556
rect 50477 55454 50511 55488
rect 50563 55726 50597 55760
rect 50563 55658 50597 55692
rect 50563 55590 50597 55624
rect 50563 55522 50597 55556
rect 50563 55454 50597 55488
rect 50649 55726 50683 55760
rect 50649 55658 50683 55692
rect 50649 55590 50683 55624
rect 50649 55522 50683 55556
rect 50649 55454 50683 55488
rect 59677 55726 59711 55760
rect 59677 55658 59711 55692
rect 59677 55590 59711 55624
rect 59677 55522 59711 55556
rect 59677 55454 59711 55488
rect 59763 55726 59797 55760
rect 59763 55658 59797 55692
rect 59763 55590 59797 55624
rect 59763 55522 59797 55556
rect 59763 55454 59797 55488
rect 59849 55726 59883 55760
rect 59849 55658 59883 55692
rect 59849 55590 59883 55624
rect 59849 55522 59883 55556
rect 59849 55454 59883 55488
rect 68877 55726 68911 55760
rect 68877 55658 68911 55692
rect 68877 55590 68911 55624
rect 68877 55522 68911 55556
rect 68877 55454 68911 55488
rect 68963 55726 68997 55760
rect 68963 55658 68997 55692
rect 68963 55590 68997 55624
rect 68963 55522 68997 55556
rect 68963 55454 68997 55488
rect 69049 55726 69083 55760
rect 69049 55658 69083 55692
rect 69049 55590 69083 55624
rect 69049 55522 69083 55556
rect 69049 55454 69083 55488
rect 4477 45846 4511 45880
rect 4477 45778 4511 45812
rect 4477 45710 4511 45744
rect 4477 45642 4511 45676
rect 4477 45574 4511 45608
rect 4563 45846 4597 45880
rect 4563 45778 4597 45812
rect 4563 45710 4597 45744
rect 4563 45642 4597 45676
rect 4563 45574 4597 45608
rect 4649 45846 4683 45880
rect 4649 45778 4683 45812
rect 4649 45710 4683 45744
rect 4649 45642 4683 45676
rect 4649 45574 4683 45608
rect 13677 45846 13711 45880
rect 13677 45778 13711 45812
rect 13677 45710 13711 45744
rect 13677 45642 13711 45676
rect 13677 45574 13711 45608
rect 13763 45846 13797 45880
rect 13763 45778 13797 45812
rect 13763 45710 13797 45744
rect 13763 45642 13797 45676
rect 13763 45574 13797 45608
rect 13849 45846 13883 45880
rect 13849 45778 13883 45812
rect 13849 45710 13883 45744
rect 13849 45642 13883 45676
rect 13849 45574 13883 45608
rect 22877 45846 22911 45880
rect 22877 45778 22911 45812
rect 22877 45710 22911 45744
rect 22877 45642 22911 45676
rect 22877 45574 22911 45608
rect 22963 45846 22997 45880
rect 22963 45778 22997 45812
rect 22963 45710 22997 45744
rect 22963 45642 22997 45676
rect 22963 45574 22997 45608
rect 23049 45846 23083 45880
rect 23049 45778 23083 45812
rect 23049 45710 23083 45744
rect 23049 45642 23083 45676
rect 23049 45574 23083 45608
rect 32077 45846 32111 45880
rect 32077 45778 32111 45812
rect 32077 45710 32111 45744
rect 32077 45642 32111 45676
rect 32077 45574 32111 45608
rect 32163 45846 32197 45880
rect 32163 45778 32197 45812
rect 32163 45710 32197 45744
rect 32163 45642 32197 45676
rect 32163 45574 32197 45608
rect 32249 45846 32283 45880
rect 32249 45778 32283 45812
rect 32249 45710 32283 45744
rect 32249 45642 32283 45676
rect 32249 45574 32283 45608
rect 41277 45846 41311 45880
rect 41277 45778 41311 45812
rect 41277 45710 41311 45744
rect 41277 45642 41311 45676
rect 41277 45574 41311 45608
rect 41363 45846 41397 45880
rect 41363 45778 41397 45812
rect 41363 45710 41397 45744
rect 41363 45642 41397 45676
rect 41363 45574 41397 45608
rect 41449 45846 41483 45880
rect 41449 45778 41483 45812
rect 41449 45710 41483 45744
rect 41449 45642 41483 45676
rect 41449 45574 41483 45608
rect 50477 45846 50511 45880
rect 50477 45778 50511 45812
rect 50477 45710 50511 45744
rect 50477 45642 50511 45676
rect 50477 45574 50511 45608
rect 50563 45846 50597 45880
rect 50563 45778 50597 45812
rect 50563 45710 50597 45744
rect 50563 45642 50597 45676
rect 50563 45574 50597 45608
rect 50649 45846 50683 45880
rect 50649 45778 50683 45812
rect 50649 45710 50683 45744
rect 50649 45642 50683 45676
rect 50649 45574 50683 45608
rect 59677 45846 59711 45880
rect 59677 45778 59711 45812
rect 59677 45710 59711 45744
rect 59677 45642 59711 45676
rect 59677 45574 59711 45608
rect 59763 45846 59797 45880
rect 59763 45778 59797 45812
rect 59763 45710 59797 45744
rect 59763 45642 59797 45676
rect 59763 45574 59797 45608
rect 59849 45846 59883 45880
rect 59849 45778 59883 45812
rect 59849 45710 59883 45744
rect 59849 45642 59883 45676
rect 59849 45574 59883 45608
rect 68877 45846 68911 45880
rect 68877 45778 68911 45812
rect 68877 45710 68911 45744
rect 68877 45642 68911 45676
rect 68877 45574 68911 45608
rect 68963 45846 68997 45880
rect 68963 45778 68997 45812
rect 68963 45710 68997 45744
rect 68963 45642 68997 45676
rect 68963 45574 68997 45608
rect 69049 45846 69083 45880
rect 69049 45778 69083 45812
rect 69049 45710 69083 45744
rect 69049 45642 69083 45676
rect 69049 45574 69083 45608
rect -424 44978 -390 45254
rect -336 44978 -302 45254
rect 4477 35966 4511 36000
rect 4477 35898 4511 35932
rect 4477 35830 4511 35864
rect 4477 35762 4511 35796
rect 4477 35694 4511 35728
rect 4563 35966 4597 36000
rect 4563 35898 4597 35932
rect 4563 35830 4597 35864
rect 4563 35762 4597 35796
rect 4563 35694 4597 35728
rect 4649 35966 4683 36000
rect 4649 35898 4683 35932
rect 4649 35830 4683 35864
rect 4649 35762 4683 35796
rect 4649 35694 4683 35728
rect 13677 35966 13711 36000
rect 13677 35898 13711 35932
rect 13677 35830 13711 35864
rect 13677 35762 13711 35796
rect 13677 35694 13711 35728
rect 13763 35966 13797 36000
rect 13763 35898 13797 35932
rect 13763 35830 13797 35864
rect 13763 35762 13797 35796
rect 13763 35694 13797 35728
rect 13849 35966 13883 36000
rect 13849 35898 13883 35932
rect 13849 35830 13883 35864
rect 13849 35762 13883 35796
rect 13849 35694 13883 35728
rect 22877 35966 22911 36000
rect 22877 35898 22911 35932
rect 22877 35830 22911 35864
rect 22877 35762 22911 35796
rect 22877 35694 22911 35728
rect 22963 35966 22997 36000
rect 22963 35898 22997 35932
rect 22963 35830 22997 35864
rect 22963 35762 22997 35796
rect 22963 35694 22997 35728
rect 23049 35966 23083 36000
rect 23049 35898 23083 35932
rect 23049 35830 23083 35864
rect 23049 35762 23083 35796
rect 23049 35694 23083 35728
rect 32077 35966 32111 36000
rect 32077 35898 32111 35932
rect 32077 35830 32111 35864
rect 32077 35762 32111 35796
rect 32077 35694 32111 35728
rect 32163 35966 32197 36000
rect 32163 35898 32197 35932
rect 32163 35830 32197 35864
rect 32163 35762 32197 35796
rect 32163 35694 32197 35728
rect 32249 35966 32283 36000
rect 32249 35898 32283 35932
rect 32249 35830 32283 35864
rect 32249 35762 32283 35796
rect 32249 35694 32283 35728
rect 41277 35966 41311 36000
rect 41277 35898 41311 35932
rect 41277 35830 41311 35864
rect 41277 35762 41311 35796
rect 41277 35694 41311 35728
rect 41363 35966 41397 36000
rect 41363 35898 41397 35932
rect 41363 35830 41397 35864
rect 41363 35762 41397 35796
rect 41363 35694 41397 35728
rect 41449 35966 41483 36000
rect 41449 35898 41483 35932
rect 41449 35830 41483 35864
rect 41449 35762 41483 35796
rect 41449 35694 41483 35728
rect 50477 35966 50511 36000
rect 50477 35898 50511 35932
rect 50477 35830 50511 35864
rect 50477 35762 50511 35796
rect 50477 35694 50511 35728
rect 50563 35966 50597 36000
rect 50563 35898 50597 35932
rect 50563 35830 50597 35864
rect 50563 35762 50597 35796
rect 50563 35694 50597 35728
rect 50649 35966 50683 36000
rect 50649 35898 50683 35932
rect 50649 35830 50683 35864
rect 50649 35762 50683 35796
rect 50649 35694 50683 35728
rect 59677 35966 59711 36000
rect 59677 35898 59711 35932
rect 59677 35830 59711 35864
rect 59677 35762 59711 35796
rect 59677 35694 59711 35728
rect 59763 35966 59797 36000
rect 59763 35898 59797 35932
rect 59763 35830 59797 35864
rect 59763 35762 59797 35796
rect 59763 35694 59797 35728
rect 59849 35966 59883 36000
rect 59849 35898 59883 35932
rect 59849 35830 59883 35864
rect 59849 35762 59883 35796
rect 59849 35694 59883 35728
rect 68877 35966 68911 36000
rect 68877 35898 68911 35932
rect 68877 35830 68911 35864
rect 68877 35762 68911 35796
rect 68877 35694 68911 35728
rect 68963 35966 68997 36000
rect 68963 35898 68997 35932
rect 68963 35830 68997 35864
rect 68963 35762 68997 35796
rect 68963 35694 68997 35728
rect 69049 35966 69083 36000
rect 69049 35898 69083 35932
rect 69049 35830 69083 35864
rect 69049 35762 69083 35796
rect 69049 35694 69083 35728
rect 4477 26086 4511 26120
rect 4477 26018 4511 26052
rect 4477 25950 4511 25984
rect 4477 25882 4511 25916
rect 4477 25814 4511 25848
rect 4563 26086 4597 26120
rect 4563 26018 4597 26052
rect 4563 25950 4597 25984
rect 4563 25882 4597 25916
rect 4563 25814 4597 25848
rect 4649 26086 4683 26120
rect 4649 26018 4683 26052
rect 4649 25950 4683 25984
rect 4649 25882 4683 25916
rect 4649 25814 4683 25848
rect 13677 26086 13711 26120
rect 13677 26018 13711 26052
rect 13677 25950 13711 25984
rect 13677 25882 13711 25916
rect 13677 25814 13711 25848
rect 13763 26086 13797 26120
rect 13763 26018 13797 26052
rect 13763 25950 13797 25984
rect 13763 25882 13797 25916
rect 13763 25814 13797 25848
rect 13849 26086 13883 26120
rect 13849 26018 13883 26052
rect 13849 25950 13883 25984
rect 13849 25882 13883 25916
rect 13849 25814 13883 25848
rect 22877 26086 22911 26120
rect 22877 26018 22911 26052
rect 22877 25950 22911 25984
rect 22877 25882 22911 25916
rect 22877 25814 22911 25848
rect 22963 26086 22997 26120
rect 22963 26018 22997 26052
rect 22963 25950 22997 25984
rect 22963 25882 22997 25916
rect 22963 25814 22997 25848
rect 23049 26086 23083 26120
rect 23049 26018 23083 26052
rect 23049 25950 23083 25984
rect 23049 25882 23083 25916
rect 23049 25814 23083 25848
rect 32077 26086 32111 26120
rect 32077 26018 32111 26052
rect 32077 25950 32111 25984
rect 32077 25882 32111 25916
rect 32077 25814 32111 25848
rect 32163 26086 32197 26120
rect 32163 26018 32197 26052
rect 32163 25950 32197 25984
rect 32163 25882 32197 25916
rect 32163 25814 32197 25848
rect 32249 26086 32283 26120
rect 32249 26018 32283 26052
rect 32249 25950 32283 25984
rect 32249 25882 32283 25916
rect 32249 25814 32283 25848
rect 41277 26086 41311 26120
rect 41277 26018 41311 26052
rect 41277 25950 41311 25984
rect 41277 25882 41311 25916
rect 41277 25814 41311 25848
rect 41363 26086 41397 26120
rect 41363 26018 41397 26052
rect 41363 25950 41397 25984
rect 41363 25882 41397 25916
rect 41363 25814 41397 25848
rect 41449 26086 41483 26120
rect 41449 26018 41483 26052
rect 41449 25950 41483 25984
rect 41449 25882 41483 25916
rect 41449 25814 41483 25848
rect 50477 26086 50511 26120
rect 50477 26018 50511 26052
rect 50477 25950 50511 25984
rect 50477 25882 50511 25916
rect 50477 25814 50511 25848
rect 50563 26086 50597 26120
rect 50563 26018 50597 26052
rect 50563 25950 50597 25984
rect 50563 25882 50597 25916
rect 50563 25814 50597 25848
rect 50649 26086 50683 26120
rect 50649 26018 50683 26052
rect 50649 25950 50683 25984
rect 50649 25882 50683 25916
rect 50649 25814 50683 25848
rect 59677 26086 59711 26120
rect 59677 26018 59711 26052
rect 59677 25950 59711 25984
rect 59677 25882 59711 25916
rect 59677 25814 59711 25848
rect 59763 26086 59797 26120
rect 59763 26018 59797 26052
rect 59763 25950 59797 25984
rect 59763 25882 59797 25916
rect 59763 25814 59797 25848
rect 59849 26086 59883 26120
rect 59849 26018 59883 26052
rect 59849 25950 59883 25984
rect 59849 25882 59883 25916
rect 59849 25814 59883 25848
rect 68877 26086 68911 26120
rect 68877 26018 68911 26052
rect 68877 25950 68911 25984
rect 68877 25882 68911 25916
rect 68877 25814 68911 25848
rect 68963 26086 68997 26120
rect 68963 26018 68997 26052
rect 68963 25950 68997 25984
rect 68963 25882 68997 25916
rect 68963 25814 68997 25848
rect 69049 26086 69083 26120
rect 69049 26018 69083 26052
rect 69049 25950 69083 25984
rect 69049 25882 69083 25916
rect 69049 25814 69083 25848
rect 4477 16206 4511 16240
rect 4477 16138 4511 16172
rect 4477 16070 4511 16104
rect 4477 16002 4511 16036
rect 4477 15934 4511 15968
rect 4563 16206 4597 16240
rect 4563 16138 4597 16172
rect 4563 16070 4597 16104
rect 4563 16002 4597 16036
rect 4563 15934 4597 15968
rect 4649 16206 4683 16240
rect 4649 16138 4683 16172
rect 4649 16070 4683 16104
rect 4649 16002 4683 16036
rect 4649 15934 4683 15968
rect 13677 16206 13711 16240
rect 13677 16138 13711 16172
rect 13677 16070 13711 16104
rect 13677 16002 13711 16036
rect 13677 15934 13711 15968
rect 13763 16206 13797 16240
rect 13763 16138 13797 16172
rect 13763 16070 13797 16104
rect 13763 16002 13797 16036
rect 13763 15934 13797 15968
rect 13849 16206 13883 16240
rect 13849 16138 13883 16172
rect 13849 16070 13883 16104
rect 13849 16002 13883 16036
rect 13849 15934 13883 15968
rect 22877 16206 22911 16240
rect 22877 16138 22911 16172
rect 22877 16070 22911 16104
rect 22877 16002 22911 16036
rect 22877 15934 22911 15968
rect 22963 16206 22997 16240
rect 22963 16138 22997 16172
rect 22963 16070 22997 16104
rect 22963 16002 22997 16036
rect 22963 15934 22997 15968
rect 23049 16206 23083 16240
rect 23049 16138 23083 16172
rect 23049 16070 23083 16104
rect 23049 16002 23083 16036
rect 23049 15934 23083 15968
rect 32077 16206 32111 16240
rect 32077 16138 32111 16172
rect 32077 16070 32111 16104
rect 32077 16002 32111 16036
rect 32077 15934 32111 15968
rect 32163 16206 32197 16240
rect 32163 16138 32197 16172
rect 32163 16070 32197 16104
rect 32163 16002 32197 16036
rect 32163 15934 32197 15968
rect 32249 16206 32283 16240
rect 32249 16138 32283 16172
rect 32249 16070 32283 16104
rect 32249 16002 32283 16036
rect 32249 15934 32283 15968
rect 41277 16206 41311 16240
rect 41277 16138 41311 16172
rect 41277 16070 41311 16104
rect 41277 16002 41311 16036
rect 41277 15934 41311 15968
rect 41363 16206 41397 16240
rect 41363 16138 41397 16172
rect 41363 16070 41397 16104
rect 41363 16002 41397 16036
rect 41363 15934 41397 15968
rect 41449 16206 41483 16240
rect 41449 16138 41483 16172
rect 41449 16070 41483 16104
rect 41449 16002 41483 16036
rect 41449 15934 41483 15968
rect 50477 16206 50511 16240
rect 50477 16138 50511 16172
rect 50477 16070 50511 16104
rect 50477 16002 50511 16036
rect 50477 15934 50511 15968
rect 50563 16206 50597 16240
rect 50563 16138 50597 16172
rect 50563 16070 50597 16104
rect 50563 16002 50597 16036
rect 50563 15934 50597 15968
rect 50649 16206 50683 16240
rect 50649 16138 50683 16172
rect 50649 16070 50683 16104
rect 50649 16002 50683 16036
rect 50649 15934 50683 15968
rect 59677 16206 59711 16240
rect 59677 16138 59711 16172
rect 59677 16070 59711 16104
rect 59677 16002 59711 16036
rect 59677 15934 59711 15968
rect 59763 16206 59797 16240
rect 59763 16138 59797 16172
rect 59763 16070 59797 16104
rect 59763 16002 59797 16036
rect 59763 15934 59797 15968
rect 59849 16206 59883 16240
rect 59849 16138 59883 16172
rect 59849 16070 59883 16104
rect 59849 16002 59883 16036
rect 59849 15934 59883 15968
rect 68877 16206 68911 16240
rect 68877 16138 68911 16172
rect 68877 16070 68911 16104
rect 68877 16002 68911 16036
rect 68877 15934 68911 15968
rect 68963 16206 68997 16240
rect 68963 16138 68997 16172
rect 68963 16070 68997 16104
rect 68963 16002 68997 16036
rect 68963 15934 68997 15968
rect 69049 16206 69083 16240
rect 69049 16138 69083 16172
rect 69049 16070 69083 16104
rect 69049 16002 69083 16036
rect 69049 15934 69083 15968
rect 4477 6326 4511 6360
rect 4477 6258 4511 6292
rect 4477 6190 4511 6224
rect 4477 6122 4511 6156
rect 4477 6054 4511 6088
rect 4563 6326 4597 6360
rect 4563 6258 4597 6292
rect 4563 6190 4597 6224
rect 4563 6122 4597 6156
rect 4563 6054 4597 6088
rect 4649 6326 4683 6360
rect 4649 6258 4683 6292
rect 4649 6190 4683 6224
rect 4649 6122 4683 6156
rect 4649 6054 4683 6088
rect 13677 6326 13711 6360
rect 13677 6258 13711 6292
rect 13677 6190 13711 6224
rect 13677 6122 13711 6156
rect 13677 6054 13711 6088
rect 13763 6326 13797 6360
rect 13763 6258 13797 6292
rect 13763 6190 13797 6224
rect 13763 6122 13797 6156
rect 13763 6054 13797 6088
rect 13849 6326 13883 6360
rect 13849 6258 13883 6292
rect 13849 6190 13883 6224
rect 13849 6122 13883 6156
rect 13849 6054 13883 6088
rect 22877 6326 22911 6360
rect 22877 6258 22911 6292
rect 22877 6190 22911 6224
rect 22877 6122 22911 6156
rect 22877 6054 22911 6088
rect 22963 6326 22997 6360
rect 22963 6258 22997 6292
rect 22963 6190 22997 6224
rect 22963 6122 22997 6156
rect 22963 6054 22997 6088
rect 23049 6326 23083 6360
rect 23049 6258 23083 6292
rect 23049 6190 23083 6224
rect 23049 6122 23083 6156
rect 23049 6054 23083 6088
rect 32077 6326 32111 6360
rect 32077 6258 32111 6292
rect 32077 6190 32111 6224
rect 32077 6122 32111 6156
rect 32077 6054 32111 6088
rect 32163 6326 32197 6360
rect 32163 6258 32197 6292
rect 32163 6190 32197 6224
rect 32163 6122 32197 6156
rect 32163 6054 32197 6088
rect 32249 6326 32283 6360
rect 32249 6258 32283 6292
rect 32249 6190 32283 6224
rect 32249 6122 32283 6156
rect 32249 6054 32283 6088
rect 41277 6326 41311 6360
rect 41277 6258 41311 6292
rect 41277 6190 41311 6224
rect 41277 6122 41311 6156
rect 41277 6054 41311 6088
rect 41363 6326 41397 6360
rect 41363 6258 41397 6292
rect 41363 6190 41397 6224
rect 41363 6122 41397 6156
rect 41363 6054 41397 6088
rect 41449 6326 41483 6360
rect 41449 6258 41483 6292
rect 41449 6190 41483 6224
rect 41449 6122 41483 6156
rect 41449 6054 41483 6088
rect 50477 6326 50511 6360
rect 50477 6258 50511 6292
rect 50477 6190 50511 6224
rect 50477 6122 50511 6156
rect 50477 6054 50511 6088
rect 50563 6326 50597 6360
rect 50563 6258 50597 6292
rect 50563 6190 50597 6224
rect 50563 6122 50597 6156
rect 50563 6054 50597 6088
rect 50649 6326 50683 6360
rect 50649 6258 50683 6292
rect 50649 6190 50683 6224
rect 50649 6122 50683 6156
rect 50649 6054 50683 6088
rect 59677 6326 59711 6360
rect 59677 6258 59711 6292
rect 59677 6190 59711 6224
rect 59677 6122 59711 6156
rect 59677 6054 59711 6088
rect 59763 6326 59797 6360
rect 59763 6258 59797 6292
rect 59763 6190 59797 6224
rect 59763 6122 59797 6156
rect 59763 6054 59797 6088
rect 59849 6326 59883 6360
rect 59849 6258 59883 6292
rect 59849 6190 59883 6224
rect 59849 6122 59883 6156
rect 59849 6054 59883 6088
rect 68877 6326 68911 6360
rect 68877 6258 68911 6292
rect 68877 6190 68911 6224
rect 68877 6122 68911 6156
rect 68877 6054 68911 6088
rect 68963 6326 68997 6360
rect 68963 6258 68997 6292
rect 68963 6190 68997 6224
rect 68963 6122 68997 6156
rect 68963 6054 68997 6088
rect 69049 6326 69083 6360
rect 69049 6258 69083 6292
rect 69049 6190 69083 6224
rect 69049 6122 69083 6156
rect 69049 6054 69083 6088
rect -424 5458 -390 5734
rect -336 5458 -302 5734
<< pdiffc >>
rect -424 94808 -390 95384
rect -336 94808 -302 95384
rect -424 84928 -390 85504
rect -336 84928 -302 85504
rect -424 75048 -390 75624
rect -336 75048 -302 75624
rect -424 65168 -390 65744
rect -336 65168 -302 65744
rect -424 45408 -390 45984
rect -336 45408 -302 45984
rect -424 5888 -390 6464
rect -336 5888 -302 6464
<< psubdiff >>
rect 4354 95246 4412 95292
rect 4354 95212 4366 95246
rect 4400 95212 4412 95246
rect 4354 95178 4412 95212
rect 4354 95144 4366 95178
rect 4400 95144 4412 95178
rect 4354 95110 4412 95144
rect 4354 95076 4366 95110
rect 4400 95076 4412 95110
rect 4354 95042 4412 95076
rect 4354 95008 4366 95042
rect 4400 95008 4412 95042
rect 4354 94962 4412 95008
rect 4748 95246 4806 95292
rect 4748 95212 4760 95246
rect 4794 95212 4806 95246
rect 4748 95178 4806 95212
rect 4748 95144 4760 95178
rect 4794 95144 4806 95178
rect 4748 95110 4806 95144
rect 4748 95076 4760 95110
rect 4794 95076 4806 95110
rect 4748 95042 4806 95076
rect 4748 95008 4760 95042
rect 4794 95008 4806 95042
rect 4748 94962 4806 95008
rect -458 94276 -260 94278
rect -458 94240 -434 94276
rect -398 94240 -338 94276
rect -300 94240 -260 94276
rect -458 94238 -260 94240
rect 4354 85366 4412 85412
rect 4354 85332 4366 85366
rect 4400 85332 4412 85366
rect 4354 85298 4412 85332
rect 4354 85264 4366 85298
rect 4400 85264 4412 85298
rect 4354 85230 4412 85264
rect 4354 85196 4366 85230
rect 4400 85196 4412 85230
rect 4354 85162 4412 85196
rect 4354 85128 4366 85162
rect 4400 85128 4412 85162
rect 4354 85082 4412 85128
rect 4748 85366 4806 85412
rect 4748 85332 4760 85366
rect 4794 85332 4806 85366
rect 4748 85298 4806 85332
rect 4748 85264 4760 85298
rect 4794 85264 4806 85298
rect 4748 85230 4806 85264
rect 4748 85196 4760 85230
rect 4794 85196 4806 85230
rect 4748 85162 4806 85196
rect 4748 85128 4760 85162
rect 4794 85128 4806 85162
rect 4748 85082 4806 85128
rect 13554 85366 13612 85412
rect 13554 85332 13566 85366
rect 13600 85332 13612 85366
rect 13554 85298 13612 85332
rect 13554 85264 13566 85298
rect 13600 85264 13612 85298
rect 13554 85230 13612 85264
rect 13554 85196 13566 85230
rect 13600 85196 13612 85230
rect 13554 85162 13612 85196
rect 13554 85128 13566 85162
rect 13600 85128 13612 85162
rect 13554 85082 13612 85128
rect 13948 85366 14006 85412
rect 13948 85332 13960 85366
rect 13994 85332 14006 85366
rect 13948 85298 14006 85332
rect 13948 85264 13960 85298
rect 13994 85264 14006 85298
rect 13948 85230 14006 85264
rect 13948 85196 13960 85230
rect 13994 85196 14006 85230
rect 13948 85162 14006 85196
rect 13948 85128 13960 85162
rect 13994 85128 14006 85162
rect 13948 85082 14006 85128
rect -458 84396 -260 84398
rect -458 84360 -434 84396
rect -398 84360 -338 84396
rect -300 84360 -260 84396
rect -458 84358 -260 84360
rect 4354 75486 4412 75532
rect 4354 75452 4366 75486
rect 4400 75452 4412 75486
rect 4354 75418 4412 75452
rect 4354 75384 4366 75418
rect 4400 75384 4412 75418
rect 4354 75350 4412 75384
rect 4354 75316 4366 75350
rect 4400 75316 4412 75350
rect 4354 75282 4412 75316
rect 4354 75248 4366 75282
rect 4400 75248 4412 75282
rect 4354 75202 4412 75248
rect 4748 75486 4806 75532
rect 4748 75452 4760 75486
rect 4794 75452 4806 75486
rect 4748 75418 4806 75452
rect 4748 75384 4760 75418
rect 4794 75384 4806 75418
rect 4748 75350 4806 75384
rect 4748 75316 4760 75350
rect 4794 75316 4806 75350
rect 4748 75282 4806 75316
rect 4748 75248 4760 75282
rect 4794 75248 4806 75282
rect 4748 75202 4806 75248
rect 13554 75486 13612 75532
rect 13554 75452 13566 75486
rect 13600 75452 13612 75486
rect 13554 75418 13612 75452
rect 13554 75384 13566 75418
rect 13600 75384 13612 75418
rect 13554 75350 13612 75384
rect 13554 75316 13566 75350
rect 13600 75316 13612 75350
rect 13554 75282 13612 75316
rect 13554 75248 13566 75282
rect 13600 75248 13612 75282
rect 13554 75202 13612 75248
rect 13948 75486 14006 75532
rect 13948 75452 13960 75486
rect 13994 75452 14006 75486
rect 13948 75418 14006 75452
rect 13948 75384 13960 75418
rect 13994 75384 14006 75418
rect 13948 75350 14006 75384
rect 13948 75316 13960 75350
rect 13994 75316 14006 75350
rect 13948 75282 14006 75316
rect 13948 75248 13960 75282
rect 13994 75248 14006 75282
rect 13948 75202 14006 75248
rect 22754 75486 22812 75532
rect 22754 75452 22766 75486
rect 22800 75452 22812 75486
rect 22754 75418 22812 75452
rect 22754 75384 22766 75418
rect 22800 75384 22812 75418
rect 22754 75350 22812 75384
rect 22754 75316 22766 75350
rect 22800 75316 22812 75350
rect 22754 75282 22812 75316
rect 22754 75248 22766 75282
rect 22800 75248 22812 75282
rect 22754 75202 22812 75248
rect 23148 75486 23206 75532
rect 23148 75452 23160 75486
rect 23194 75452 23206 75486
rect 23148 75418 23206 75452
rect 23148 75384 23160 75418
rect 23194 75384 23206 75418
rect 23148 75350 23206 75384
rect 23148 75316 23160 75350
rect 23194 75316 23206 75350
rect 23148 75282 23206 75316
rect 23148 75248 23160 75282
rect 23194 75248 23206 75282
rect 23148 75202 23206 75248
rect 31954 75486 32012 75532
rect 31954 75452 31966 75486
rect 32000 75452 32012 75486
rect 31954 75418 32012 75452
rect 31954 75384 31966 75418
rect 32000 75384 32012 75418
rect 31954 75350 32012 75384
rect 31954 75316 31966 75350
rect 32000 75316 32012 75350
rect 31954 75282 32012 75316
rect 31954 75248 31966 75282
rect 32000 75248 32012 75282
rect 31954 75202 32012 75248
rect 32348 75486 32406 75532
rect 32348 75452 32360 75486
rect 32394 75452 32406 75486
rect 32348 75418 32406 75452
rect 32348 75384 32360 75418
rect 32394 75384 32406 75418
rect 32348 75350 32406 75384
rect 32348 75316 32360 75350
rect 32394 75316 32406 75350
rect 32348 75282 32406 75316
rect 32348 75248 32360 75282
rect 32394 75248 32406 75282
rect 32348 75202 32406 75248
rect -458 74516 -260 74518
rect -458 74480 -434 74516
rect -398 74480 -338 74516
rect -300 74480 -260 74516
rect -458 74478 -260 74480
rect 4354 65606 4412 65652
rect 4354 65572 4366 65606
rect 4400 65572 4412 65606
rect 4354 65538 4412 65572
rect 4354 65504 4366 65538
rect 4400 65504 4412 65538
rect 4354 65470 4412 65504
rect 4354 65436 4366 65470
rect 4400 65436 4412 65470
rect 4354 65402 4412 65436
rect 4354 65368 4366 65402
rect 4400 65368 4412 65402
rect 4354 65322 4412 65368
rect 4748 65606 4806 65652
rect 4748 65572 4760 65606
rect 4794 65572 4806 65606
rect 4748 65538 4806 65572
rect 4748 65504 4760 65538
rect 4794 65504 4806 65538
rect 4748 65470 4806 65504
rect 4748 65436 4760 65470
rect 4794 65436 4806 65470
rect 4748 65402 4806 65436
rect 4748 65368 4760 65402
rect 4794 65368 4806 65402
rect 4748 65322 4806 65368
rect 13554 65606 13612 65652
rect 13554 65572 13566 65606
rect 13600 65572 13612 65606
rect 13554 65538 13612 65572
rect 13554 65504 13566 65538
rect 13600 65504 13612 65538
rect 13554 65470 13612 65504
rect 13554 65436 13566 65470
rect 13600 65436 13612 65470
rect 13554 65402 13612 65436
rect 13554 65368 13566 65402
rect 13600 65368 13612 65402
rect 13554 65322 13612 65368
rect 13948 65606 14006 65652
rect 13948 65572 13960 65606
rect 13994 65572 14006 65606
rect 13948 65538 14006 65572
rect 13948 65504 13960 65538
rect 13994 65504 14006 65538
rect 13948 65470 14006 65504
rect 13948 65436 13960 65470
rect 13994 65436 14006 65470
rect 13948 65402 14006 65436
rect 13948 65368 13960 65402
rect 13994 65368 14006 65402
rect 13948 65322 14006 65368
rect 22754 65606 22812 65652
rect 22754 65572 22766 65606
rect 22800 65572 22812 65606
rect 22754 65538 22812 65572
rect 22754 65504 22766 65538
rect 22800 65504 22812 65538
rect 22754 65470 22812 65504
rect 22754 65436 22766 65470
rect 22800 65436 22812 65470
rect 22754 65402 22812 65436
rect 22754 65368 22766 65402
rect 22800 65368 22812 65402
rect 22754 65322 22812 65368
rect 23148 65606 23206 65652
rect 23148 65572 23160 65606
rect 23194 65572 23206 65606
rect 23148 65538 23206 65572
rect 23148 65504 23160 65538
rect 23194 65504 23206 65538
rect 23148 65470 23206 65504
rect 23148 65436 23160 65470
rect 23194 65436 23206 65470
rect 23148 65402 23206 65436
rect 23148 65368 23160 65402
rect 23194 65368 23206 65402
rect 23148 65322 23206 65368
rect 31954 65606 32012 65652
rect 31954 65572 31966 65606
rect 32000 65572 32012 65606
rect 31954 65538 32012 65572
rect 31954 65504 31966 65538
rect 32000 65504 32012 65538
rect 31954 65470 32012 65504
rect 31954 65436 31966 65470
rect 32000 65436 32012 65470
rect 31954 65402 32012 65436
rect 31954 65368 31966 65402
rect 32000 65368 32012 65402
rect 31954 65322 32012 65368
rect 32348 65606 32406 65652
rect 32348 65572 32360 65606
rect 32394 65572 32406 65606
rect 32348 65538 32406 65572
rect 32348 65504 32360 65538
rect 32394 65504 32406 65538
rect 32348 65470 32406 65504
rect 32348 65436 32360 65470
rect 32394 65436 32406 65470
rect 32348 65402 32406 65436
rect 32348 65368 32360 65402
rect 32394 65368 32406 65402
rect 32348 65322 32406 65368
rect 41154 65606 41212 65652
rect 41154 65572 41166 65606
rect 41200 65572 41212 65606
rect 41154 65538 41212 65572
rect 41154 65504 41166 65538
rect 41200 65504 41212 65538
rect 41154 65470 41212 65504
rect 41154 65436 41166 65470
rect 41200 65436 41212 65470
rect 41154 65402 41212 65436
rect 41154 65368 41166 65402
rect 41200 65368 41212 65402
rect 41154 65322 41212 65368
rect 41548 65606 41606 65652
rect 41548 65572 41560 65606
rect 41594 65572 41606 65606
rect 41548 65538 41606 65572
rect 41548 65504 41560 65538
rect 41594 65504 41606 65538
rect 41548 65470 41606 65504
rect 41548 65436 41560 65470
rect 41594 65436 41606 65470
rect 41548 65402 41606 65436
rect 41548 65368 41560 65402
rect 41594 65368 41606 65402
rect 41548 65322 41606 65368
rect 50354 65606 50412 65652
rect 50354 65572 50366 65606
rect 50400 65572 50412 65606
rect 50354 65538 50412 65572
rect 50354 65504 50366 65538
rect 50400 65504 50412 65538
rect 50354 65470 50412 65504
rect 50354 65436 50366 65470
rect 50400 65436 50412 65470
rect 50354 65402 50412 65436
rect 50354 65368 50366 65402
rect 50400 65368 50412 65402
rect 50354 65322 50412 65368
rect 50748 65606 50806 65652
rect 50748 65572 50760 65606
rect 50794 65572 50806 65606
rect 50748 65538 50806 65572
rect 50748 65504 50760 65538
rect 50794 65504 50806 65538
rect 50748 65470 50806 65504
rect 50748 65436 50760 65470
rect 50794 65436 50806 65470
rect 50748 65402 50806 65436
rect 50748 65368 50760 65402
rect 50794 65368 50806 65402
rect 50748 65322 50806 65368
rect 59554 65606 59612 65652
rect 59554 65572 59566 65606
rect 59600 65572 59612 65606
rect 59554 65538 59612 65572
rect 59554 65504 59566 65538
rect 59600 65504 59612 65538
rect 59554 65470 59612 65504
rect 59554 65436 59566 65470
rect 59600 65436 59612 65470
rect 59554 65402 59612 65436
rect 59554 65368 59566 65402
rect 59600 65368 59612 65402
rect 59554 65322 59612 65368
rect 59948 65606 60006 65652
rect 59948 65572 59960 65606
rect 59994 65572 60006 65606
rect 59948 65538 60006 65572
rect 59948 65504 59960 65538
rect 59994 65504 60006 65538
rect 59948 65470 60006 65504
rect 59948 65436 59960 65470
rect 59994 65436 60006 65470
rect 59948 65402 60006 65436
rect 59948 65368 59960 65402
rect 59994 65368 60006 65402
rect 59948 65322 60006 65368
rect 68754 65606 68812 65652
rect 68754 65572 68766 65606
rect 68800 65572 68812 65606
rect 68754 65538 68812 65572
rect 68754 65504 68766 65538
rect 68800 65504 68812 65538
rect 68754 65470 68812 65504
rect 68754 65436 68766 65470
rect 68800 65436 68812 65470
rect 68754 65402 68812 65436
rect 68754 65368 68766 65402
rect 68800 65368 68812 65402
rect 68754 65322 68812 65368
rect 69148 65606 69206 65652
rect 69148 65572 69160 65606
rect 69194 65572 69206 65606
rect 69148 65538 69206 65572
rect 69148 65504 69160 65538
rect 69194 65504 69206 65538
rect 69148 65470 69206 65504
rect 69148 65436 69160 65470
rect 69194 65436 69206 65470
rect 69148 65402 69206 65436
rect 69148 65368 69160 65402
rect 69194 65368 69206 65402
rect 69148 65322 69206 65368
rect -458 64636 -260 64638
rect -458 64600 -434 64636
rect -398 64600 -338 64636
rect -300 64600 -260 64636
rect -458 64598 -260 64600
rect 4354 55726 4412 55772
rect 4354 55692 4366 55726
rect 4400 55692 4412 55726
rect 4354 55658 4412 55692
rect 4354 55624 4366 55658
rect 4400 55624 4412 55658
rect 4354 55590 4412 55624
rect 4354 55556 4366 55590
rect 4400 55556 4412 55590
rect 4354 55522 4412 55556
rect 4354 55488 4366 55522
rect 4400 55488 4412 55522
rect 4354 55442 4412 55488
rect 4748 55726 4806 55772
rect 4748 55692 4760 55726
rect 4794 55692 4806 55726
rect 4748 55658 4806 55692
rect 4748 55624 4760 55658
rect 4794 55624 4806 55658
rect 4748 55590 4806 55624
rect 4748 55556 4760 55590
rect 4794 55556 4806 55590
rect 4748 55522 4806 55556
rect 4748 55488 4760 55522
rect 4794 55488 4806 55522
rect 4748 55442 4806 55488
rect 13554 55726 13612 55772
rect 13554 55692 13566 55726
rect 13600 55692 13612 55726
rect 13554 55658 13612 55692
rect 13554 55624 13566 55658
rect 13600 55624 13612 55658
rect 13554 55590 13612 55624
rect 13554 55556 13566 55590
rect 13600 55556 13612 55590
rect 13554 55522 13612 55556
rect 13554 55488 13566 55522
rect 13600 55488 13612 55522
rect 13554 55442 13612 55488
rect 13948 55726 14006 55772
rect 13948 55692 13960 55726
rect 13994 55692 14006 55726
rect 13948 55658 14006 55692
rect 13948 55624 13960 55658
rect 13994 55624 14006 55658
rect 13948 55590 14006 55624
rect 13948 55556 13960 55590
rect 13994 55556 14006 55590
rect 13948 55522 14006 55556
rect 13948 55488 13960 55522
rect 13994 55488 14006 55522
rect 13948 55442 14006 55488
rect 22754 55726 22812 55772
rect 22754 55692 22766 55726
rect 22800 55692 22812 55726
rect 22754 55658 22812 55692
rect 22754 55624 22766 55658
rect 22800 55624 22812 55658
rect 22754 55590 22812 55624
rect 22754 55556 22766 55590
rect 22800 55556 22812 55590
rect 22754 55522 22812 55556
rect 22754 55488 22766 55522
rect 22800 55488 22812 55522
rect 22754 55442 22812 55488
rect 23148 55726 23206 55772
rect 23148 55692 23160 55726
rect 23194 55692 23206 55726
rect 23148 55658 23206 55692
rect 23148 55624 23160 55658
rect 23194 55624 23206 55658
rect 23148 55590 23206 55624
rect 23148 55556 23160 55590
rect 23194 55556 23206 55590
rect 23148 55522 23206 55556
rect 23148 55488 23160 55522
rect 23194 55488 23206 55522
rect 23148 55442 23206 55488
rect 31954 55726 32012 55772
rect 31954 55692 31966 55726
rect 32000 55692 32012 55726
rect 31954 55658 32012 55692
rect 31954 55624 31966 55658
rect 32000 55624 32012 55658
rect 31954 55590 32012 55624
rect 31954 55556 31966 55590
rect 32000 55556 32012 55590
rect 31954 55522 32012 55556
rect 31954 55488 31966 55522
rect 32000 55488 32012 55522
rect 31954 55442 32012 55488
rect 32348 55726 32406 55772
rect 32348 55692 32360 55726
rect 32394 55692 32406 55726
rect 32348 55658 32406 55692
rect 32348 55624 32360 55658
rect 32394 55624 32406 55658
rect 32348 55590 32406 55624
rect 32348 55556 32360 55590
rect 32394 55556 32406 55590
rect 32348 55522 32406 55556
rect 32348 55488 32360 55522
rect 32394 55488 32406 55522
rect 32348 55442 32406 55488
rect 41154 55726 41212 55772
rect 41154 55692 41166 55726
rect 41200 55692 41212 55726
rect 41154 55658 41212 55692
rect 41154 55624 41166 55658
rect 41200 55624 41212 55658
rect 41154 55590 41212 55624
rect 41154 55556 41166 55590
rect 41200 55556 41212 55590
rect 41154 55522 41212 55556
rect 41154 55488 41166 55522
rect 41200 55488 41212 55522
rect 41154 55442 41212 55488
rect 41548 55726 41606 55772
rect 41548 55692 41560 55726
rect 41594 55692 41606 55726
rect 41548 55658 41606 55692
rect 41548 55624 41560 55658
rect 41594 55624 41606 55658
rect 41548 55590 41606 55624
rect 41548 55556 41560 55590
rect 41594 55556 41606 55590
rect 41548 55522 41606 55556
rect 41548 55488 41560 55522
rect 41594 55488 41606 55522
rect 41548 55442 41606 55488
rect 50354 55726 50412 55772
rect 50354 55692 50366 55726
rect 50400 55692 50412 55726
rect 50354 55658 50412 55692
rect 50354 55624 50366 55658
rect 50400 55624 50412 55658
rect 50354 55590 50412 55624
rect 50354 55556 50366 55590
rect 50400 55556 50412 55590
rect 50354 55522 50412 55556
rect 50354 55488 50366 55522
rect 50400 55488 50412 55522
rect 50354 55442 50412 55488
rect 50748 55726 50806 55772
rect 50748 55692 50760 55726
rect 50794 55692 50806 55726
rect 50748 55658 50806 55692
rect 50748 55624 50760 55658
rect 50794 55624 50806 55658
rect 50748 55590 50806 55624
rect 50748 55556 50760 55590
rect 50794 55556 50806 55590
rect 50748 55522 50806 55556
rect 50748 55488 50760 55522
rect 50794 55488 50806 55522
rect 50748 55442 50806 55488
rect 59554 55726 59612 55772
rect 59554 55692 59566 55726
rect 59600 55692 59612 55726
rect 59554 55658 59612 55692
rect 59554 55624 59566 55658
rect 59600 55624 59612 55658
rect 59554 55590 59612 55624
rect 59554 55556 59566 55590
rect 59600 55556 59612 55590
rect 59554 55522 59612 55556
rect 59554 55488 59566 55522
rect 59600 55488 59612 55522
rect 59554 55442 59612 55488
rect 59948 55726 60006 55772
rect 59948 55692 59960 55726
rect 59994 55692 60006 55726
rect 59948 55658 60006 55692
rect 59948 55624 59960 55658
rect 59994 55624 60006 55658
rect 59948 55590 60006 55624
rect 59948 55556 59960 55590
rect 59994 55556 60006 55590
rect 59948 55522 60006 55556
rect 59948 55488 59960 55522
rect 59994 55488 60006 55522
rect 59948 55442 60006 55488
rect 68754 55726 68812 55772
rect 68754 55692 68766 55726
rect 68800 55692 68812 55726
rect 68754 55658 68812 55692
rect 68754 55624 68766 55658
rect 68800 55624 68812 55658
rect 68754 55590 68812 55624
rect 68754 55556 68766 55590
rect 68800 55556 68812 55590
rect 68754 55522 68812 55556
rect 68754 55488 68766 55522
rect 68800 55488 68812 55522
rect 68754 55442 68812 55488
rect 69148 55726 69206 55772
rect 69148 55692 69160 55726
rect 69194 55692 69206 55726
rect 69148 55658 69206 55692
rect 69148 55624 69160 55658
rect 69194 55624 69206 55658
rect 69148 55590 69206 55624
rect 69148 55556 69160 55590
rect 69194 55556 69206 55590
rect 69148 55522 69206 55556
rect 69148 55488 69160 55522
rect 69194 55488 69206 55522
rect 69148 55442 69206 55488
rect 4354 45846 4412 45892
rect 4354 45812 4366 45846
rect 4400 45812 4412 45846
rect 4354 45778 4412 45812
rect 4354 45744 4366 45778
rect 4400 45744 4412 45778
rect 4354 45710 4412 45744
rect 4354 45676 4366 45710
rect 4400 45676 4412 45710
rect 4354 45642 4412 45676
rect 4354 45608 4366 45642
rect 4400 45608 4412 45642
rect 4354 45562 4412 45608
rect 4748 45846 4806 45892
rect 4748 45812 4760 45846
rect 4794 45812 4806 45846
rect 4748 45778 4806 45812
rect 4748 45744 4760 45778
rect 4794 45744 4806 45778
rect 4748 45710 4806 45744
rect 4748 45676 4760 45710
rect 4794 45676 4806 45710
rect 4748 45642 4806 45676
rect 4748 45608 4760 45642
rect 4794 45608 4806 45642
rect 4748 45562 4806 45608
rect 13554 45846 13612 45892
rect 13554 45812 13566 45846
rect 13600 45812 13612 45846
rect 13554 45778 13612 45812
rect 13554 45744 13566 45778
rect 13600 45744 13612 45778
rect 13554 45710 13612 45744
rect 13554 45676 13566 45710
rect 13600 45676 13612 45710
rect 13554 45642 13612 45676
rect 13554 45608 13566 45642
rect 13600 45608 13612 45642
rect 13554 45562 13612 45608
rect 13948 45846 14006 45892
rect 13948 45812 13960 45846
rect 13994 45812 14006 45846
rect 13948 45778 14006 45812
rect 13948 45744 13960 45778
rect 13994 45744 14006 45778
rect 13948 45710 14006 45744
rect 13948 45676 13960 45710
rect 13994 45676 14006 45710
rect 13948 45642 14006 45676
rect 13948 45608 13960 45642
rect 13994 45608 14006 45642
rect 13948 45562 14006 45608
rect 22754 45846 22812 45892
rect 22754 45812 22766 45846
rect 22800 45812 22812 45846
rect 22754 45778 22812 45812
rect 22754 45744 22766 45778
rect 22800 45744 22812 45778
rect 22754 45710 22812 45744
rect 22754 45676 22766 45710
rect 22800 45676 22812 45710
rect 22754 45642 22812 45676
rect 22754 45608 22766 45642
rect 22800 45608 22812 45642
rect 22754 45562 22812 45608
rect 23148 45846 23206 45892
rect 23148 45812 23160 45846
rect 23194 45812 23206 45846
rect 23148 45778 23206 45812
rect 23148 45744 23160 45778
rect 23194 45744 23206 45778
rect 23148 45710 23206 45744
rect 23148 45676 23160 45710
rect 23194 45676 23206 45710
rect 23148 45642 23206 45676
rect 23148 45608 23160 45642
rect 23194 45608 23206 45642
rect 23148 45562 23206 45608
rect 31954 45846 32012 45892
rect 31954 45812 31966 45846
rect 32000 45812 32012 45846
rect 31954 45778 32012 45812
rect 31954 45744 31966 45778
rect 32000 45744 32012 45778
rect 31954 45710 32012 45744
rect 31954 45676 31966 45710
rect 32000 45676 32012 45710
rect 31954 45642 32012 45676
rect 31954 45608 31966 45642
rect 32000 45608 32012 45642
rect 31954 45562 32012 45608
rect 32348 45846 32406 45892
rect 32348 45812 32360 45846
rect 32394 45812 32406 45846
rect 32348 45778 32406 45812
rect 32348 45744 32360 45778
rect 32394 45744 32406 45778
rect 32348 45710 32406 45744
rect 32348 45676 32360 45710
rect 32394 45676 32406 45710
rect 32348 45642 32406 45676
rect 32348 45608 32360 45642
rect 32394 45608 32406 45642
rect 32348 45562 32406 45608
rect 41154 45846 41212 45892
rect 41154 45812 41166 45846
rect 41200 45812 41212 45846
rect 41154 45778 41212 45812
rect 41154 45744 41166 45778
rect 41200 45744 41212 45778
rect 41154 45710 41212 45744
rect 41154 45676 41166 45710
rect 41200 45676 41212 45710
rect 41154 45642 41212 45676
rect 41154 45608 41166 45642
rect 41200 45608 41212 45642
rect 41154 45562 41212 45608
rect 41548 45846 41606 45892
rect 41548 45812 41560 45846
rect 41594 45812 41606 45846
rect 41548 45778 41606 45812
rect 41548 45744 41560 45778
rect 41594 45744 41606 45778
rect 41548 45710 41606 45744
rect 41548 45676 41560 45710
rect 41594 45676 41606 45710
rect 41548 45642 41606 45676
rect 41548 45608 41560 45642
rect 41594 45608 41606 45642
rect 41548 45562 41606 45608
rect 50354 45846 50412 45892
rect 50354 45812 50366 45846
rect 50400 45812 50412 45846
rect 50354 45778 50412 45812
rect 50354 45744 50366 45778
rect 50400 45744 50412 45778
rect 50354 45710 50412 45744
rect 50354 45676 50366 45710
rect 50400 45676 50412 45710
rect 50354 45642 50412 45676
rect 50354 45608 50366 45642
rect 50400 45608 50412 45642
rect 50354 45562 50412 45608
rect 50748 45846 50806 45892
rect 50748 45812 50760 45846
rect 50794 45812 50806 45846
rect 50748 45778 50806 45812
rect 50748 45744 50760 45778
rect 50794 45744 50806 45778
rect 50748 45710 50806 45744
rect 50748 45676 50760 45710
rect 50794 45676 50806 45710
rect 50748 45642 50806 45676
rect 50748 45608 50760 45642
rect 50794 45608 50806 45642
rect 50748 45562 50806 45608
rect 59554 45846 59612 45892
rect 59554 45812 59566 45846
rect 59600 45812 59612 45846
rect 59554 45778 59612 45812
rect 59554 45744 59566 45778
rect 59600 45744 59612 45778
rect 59554 45710 59612 45744
rect 59554 45676 59566 45710
rect 59600 45676 59612 45710
rect 59554 45642 59612 45676
rect 59554 45608 59566 45642
rect 59600 45608 59612 45642
rect 59554 45562 59612 45608
rect 59948 45846 60006 45892
rect 59948 45812 59960 45846
rect 59994 45812 60006 45846
rect 59948 45778 60006 45812
rect 59948 45744 59960 45778
rect 59994 45744 60006 45778
rect 59948 45710 60006 45744
rect 59948 45676 59960 45710
rect 59994 45676 60006 45710
rect 59948 45642 60006 45676
rect 59948 45608 59960 45642
rect 59994 45608 60006 45642
rect 59948 45562 60006 45608
rect 68754 45846 68812 45892
rect 68754 45812 68766 45846
rect 68800 45812 68812 45846
rect 68754 45778 68812 45812
rect 68754 45744 68766 45778
rect 68800 45744 68812 45778
rect 68754 45710 68812 45744
rect 68754 45676 68766 45710
rect 68800 45676 68812 45710
rect 68754 45642 68812 45676
rect 68754 45608 68766 45642
rect 68800 45608 68812 45642
rect 68754 45562 68812 45608
rect 69148 45846 69206 45892
rect 69148 45812 69160 45846
rect 69194 45812 69206 45846
rect 69148 45778 69206 45812
rect 69148 45744 69160 45778
rect 69194 45744 69206 45778
rect 69148 45710 69206 45744
rect 69148 45676 69160 45710
rect 69194 45676 69206 45710
rect 69148 45642 69206 45676
rect 69148 45608 69160 45642
rect 69194 45608 69206 45642
rect 69148 45562 69206 45608
rect -458 44876 -260 44878
rect -458 44840 -434 44876
rect -398 44840 -338 44876
rect -300 44840 -260 44876
rect -458 44838 -260 44840
rect 4354 35966 4412 36012
rect 4354 35932 4366 35966
rect 4400 35932 4412 35966
rect 4354 35898 4412 35932
rect 4354 35864 4366 35898
rect 4400 35864 4412 35898
rect 4354 35830 4412 35864
rect 4354 35796 4366 35830
rect 4400 35796 4412 35830
rect 4354 35762 4412 35796
rect 4354 35728 4366 35762
rect 4400 35728 4412 35762
rect 4354 35682 4412 35728
rect 4748 35966 4806 36012
rect 4748 35932 4760 35966
rect 4794 35932 4806 35966
rect 4748 35898 4806 35932
rect 4748 35864 4760 35898
rect 4794 35864 4806 35898
rect 4748 35830 4806 35864
rect 4748 35796 4760 35830
rect 4794 35796 4806 35830
rect 4748 35762 4806 35796
rect 4748 35728 4760 35762
rect 4794 35728 4806 35762
rect 4748 35682 4806 35728
rect 13554 35966 13612 36012
rect 13554 35932 13566 35966
rect 13600 35932 13612 35966
rect 13554 35898 13612 35932
rect 13554 35864 13566 35898
rect 13600 35864 13612 35898
rect 13554 35830 13612 35864
rect 13554 35796 13566 35830
rect 13600 35796 13612 35830
rect 13554 35762 13612 35796
rect 13554 35728 13566 35762
rect 13600 35728 13612 35762
rect 13554 35682 13612 35728
rect 13948 35966 14006 36012
rect 13948 35932 13960 35966
rect 13994 35932 14006 35966
rect 13948 35898 14006 35932
rect 13948 35864 13960 35898
rect 13994 35864 14006 35898
rect 13948 35830 14006 35864
rect 13948 35796 13960 35830
rect 13994 35796 14006 35830
rect 13948 35762 14006 35796
rect 13948 35728 13960 35762
rect 13994 35728 14006 35762
rect 13948 35682 14006 35728
rect 22754 35966 22812 36012
rect 22754 35932 22766 35966
rect 22800 35932 22812 35966
rect 22754 35898 22812 35932
rect 22754 35864 22766 35898
rect 22800 35864 22812 35898
rect 22754 35830 22812 35864
rect 22754 35796 22766 35830
rect 22800 35796 22812 35830
rect 22754 35762 22812 35796
rect 22754 35728 22766 35762
rect 22800 35728 22812 35762
rect 22754 35682 22812 35728
rect 23148 35966 23206 36012
rect 23148 35932 23160 35966
rect 23194 35932 23206 35966
rect 23148 35898 23206 35932
rect 23148 35864 23160 35898
rect 23194 35864 23206 35898
rect 23148 35830 23206 35864
rect 23148 35796 23160 35830
rect 23194 35796 23206 35830
rect 23148 35762 23206 35796
rect 23148 35728 23160 35762
rect 23194 35728 23206 35762
rect 23148 35682 23206 35728
rect 31954 35966 32012 36012
rect 31954 35932 31966 35966
rect 32000 35932 32012 35966
rect 31954 35898 32012 35932
rect 31954 35864 31966 35898
rect 32000 35864 32012 35898
rect 31954 35830 32012 35864
rect 31954 35796 31966 35830
rect 32000 35796 32012 35830
rect 31954 35762 32012 35796
rect 31954 35728 31966 35762
rect 32000 35728 32012 35762
rect 31954 35682 32012 35728
rect 32348 35966 32406 36012
rect 32348 35932 32360 35966
rect 32394 35932 32406 35966
rect 32348 35898 32406 35932
rect 32348 35864 32360 35898
rect 32394 35864 32406 35898
rect 32348 35830 32406 35864
rect 32348 35796 32360 35830
rect 32394 35796 32406 35830
rect 32348 35762 32406 35796
rect 32348 35728 32360 35762
rect 32394 35728 32406 35762
rect 32348 35682 32406 35728
rect 41154 35966 41212 36012
rect 41154 35932 41166 35966
rect 41200 35932 41212 35966
rect 41154 35898 41212 35932
rect 41154 35864 41166 35898
rect 41200 35864 41212 35898
rect 41154 35830 41212 35864
rect 41154 35796 41166 35830
rect 41200 35796 41212 35830
rect 41154 35762 41212 35796
rect 41154 35728 41166 35762
rect 41200 35728 41212 35762
rect 41154 35682 41212 35728
rect 41548 35966 41606 36012
rect 41548 35932 41560 35966
rect 41594 35932 41606 35966
rect 41548 35898 41606 35932
rect 41548 35864 41560 35898
rect 41594 35864 41606 35898
rect 41548 35830 41606 35864
rect 41548 35796 41560 35830
rect 41594 35796 41606 35830
rect 41548 35762 41606 35796
rect 41548 35728 41560 35762
rect 41594 35728 41606 35762
rect 41548 35682 41606 35728
rect 50354 35966 50412 36012
rect 50354 35932 50366 35966
rect 50400 35932 50412 35966
rect 50354 35898 50412 35932
rect 50354 35864 50366 35898
rect 50400 35864 50412 35898
rect 50354 35830 50412 35864
rect 50354 35796 50366 35830
rect 50400 35796 50412 35830
rect 50354 35762 50412 35796
rect 50354 35728 50366 35762
rect 50400 35728 50412 35762
rect 50354 35682 50412 35728
rect 50748 35966 50806 36012
rect 50748 35932 50760 35966
rect 50794 35932 50806 35966
rect 50748 35898 50806 35932
rect 50748 35864 50760 35898
rect 50794 35864 50806 35898
rect 50748 35830 50806 35864
rect 50748 35796 50760 35830
rect 50794 35796 50806 35830
rect 50748 35762 50806 35796
rect 50748 35728 50760 35762
rect 50794 35728 50806 35762
rect 50748 35682 50806 35728
rect 59554 35966 59612 36012
rect 59554 35932 59566 35966
rect 59600 35932 59612 35966
rect 59554 35898 59612 35932
rect 59554 35864 59566 35898
rect 59600 35864 59612 35898
rect 59554 35830 59612 35864
rect 59554 35796 59566 35830
rect 59600 35796 59612 35830
rect 59554 35762 59612 35796
rect 59554 35728 59566 35762
rect 59600 35728 59612 35762
rect 59554 35682 59612 35728
rect 59948 35966 60006 36012
rect 59948 35932 59960 35966
rect 59994 35932 60006 35966
rect 59948 35898 60006 35932
rect 59948 35864 59960 35898
rect 59994 35864 60006 35898
rect 59948 35830 60006 35864
rect 59948 35796 59960 35830
rect 59994 35796 60006 35830
rect 59948 35762 60006 35796
rect 59948 35728 59960 35762
rect 59994 35728 60006 35762
rect 59948 35682 60006 35728
rect 68754 35966 68812 36012
rect 68754 35932 68766 35966
rect 68800 35932 68812 35966
rect 68754 35898 68812 35932
rect 68754 35864 68766 35898
rect 68800 35864 68812 35898
rect 68754 35830 68812 35864
rect 68754 35796 68766 35830
rect 68800 35796 68812 35830
rect 68754 35762 68812 35796
rect 68754 35728 68766 35762
rect 68800 35728 68812 35762
rect 68754 35682 68812 35728
rect 69148 35966 69206 36012
rect 69148 35932 69160 35966
rect 69194 35932 69206 35966
rect 69148 35898 69206 35932
rect 69148 35864 69160 35898
rect 69194 35864 69206 35898
rect 69148 35830 69206 35864
rect 69148 35796 69160 35830
rect 69194 35796 69206 35830
rect 69148 35762 69206 35796
rect 69148 35728 69160 35762
rect 69194 35728 69206 35762
rect 69148 35682 69206 35728
rect 4354 26086 4412 26132
rect 4354 26052 4366 26086
rect 4400 26052 4412 26086
rect 4354 26018 4412 26052
rect 4354 25984 4366 26018
rect 4400 25984 4412 26018
rect 4354 25950 4412 25984
rect 4354 25916 4366 25950
rect 4400 25916 4412 25950
rect 4354 25882 4412 25916
rect 4354 25848 4366 25882
rect 4400 25848 4412 25882
rect 4354 25802 4412 25848
rect 4748 26086 4806 26132
rect 4748 26052 4760 26086
rect 4794 26052 4806 26086
rect 4748 26018 4806 26052
rect 4748 25984 4760 26018
rect 4794 25984 4806 26018
rect 4748 25950 4806 25984
rect 4748 25916 4760 25950
rect 4794 25916 4806 25950
rect 4748 25882 4806 25916
rect 4748 25848 4760 25882
rect 4794 25848 4806 25882
rect 4748 25802 4806 25848
rect 13554 26086 13612 26132
rect 13554 26052 13566 26086
rect 13600 26052 13612 26086
rect 13554 26018 13612 26052
rect 13554 25984 13566 26018
rect 13600 25984 13612 26018
rect 13554 25950 13612 25984
rect 13554 25916 13566 25950
rect 13600 25916 13612 25950
rect 13554 25882 13612 25916
rect 13554 25848 13566 25882
rect 13600 25848 13612 25882
rect 13554 25802 13612 25848
rect 13948 26086 14006 26132
rect 13948 26052 13960 26086
rect 13994 26052 14006 26086
rect 13948 26018 14006 26052
rect 13948 25984 13960 26018
rect 13994 25984 14006 26018
rect 13948 25950 14006 25984
rect 13948 25916 13960 25950
rect 13994 25916 14006 25950
rect 13948 25882 14006 25916
rect 13948 25848 13960 25882
rect 13994 25848 14006 25882
rect 13948 25802 14006 25848
rect 22754 26086 22812 26132
rect 22754 26052 22766 26086
rect 22800 26052 22812 26086
rect 22754 26018 22812 26052
rect 22754 25984 22766 26018
rect 22800 25984 22812 26018
rect 22754 25950 22812 25984
rect 22754 25916 22766 25950
rect 22800 25916 22812 25950
rect 22754 25882 22812 25916
rect 22754 25848 22766 25882
rect 22800 25848 22812 25882
rect 22754 25802 22812 25848
rect 23148 26086 23206 26132
rect 23148 26052 23160 26086
rect 23194 26052 23206 26086
rect 23148 26018 23206 26052
rect 23148 25984 23160 26018
rect 23194 25984 23206 26018
rect 23148 25950 23206 25984
rect 23148 25916 23160 25950
rect 23194 25916 23206 25950
rect 23148 25882 23206 25916
rect 23148 25848 23160 25882
rect 23194 25848 23206 25882
rect 23148 25802 23206 25848
rect 31954 26086 32012 26132
rect 31954 26052 31966 26086
rect 32000 26052 32012 26086
rect 31954 26018 32012 26052
rect 31954 25984 31966 26018
rect 32000 25984 32012 26018
rect 31954 25950 32012 25984
rect 31954 25916 31966 25950
rect 32000 25916 32012 25950
rect 31954 25882 32012 25916
rect 31954 25848 31966 25882
rect 32000 25848 32012 25882
rect 31954 25802 32012 25848
rect 32348 26086 32406 26132
rect 32348 26052 32360 26086
rect 32394 26052 32406 26086
rect 32348 26018 32406 26052
rect 32348 25984 32360 26018
rect 32394 25984 32406 26018
rect 32348 25950 32406 25984
rect 32348 25916 32360 25950
rect 32394 25916 32406 25950
rect 32348 25882 32406 25916
rect 32348 25848 32360 25882
rect 32394 25848 32406 25882
rect 32348 25802 32406 25848
rect 41154 26086 41212 26132
rect 41154 26052 41166 26086
rect 41200 26052 41212 26086
rect 41154 26018 41212 26052
rect 41154 25984 41166 26018
rect 41200 25984 41212 26018
rect 41154 25950 41212 25984
rect 41154 25916 41166 25950
rect 41200 25916 41212 25950
rect 41154 25882 41212 25916
rect 41154 25848 41166 25882
rect 41200 25848 41212 25882
rect 41154 25802 41212 25848
rect 41548 26086 41606 26132
rect 41548 26052 41560 26086
rect 41594 26052 41606 26086
rect 41548 26018 41606 26052
rect 41548 25984 41560 26018
rect 41594 25984 41606 26018
rect 41548 25950 41606 25984
rect 41548 25916 41560 25950
rect 41594 25916 41606 25950
rect 41548 25882 41606 25916
rect 41548 25848 41560 25882
rect 41594 25848 41606 25882
rect 41548 25802 41606 25848
rect 50354 26086 50412 26132
rect 50354 26052 50366 26086
rect 50400 26052 50412 26086
rect 50354 26018 50412 26052
rect 50354 25984 50366 26018
rect 50400 25984 50412 26018
rect 50354 25950 50412 25984
rect 50354 25916 50366 25950
rect 50400 25916 50412 25950
rect 50354 25882 50412 25916
rect 50354 25848 50366 25882
rect 50400 25848 50412 25882
rect 50354 25802 50412 25848
rect 50748 26086 50806 26132
rect 50748 26052 50760 26086
rect 50794 26052 50806 26086
rect 50748 26018 50806 26052
rect 50748 25984 50760 26018
rect 50794 25984 50806 26018
rect 50748 25950 50806 25984
rect 50748 25916 50760 25950
rect 50794 25916 50806 25950
rect 50748 25882 50806 25916
rect 50748 25848 50760 25882
rect 50794 25848 50806 25882
rect 50748 25802 50806 25848
rect 59554 26086 59612 26132
rect 59554 26052 59566 26086
rect 59600 26052 59612 26086
rect 59554 26018 59612 26052
rect 59554 25984 59566 26018
rect 59600 25984 59612 26018
rect 59554 25950 59612 25984
rect 59554 25916 59566 25950
rect 59600 25916 59612 25950
rect 59554 25882 59612 25916
rect 59554 25848 59566 25882
rect 59600 25848 59612 25882
rect 59554 25802 59612 25848
rect 59948 26086 60006 26132
rect 59948 26052 59960 26086
rect 59994 26052 60006 26086
rect 59948 26018 60006 26052
rect 59948 25984 59960 26018
rect 59994 25984 60006 26018
rect 59948 25950 60006 25984
rect 59948 25916 59960 25950
rect 59994 25916 60006 25950
rect 59948 25882 60006 25916
rect 59948 25848 59960 25882
rect 59994 25848 60006 25882
rect 59948 25802 60006 25848
rect 68754 26086 68812 26132
rect 68754 26052 68766 26086
rect 68800 26052 68812 26086
rect 68754 26018 68812 26052
rect 68754 25984 68766 26018
rect 68800 25984 68812 26018
rect 68754 25950 68812 25984
rect 68754 25916 68766 25950
rect 68800 25916 68812 25950
rect 68754 25882 68812 25916
rect 68754 25848 68766 25882
rect 68800 25848 68812 25882
rect 68754 25802 68812 25848
rect 69148 26086 69206 26132
rect 69148 26052 69160 26086
rect 69194 26052 69206 26086
rect 69148 26018 69206 26052
rect 69148 25984 69160 26018
rect 69194 25984 69206 26018
rect 69148 25950 69206 25984
rect 69148 25916 69160 25950
rect 69194 25916 69206 25950
rect 69148 25882 69206 25916
rect 69148 25848 69160 25882
rect 69194 25848 69206 25882
rect 69148 25802 69206 25848
rect 4354 16206 4412 16252
rect 4354 16172 4366 16206
rect 4400 16172 4412 16206
rect 4354 16138 4412 16172
rect 4354 16104 4366 16138
rect 4400 16104 4412 16138
rect 4354 16070 4412 16104
rect 4354 16036 4366 16070
rect 4400 16036 4412 16070
rect 4354 16002 4412 16036
rect 4354 15968 4366 16002
rect 4400 15968 4412 16002
rect 4354 15922 4412 15968
rect 4748 16206 4806 16252
rect 4748 16172 4760 16206
rect 4794 16172 4806 16206
rect 4748 16138 4806 16172
rect 4748 16104 4760 16138
rect 4794 16104 4806 16138
rect 4748 16070 4806 16104
rect 4748 16036 4760 16070
rect 4794 16036 4806 16070
rect 4748 16002 4806 16036
rect 4748 15968 4760 16002
rect 4794 15968 4806 16002
rect 4748 15922 4806 15968
rect 13554 16206 13612 16252
rect 13554 16172 13566 16206
rect 13600 16172 13612 16206
rect 13554 16138 13612 16172
rect 13554 16104 13566 16138
rect 13600 16104 13612 16138
rect 13554 16070 13612 16104
rect 13554 16036 13566 16070
rect 13600 16036 13612 16070
rect 13554 16002 13612 16036
rect 13554 15968 13566 16002
rect 13600 15968 13612 16002
rect 13554 15922 13612 15968
rect 13948 16206 14006 16252
rect 13948 16172 13960 16206
rect 13994 16172 14006 16206
rect 13948 16138 14006 16172
rect 13948 16104 13960 16138
rect 13994 16104 14006 16138
rect 13948 16070 14006 16104
rect 13948 16036 13960 16070
rect 13994 16036 14006 16070
rect 13948 16002 14006 16036
rect 13948 15968 13960 16002
rect 13994 15968 14006 16002
rect 13948 15922 14006 15968
rect 22754 16206 22812 16252
rect 22754 16172 22766 16206
rect 22800 16172 22812 16206
rect 22754 16138 22812 16172
rect 22754 16104 22766 16138
rect 22800 16104 22812 16138
rect 22754 16070 22812 16104
rect 22754 16036 22766 16070
rect 22800 16036 22812 16070
rect 22754 16002 22812 16036
rect 22754 15968 22766 16002
rect 22800 15968 22812 16002
rect 22754 15922 22812 15968
rect 23148 16206 23206 16252
rect 23148 16172 23160 16206
rect 23194 16172 23206 16206
rect 23148 16138 23206 16172
rect 23148 16104 23160 16138
rect 23194 16104 23206 16138
rect 23148 16070 23206 16104
rect 23148 16036 23160 16070
rect 23194 16036 23206 16070
rect 23148 16002 23206 16036
rect 23148 15968 23160 16002
rect 23194 15968 23206 16002
rect 23148 15922 23206 15968
rect 31954 16206 32012 16252
rect 31954 16172 31966 16206
rect 32000 16172 32012 16206
rect 31954 16138 32012 16172
rect 31954 16104 31966 16138
rect 32000 16104 32012 16138
rect 31954 16070 32012 16104
rect 31954 16036 31966 16070
rect 32000 16036 32012 16070
rect 31954 16002 32012 16036
rect 31954 15968 31966 16002
rect 32000 15968 32012 16002
rect 31954 15922 32012 15968
rect 32348 16206 32406 16252
rect 32348 16172 32360 16206
rect 32394 16172 32406 16206
rect 32348 16138 32406 16172
rect 32348 16104 32360 16138
rect 32394 16104 32406 16138
rect 32348 16070 32406 16104
rect 32348 16036 32360 16070
rect 32394 16036 32406 16070
rect 32348 16002 32406 16036
rect 32348 15968 32360 16002
rect 32394 15968 32406 16002
rect 32348 15922 32406 15968
rect 41154 16206 41212 16252
rect 41154 16172 41166 16206
rect 41200 16172 41212 16206
rect 41154 16138 41212 16172
rect 41154 16104 41166 16138
rect 41200 16104 41212 16138
rect 41154 16070 41212 16104
rect 41154 16036 41166 16070
rect 41200 16036 41212 16070
rect 41154 16002 41212 16036
rect 41154 15968 41166 16002
rect 41200 15968 41212 16002
rect 41154 15922 41212 15968
rect 41548 16206 41606 16252
rect 41548 16172 41560 16206
rect 41594 16172 41606 16206
rect 41548 16138 41606 16172
rect 41548 16104 41560 16138
rect 41594 16104 41606 16138
rect 41548 16070 41606 16104
rect 41548 16036 41560 16070
rect 41594 16036 41606 16070
rect 41548 16002 41606 16036
rect 41548 15968 41560 16002
rect 41594 15968 41606 16002
rect 41548 15922 41606 15968
rect 50354 16206 50412 16252
rect 50354 16172 50366 16206
rect 50400 16172 50412 16206
rect 50354 16138 50412 16172
rect 50354 16104 50366 16138
rect 50400 16104 50412 16138
rect 50354 16070 50412 16104
rect 50354 16036 50366 16070
rect 50400 16036 50412 16070
rect 50354 16002 50412 16036
rect 50354 15968 50366 16002
rect 50400 15968 50412 16002
rect 50354 15922 50412 15968
rect 50748 16206 50806 16252
rect 50748 16172 50760 16206
rect 50794 16172 50806 16206
rect 50748 16138 50806 16172
rect 50748 16104 50760 16138
rect 50794 16104 50806 16138
rect 50748 16070 50806 16104
rect 50748 16036 50760 16070
rect 50794 16036 50806 16070
rect 50748 16002 50806 16036
rect 50748 15968 50760 16002
rect 50794 15968 50806 16002
rect 50748 15922 50806 15968
rect 59554 16206 59612 16252
rect 59554 16172 59566 16206
rect 59600 16172 59612 16206
rect 59554 16138 59612 16172
rect 59554 16104 59566 16138
rect 59600 16104 59612 16138
rect 59554 16070 59612 16104
rect 59554 16036 59566 16070
rect 59600 16036 59612 16070
rect 59554 16002 59612 16036
rect 59554 15968 59566 16002
rect 59600 15968 59612 16002
rect 59554 15922 59612 15968
rect 59948 16206 60006 16252
rect 59948 16172 59960 16206
rect 59994 16172 60006 16206
rect 59948 16138 60006 16172
rect 59948 16104 59960 16138
rect 59994 16104 60006 16138
rect 59948 16070 60006 16104
rect 59948 16036 59960 16070
rect 59994 16036 60006 16070
rect 59948 16002 60006 16036
rect 59948 15968 59960 16002
rect 59994 15968 60006 16002
rect 59948 15922 60006 15968
rect 68754 16206 68812 16252
rect 68754 16172 68766 16206
rect 68800 16172 68812 16206
rect 68754 16138 68812 16172
rect 68754 16104 68766 16138
rect 68800 16104 68812 16138
rect 68754 16070 68812 16104
rect 68754 16036 68766 16070
rect 68800 16036 68812 16070
rect 68754 16002 68812 16036
rect 68754 15968 68766 16002
rect 68800 15968 68812 16002
rect 68754 15922 68812 15968
rect 69148 16206 69206 16252
rect 69148 16172 69160 16206
rect 69194 16172 69206 16206
rect 69148 16138 69206 16172
rect 69148 16104 69160 16138
rect 69194 16104 69206 16138
rect 69148 16070 69206 16104
rect 69148 16036 69160 16070
rect 69194 16036 69206 16070
rect 69148 16002 69206 16036
rect 69148 15968 69160 16002
rect 69194 15968 69206 16002
rect 69148 15922 69206 15968
rect 4354 6326 4412 6372
rect 4354 6292 4366 6326
rect 4400 6292 4412 6326
rect 4354 6258 4412 6292
rect 4354 6224 4366 6258
rect 4400 6224 4412 6258
rect 4354 6190 4412 6224
rect 4354 6156 4366 6190
rect 4400 6156 4412 6190
rect 4354 6122 4412 6156
rect 4354 6088 4366 6122
rect 4400 6088 4412 6122
rect 4354 6042 4412 6088
rect 4748 6326 4806 6372
rect 4748 6292 4760 6326
rect 4794 6292 4806 6326
rect 4748 6258 4806 6292
rect 4748 6224 4760 6258
rect 4794 6224 4806 6258
rect 4748 6190 4806 6224
rect 4748 6156 4760 6190
rect 4794 6156 4806 6190
rect 4748 6122 4806 6156
rect 4748 6088 4760 6122
rect 4794 6088 4806 6122
rect 4748 6042 4806 6088
rect 13554 6326 13612 6372
rect 13554 6292 13566 6326
rect 13600 6292 13612 6326
rect 13554 6258 13612 6292
rect 13554 6224 13566 6258
rect 13600 6224 13612 6258
rect 13554 6190 13612 6224
rect 13554 6156 13566 6190
rect 13600 6156 13612 6190
rect 13554 6122 13612 6156
rect 13554 6088 13566 6122
rect 13600 6088 13612 6122
rect 13554 6042 13612 6088
rect 13948 6326 14006 6372
rect 13948 6292 13960 6326
rect 13994 6292 14006 6326
rect 13948 6258 14006 6292
rect 13948 6224 13960 6258
rect 13994 6224 14006 6258
rect 13948 6190 14006 6224
rect 13948 6156 13960 6190
rect 13994 6156 14006 6190
rect 13948 6122 14006 6156
rect 13948 6088 13960 6122
rect 13994 6088 14006 6122
rect 13948 6042 14006 6088
rect 22754 6326 22812 6372
rect 22754 6292 22766 6326
rect 22800 6292 22812 6326
rect 22754 6258 22812 6292
rect 22754 6224 22766 6258
rect 22800 6224 22812 6258
rect 22754 6190 22812 6224
rect 22754 6156 22766 6190
rect 22800 6156 22812 6190
rect 22754 6122 22812 6156
rect 22754 6088 22766 6122
rect 22800 6088 22812 6122
rect 22754 6042 22812 6088
rect 23148 6326 23206 6372
rect 23148 6292 23160 6326
rect 23194 6292 23206 6326
rect 23148 6258 23206 6292
rect 23148 6224 23160 6258
rect 23194 6224 23206 6258
rect 23148 6190 23206 6224
rect 23148 6156 23160 6190
rect 23194 6156 23206 6190
rect 23148 6122 23206 6156
rect 23148 6088 23160 6122
rect 23194 6088 23206 6122
rect 23148 6042 23206 6088
rect 31954 6326 32012 6372
rect 31954 6292 31966 6326
rect 32000 6292 32012 6326
rect 31954 6258 32012 6292
rect 31954 6224 31966 6258
rect 32000 6224 32012 6258
rect 31954 6190 32012 6224
rect 31954 6156 31966 6190
rect 32000 6156 32012 6190
rect 31954 6122 32012 6156
rect 31954 6088 31966 6122
rect 32000 6088 32012 6122
rect 31954 6042 32012 6088
rect 32348 6326 32406 6372
rect 32348 6292 32360 6326
rect 32394 6292 32406 6326
rect 32348 6258 32406 6292
rect 32348 6224 32360 6258
rect 32394 6224 32406 6258
rect 32348 6190 32406 6224
rect 32348 6156 32360 6190
rect 32394 6156 32406 6190
rect 32348 6122 32406 6156
rect 32348 6088 32360 6122
rect 32394 6088 32406 6122
rect 32348 6042 32406 6088
rect 41154 6326 41212 6372
rect 41154 6292 41166 6326
rect 41200 6292 41212 6326
rect 41154 6258 41212 6292
rect 41154 6224 41166 6258
rect 41200 6224 41212 6258
rect 41154 6190 41212 6224
rect 41154 6156 41166 6190
rect 41200 6156 41212 6190
rect 41154 6122 41212 6156
rect 41154 6088 41166 6122
rect 41200 6088 41212 6122
rect 41154 6042 41212 6088
rect 41548 6326 41606 6372
rect 41548 6292 41560 6326
rect 41594 6292 41606 6326
rect 41548 6258 41606 6292
rect 41548 6224 41560 6258
rect 41594 6224 41606 6258
rect 41548 6190 41606 6224
rect 41548 6156 41560 6190
rect 41594 6156 41606 6190
rect 41548 6122 41606 6156
rect 41548 6088 41560 6122
rect 41594 6088 41606 6122
rect 41548 6042 41606 6088
rect 50354 6326 50412 6372
rect 50354 6292 50366 6326
rect 50400 6292 50412 6326
rect 50354 6258 50412 6292
rect 50354 6224 50366 6258
rect 50400 6224 50412 6258
rect 50354 6190 50412 6224
rect 50354 6156 50366 6190
rect 50400 6156 50412 6190
rect 50354 6122 50412 6156
rect 50354 6088 50366 6122
rect 50400 6088 50412 6122
rect 50354 6042 50412 6088
rect 50748 6326 50806 6372
rect 50748 6292 50760 6326
rect 50794 6292 50806 6326
rect 50748 6258 50806 6292
rect 50748 6224 50760 6258
rect 50794 6224 50806 6258
rect 50748 6190 50806 6224
rect 50748 6156 50760 6190
rect 50794 6156 50806 6190
rect 50748 6122 50806 6156
rect 50748 6088 50760 6122
rect 50794 6088 50806 6122
rect 50748 6042 50806 6088
rect 59554 6326 59612 6372
rect 59554 6292 59566 6326
rect 59600 6292 59612 6326
rect 59554 6258 59612 6292
rect 59554 6224 59566 6258
rect 59600 6224 59612 6258
rect 59554 6190 59612 6224
rect 59554 6156 59566 6190
rect 59600 6156 59612 6190
rect 59554 6122 59612 6156
rect 59554 6088 59566 6122
rect 59600 6088 59612 6122
rect 59554 6042 59612 6088
rect 59948 6326 60006 6372
rect 59948 6292 59960 6326
rect 59994 6292 60006 6326
rect 59948 6258 60006 6292
rect 59948 6224 59960 6258
rect 59994 6224 60006 6258
rect 59948 6190 60006 6224
rect 59948 6156 59960 6190
rect 59994 6156 60006 6190
rect 59948 6122 60006 6156
rect 59948 6088 59960 6122
rect 59994 6088 60006 6122
rect 59948 6042 60006 6088
rect 68754 6326 68812 6372
rect 68754 6292 68766 6326
rect 68800 6292 68812 6326
rect 68754 6258 68812 6292
rect 68754 6224 68766 6258
rect 68800 6224 68812 6258
rect 68754 6190 68812 6224
rect 68754 6156 68766 6190
rect 68800 6156 68812 6190
rect 68754 6122 68812 6156
rect 68754 6088 68766 6122
rect 68800 6088 68812 6122
rect 68754 6042 68812 6088
rect 69148 6326 69206 6372
rect 69148 6292 69160 6326
rect 69194 6292 69206 6326
rect 69148 6258 69206 6292
rect 69148 6224 69160 6258
rect 69194 6224 69206 6258
rect 69148 6190 69206 6224
rect 69148 6156 69160 6190
rect 69194 6156 69206 6190
rect 69148 6122 69206 6156
rect 69148 6088 69160 6122
rect 69194 6088 69206 6122
rect 69148 6042 69206 6088
rect -458 5356 -260 5358
rect -458 5320 -434 5356
rect -398 5320 -338 5356
rect -300 5320 -260 5356
rect -458 5318 -260 5320
<< nsubdiff >>
rect -464 95532 -254 95540
rect -464 95494 -440 95532
rect -392 95494 -326 95532
rect -278 95494 -254 95532
rect -464 95486 -254 95494
rect -464 85652 -254 85660
rect -464 85614 -440 85652
rect -392 85614 -326 85652
rect -278 85614 -254 85652
rect -464 85606 -254 85614
rect -464 75772 -254 75780
rect -464 75734 -440 75772
rect -392 75734 -326 75772
rect -278 75734 -254 75772
rect -464 75726 -254 75734
rect -464 65892 -254 65900
rect -464 65854 -440 65892
rect -392 65854 -326 65892
rect -278 65854 -254 65892
rect -464 65846 -254 65854
rect -464 46132 -254 46140
rect -464 46094 -440 46132
rect -392 46094 -326 46132
rect -278 46094 -254 46132
rect -464 46086 -254 46094
rect -464 6612 -254 6620
rect -464 6574 -440 6612
rect -392 6574 -326 6612
rect -278 6574 -254 6612
rect -464 6566 -254 6574
<< psubdiffcont >>
rect 4366 95212 4400 95246
rect 4366 95144 4400 95178
rect 4366 95076 4400 95110
rect 4366 95008 4400 95042
rect 4760 95212 4794 95246
rect 4760 95144 4794 95178
rect 4760 95076 4794 95110
rect 4760 95008 4794 95042
rect -434 94240 -398 94276
rect -338 94240 -300 94276
rect 4366 85332 4400 85366
rect 4366 85264 4400 85298
rect 4366 85196 4400 85230
rect 4366 85128 4400 85162
rect 4760 85332 4794 85366
rect 4760 85264 4794 85298
rect 4760 85196 4794 85230
rect 4760 85128 4794 85162
rect 13566 85332 13600 85366
rect 13566 85264 13600 85298
rect 13566 85196 13600 85230
rect 13566 85128 13600 85162
rect 13960 85332 13994 85366
rect 13960 85264 13994 85298
rect 13960 85196 13994 85230
rect 13960 85128 13994 85162
rect -434 84360 -398 84396
rect -338 84360 -300 84396
rect 4366 75452 4400 75486
rect 4366 75384 4400 75418
rect 4366 75316 4400 75350
rect 4366 75248 4400 75282
rect 4760 75452 4794 75486
rect 4760 75384 4794 75418
rect 4760 75316 4794 75350
rect 4760 75248 4794 75282
rect 13566 75452 13600 75486
rect 13566 75384 13600 75418
rect 13566 75316 13600 75350
rect 13566 75248 13600 75282
rect 13960 75452 13994 75486
rect 13960 75384 13994 75418
rect 13960 75316 13994 75350
rect 13960 75248 13994 75282
rect 22766 75452 22800 75486
rect 22766 75384 22800 75418
rect 22766 75316 22800 75350
rect 22766 75248 22800 75282
rect 23160 75452 23194 75486
rect 23160 75384 23194 75418
rect 23160 75316 23194 75350
rect 23160 75248 23194 75282
rect 31966 75452 32000 75486
rect 31966 75384 32000 75418
rect 31966 75316 32000 75350
rect 31966 75248 32000 75282
rect 32360 75452 32394 75486
rect 32360 75384 32394 75418
rect 32360 75316 32394 75350
rect 32360 75248 32394 75282
rect -434 74480 -398 74516
rect -338 74480 -300 74516
rect 4366 65572 4400 65606
rect 4366 65504 4400 65538
rect 4366 65436 4400 65470
rect 4366 65368 4400 65402
rect 4760 65572 4794 65606
rect 4760 65504 4794 65538
rect 4760 65436 4794 65470
rect 4760 65368 4794 65402
rect 13566 65572 13600 65606
rect 13566 65504 13600 65538
rect 13566 65436 13600 65470
rect 13566 65368 13600 65402
rect 13960 65572 13994 65606
rect 13960 65504 13994 65538
rect 13960 65436 13994 65470
rect 13960 65368 13994 65402
rect 22766 65572 22800 65606
rect 22766 65504 22800 65538
rect 22766 65436 22800 65470
rect 22766 65368 22800 65402
rect 23160 65572 23194 65606
rect 23160 65504 23194 65538
rect 23160 65436 23194 65470
rect 23160 65368 23194 65402
rect 31966 65572 32000 65606
rect 31966 65504 32000 65538
rect 31966 65436 32000 65470
rect 31966 65368 32000 65402
rect 32360 65572 32394 65606
rect 32360 65504 32394 65538
rect 32360 65436 32394 65470
rect 32360 65368 32394 65402
rect 41166 65572 41200 65606
rect 41166 65504 41200 65538
rect 41166 65436 41200 65470
rect 41166 65368 41200 65402
rect 41560 65572 41594 65606
rect 41560 65504 41594 65538
rect 41560 65436 41594 65470
rect 41560 65368 41594 65402
rect 50366 65572 50400 65606
rect 50366 65504 50400 65538
rect 50366 65436 50400 65470
rect 50366 65368 50400 65402
rect 50760 65572 50794 65606
rect 50760 65504 50794 65538
rect 50760 65436 50794 65470
rect 50760 65368 50794 65402
rect 59566 65572 59600 65606
rect 59566 65504 59600 65538
rect 59566 65436 59600 65470
rect 59566 65368 59600 65402
rect 59960 65572 59994 65606
rect 59960 65504 59994 65538
rect 59960 65436 59994 65470
rect 59960 65368 59994 65402
rect 68766 65572 68800 65606
rect 68766 65504 68800 65538
rect 68766 65436 68800 65470
rect 68766 65368 68800 65402
rect 69160 65572 69194 65606
rect 69160 65504 69194 65538
rect 69160 65436 69194 65470
rect 69160 65368 69194 65402
rect -434 64600 -398 64636
rect -338 64600 -300 64636
rect 4366 55692 4400 55726
rect 4366 55624 4400 55658
rect 4366 55556 4400 55590
rect 4366 55488 4400 55522
rect 4760 55692 4794 55726
rect 4760 55624 4794 55658
rect 4760 55556 4794 55590
rect 4760 55488 4794 55522
rect 13566 55692 13600 55726
rect 13566 55624 13600 55658
rect 13566 55556 13600 55590
rect 13566 55488 13600 55522
rect 13960 55692 13994 55726
rect 13960 55624 13994 55658
rect 13960 55556 13994 55590
rect 13960 55488 13994 55522
rect 22766 55692 22800 55726
rect 22766 55624 22800 55658
rect 22766 55556 22800 55590
rect 22766 55488 22800 55522
rect 23160 55692 23194 55726
rect 23160 55624 23194 55658
rect 23160 55556 23194 55590
rect 23160 55488 23194 55522
rect 31966 55692 32000 55726
rect 31966 55624 32000 55658
rect 31966 55556 32000 55590
rect 31966 55488 32000 55522
rect 32360 55692 32394 55726
rect 32360 55624 32394 55658
rect 32360 55556 32394 55590
rect 32360 55488 32394 55522
rect 41166 55692 41200 55726
rect 41166 55624 41200 55658
rect 41166 55556 41200 55590
rect 41166 55488 41200 55522
rect 41560 55692 41594 55726
rect 41560 55624 41594 55658
rect 41560 55556 41594 55590
rect 41560 55488 41594 55522
rect 50366 55692 50400 55726
rect 50366 55624 50400 55658
rect 50366 55556 50400 55590
rect 50366 55488 50400 55522
rect 50760 55692 50794 55726
rect 50760 55624 50794 55658
rect 50760 55556 50794 55590
rect 50760 55488 50794 55522
rect 59566 55692 59600 55726
rect 59566 55624 59600 55658
rect 59566 55556 59600 55590
rect 59566 55488 59600 55522
rect 59960 55692 59994 55726
rect 59960 55624 59994 55658
rect 59960 55556 59994 55590
rect 59960 55488 59994 55522
rect 68766 55692 68800 55726
rect 68766 55624 68800 55658
rect 68766 55556 68800 55590
rect 68766 55488 68800 55522
rect 69160 55692 69194 55726
rect 69160 55624 69194 55658
rect 69160 55556 69194 55590
rect 69160 55488 69194 55522
rect 4366 45812 4400 45846
rect 4366 45744 4400 45778
rect 4366 45676 4400 45710
rect 4366 45608 4400 45642
rect 4760 45812 4794 45846
rect 4760 45744 4794 45778
rect 4760 45676 4794 45710
rect 4760 45608 4794 45642
rect 13566 45812 13600 45846
rect 13566 45744 13600 45778
rect 13566 45676 13600 45710
rect 13566 45608 13600 45642
rect 13960 45812 13994 45846
rect 13960 45744 13994 45778
rect 13960 45676 13994 45710
rect 13960 45608 13994 45642
rect 22766 45812 22800 45846
rect 22766 45744 22800 45778
rect 22766 45676 22800 45710
rect 22766 45608 22800 45642
rect 23160 45812 23194 45846
rect 23160 45744 23194 45778
rect 23160 45676 23194 45710
rect 23160 45608 23194 45642
rect 31966 45812 32000 45846
rect 31966 45744 32000 45778
rect 31966 45676 32000 45710
rect 31966 45608 32000 45642
rect 32360 45812 32394 45846
rect 32360 45744 32394 45778
rect 32360 45676 32394 45710
rect 32360 45608 32394 45642
rect 41166 45812 41200 45846
rect 41166 45744 41200 45778
rect 41166 45676 41200 45710
rect 41166 45608 41200 45642
rect 41560 45812 41594 45846
rect 41560 45744 41594 45778
rect 41560 45676 41594 45710
rect 41560 45608 41594 45642
rect 50366 45812 50400 45846
rect 50366 45744 50400 45778
rect 50366 45676 50400 45710
rect 50366 45608 50400 45642
rect 50760 45812 50794 45846
rect 50760 45744 50794 45778
rect 50760 45676 50794 45710
rect 50760 45608 50794 45642
rect 59566 45812 59600 45846
rect 59566 45744 59600 45778
rect 59566 45676 59600 45710
rect 59566 45608 59600 45642
rect 59960 45812 59994 45846
rect 59960 45744 59994 45778
rect 59960 45676 59994 45710
rect 59960 45608 59994 45642
rect 68766 45812 68800 45846
rect 68766 45744 68800 45778
rect 68766 45676 68800 45710
rect 68766 45608 68800 45642
rect 69160 45812 69194 45846
rect 69160 45744 69194 45778
rect 69160 45676 69194 45710
rect 69160 45608 69194 45642
rect -434 44840 -398 44876
rect -338 44840 -300 44876
rect 4366 35932 4400 35966
rect 4366 35864 4400 35898
rect 4366 35796 4400 35830
rect 4366 35728 4400 35762
rect 4760 35932 4794 35966
rect 4760 35864 4794 35898
rect 4760 35796 4794 35830
rect 4760 35728 4794 35762
rect 13566 35932 13600 35966
rect 13566 35864 13600 35898
rect 13566 35796 13600 35830
rect 13566 35728 13600 35762
rect 13960 35932 13994 35966
rect 13960 35864 13994 35898
rect 13960 35796 13994 35830
rect 13960 35728 13994 35762
rect 22766 35932 22800 35966
rect 22766 35864 22800 35898
rect 22766 35796 22800 35830
rect 22766 35728 22800 35762
rect 23160 35932 23194 35966
rect 23160 35864 23194 35898
rect 23160 35796 23194 35830
rect 23160 35728 23194 35762
rect 31966 35932 32000 35966
rect 31966 35864 32000 35898
rect 31966 35796 32000 35830
rect 31966 35728 32000 35762
rect 32360 35932 32394 35966
rect 32360 35864 32394 35898
rect 32360 35796 32394 35830
rect 32360 35728 32394 35762
rect 41166 35932 41200 35966
rect 41166 35864 41200 35898
rect 41166 35796 41200 35830
rect 41166 35728 41200 35762
rect 41560 35932 41594 35966
rect 41560 35864 41594 35898
rect 41560 35796 41594 35830
rect 41560 35728 41594 35762
rect 50366 35932 50400 35966
rect 50366 35864 50400 35898
rect 50366 35796 50400 35830
rect 50366 35728 50400 35762
rect 50760 35932 50794 35966
rect 50760 35864 50794 35898
rect 50760 35796 50794 35830
rect 50760 35728 50794 35762
rect 59566 35932 59600 35966
rect 59566 35864 59600 35898
rect 59566 35796 59600 35830
rect 59566 35728 59600 35762
rect 59960 35932 59994 35966
rect 59960 35864 59994 35898
rect 59960 35796 59994 35830
rect 59960 35728 59994 35762
rect 68766 35932 68800 35966
rect 68766 35864 68800 35898
rect 68766 35796 68800 35830
rect 68766 35728 68800 35762
rect 69160 35932 69194 35966
rect 69160 35864 69194 35898
rect 69160 35796 69194 35830
rect 69160 35728 69194 35762
rect 4366 26052 4400 26086
rect 4366 25984 4400 26018
rect 4366 25916 4400 25950
rect 4366 25848 4400 25882
rect 4760 26052 4794 26086
rect 4760 25984 4794 26018
rect 4760 25916 4794 25950
rect 4760 25848 4794 25882
rect 13566 26052 13600 26086
rect 13566 25984 13600 26018
rect 13566 25916 13600 25950
rect 13566 25848 13600 25882
rect 13960 26052 13994 26086
rect 13960 25984 13994 26018
rect 13960 25916 13994 25950
rect 13960 25848 13994 25882
rect 22766 26052 22800 26086
rect 22766 25984 22800 26018
rect 22766 25916 22800 25950
rect 22766 25848 22800 25882
rect 23160 26052 23194 26086
rect 23160 25984 23194 26018
rect 23160 25916 23194 25950
rect 23160 25848 23194 25882
rect 31966 26052 32000 26086
rect 31966 25984 32000 26018
rect 31966 25916 32000 25950
rect 31966 25848 32000 25882
rect 32360 26052 32394 26086
rect 32360 25984 32394 26018
rect 32360 25916 32394 25950
rect 32360 25848 32394 25882
rect 41166 26052 41200 26086
rect 41166 25984 41200 26018
rect 41166 25916 41200 25950
rect 41166 25848 41200 25882
rect 41560 26052 41594 26086
rect 41560 25984 41594 26018
rect 41560 25916 41594 25950
rect 41560 25848 41594 25882
rect 50366 26052 50400 26086
rect 50366 25984 50400 26018
rect 50366 25916 50400 25950
rect 50366 25848 50400 25882
rect 50760 26052 50794 26086
rect 50760 25984 50794 26018
rect 50760 25916 50794 25950
rect 50760 25848 50794 25882
rect 59566 26052 59600 26086
rect 59566 25984 59600 26018
rect 59566 25916 59600 25950
rect 59566 25848 59600 25882
rect 59960 26052 59994 26086
rect 59960 25984 59994 26018
rect 59960 25916 59994 25950
rect 59960 25848 59994 25882
rect 68766 26052 68800 26086
rect 68766 25984 68800 26018
rect 68766 25916 68800 25950
rect 68766 25848 68800 25882
rect 69160 26052 69194 26086
rect 69160 25984 69194 26018
rect 69160 25916 69194 25950
rect 69160 25848 69194 25882
rect 4366 16172 4400 16206
rect 4366 16104 4400 16138
rect 4366 16036 4400 16070
rect 4366 15968 4400 16002
rect 4760 16172 4794 16206
rect 4760 16104 4794 16138
rect 4760 16036 4794 16070
rect 4760 15968 4794 16002
rect 13566 16172 13600 16206
rect 13566 16104 13600 16138
rect 13566 16036 13600 16070
rect 13566 15968 13600 16002
rect 13960 16172 13994 16206
rect 13960 16104 13994 16138
rect 13960 16036 13994 16070
rect 13960 15968 13994 16002
rect 22766 16172 22800 16206
rect 22766 16104 22800 16138
rect 22766 16036 22800 16070
rect 22766 15968 22800 16002
rect 23160 16172 23194 16206
rect 23160 16104 23194 16138
rect 23160 16036 23194 16070
rect 23160 15968 23194 16002
rect 31966 16172 32000 16206
rect 31966 16104 32000 16138
rect 31966 16036 32000 16070
rect 31966 15968 32000 16002
rect 32360 16172 32394 16206
rect 32360 16104 32394 16138
rect 32360 16036 32394 16070
rect 32360 15968 32394 16002
rect 41166 16172 41200 16206
rect 41166 16104 41200 16138
rect 41166 16036 41200 16070
rect 41166 15968 41200 16002
rect 41560 16172 41594 16206
rect 41560 16104 41594 16138
rect 41560 16036 41594 16070
rect 41560 15968 41594 16002
rect 50366 16172 50400 16206
rect 50366 16104 50400 16138
rect 50366 16036 50400 16070
rect 50366 15968 50400 16002
rect 50760 16172 50794 16206
rect 50760 16104 50794 16138
rect 50760 16036 50794 16070
rect 50760 15968 50794 16002
rect 59566 16172 59600 16206
rect 59566 16104 59600 16138
rect 59566 16036 59600 16070
rect 59566 15968 59600 16002
rect 59960 16172 59994 16206
rect 59960 16104 59994 16138
rect 59960 16036 59994 16070
rect 59960 15968 59994 16002
rect 68766 16172 68800 16206
rect 68766 16104 68800 16138
rect 68766 16036 68800 16070
rect 68766 15968 68800 16002
rect 69160 16172 69194 16206
rect 69160 16104 69194 16138
rect 69160 16036 69194 16070
rect 69160 15968 69194 16002
rect 4366 6292 4400 6326
rect 4366 6224 4400 6258
rect 4366 6156 4400 6190
rect 4366 6088 4400 6122
rect 4760 6292 4794 6326
rect 4760 6224 4794 6258
rect 4760 6156 4794 6190
rect 4760 6088 4794 6122
rect 13566 6292 13600 6326
rect 13566 6224 13600 6258
rect 13566 6156 13600 6190
rect 13566 6088 13600 6122
rect 13960 6292 13994 6326
rect 13960 6224 13994 6258
rect 13960 6156 13994 6190
rect 13960 6088 13994 6122
rect 22766 6292 22800 6326
rect 22766 6224 22800 6258
rect 22766 6156 22800 6190
rect 22766 6088 22800 6122
rect 23160 6292 23194 6326
rect 23160 6224 23194 6258
rect 23160 6156 23194 6190
rect 23160 6088 23194 6122
rect 31966 6292 32000 6326
rect 31966 6224 32000 6258
rect 31966 6156 32000 6190
rect 31966 6088 32000 6122
rect 32360 6292 32394 6326
rect 32360 6224 32394 6258
rect 32360 6156 32394 6190
rect 32360 6088 32394 6122
rect 41166 6292 41200 6326
rect 41166 6224 41200 6258
rect 41166 6156 41200 6190
rect 41166 6088 41200 6122
rect 41560 6292 41594 6326
rect 41560 6224 41594 6258
rect 41560 6156 41594 6190
rect 41560 6088 41594 6122
rect 50366 6292 50400 6326
rect 50366 6224 50400 6258
rect 50366 6156 50400 6190
rect 50366 6088 50400 6122
rect 50760 6292 50794 6326
rect 50760 6224 50794 6258
rect 50760 6156 50794 6190
rect 50760 6088 50794 6122
rect 59566 6292 59600 6326
rect 59566 6224 59600 6258
rect 59566 6156 59600 6190
rect 59566 6088 59600 6122
rect 59960 6292 59994 6326
rect 59960 6224 59994 6258
rect 59960 6156 59994 6190
rect 59960 6088 59994 6122
rect 68766 6292 68800 6326
rect 68766 6224 68800 6258
rect 68766 6156 68800 6190
rect 68766 6088 68800 6122
rect 69160 6292 69194 6326
rect 69160 6224 69194 6258
rect 69160 6156 69194 6190
rect 69160 6088 69194 6122
rect -434 5320 -398 5356
rect -338 5320 -300 5356
<< nsubdiffcont >>
rect -440 95494 -392 95532
rect -326 95494 -278 95532
rect -440 85614 -392 85652
rect -326 85614 -278 85652
rect -440 75734 -392 75772
rect -326 75734 -278 75772
rect -440 65854 -392 65892
rect -326 65854 -278 65892
rect -440 46094 -392 46132
rect -326 46094 -278 46132
rect -440 6574 -392 6612
rect -326 6574 -278 6612
<< poly >>
rect -378 95396 -348 95422
rect 4479 95364 4681 95384
rect 4479 95330 4495 95364
rect 4529 95330 4563 95364
rect 4597 95330 4631 95364
rect 4665 95330 4681 95364
rect 4479 95314 4681 95330
rect 4522 95292 4552 95314
rect 4608 95292 4638 95314
rect 4522 94940 4552 94962
rect 4608 94940 4638 94962
rect 4479 94924 4681 94940
rect 4479 94890 4495 94924
rect 4529 94890 4563 94924
rect 4597 94890 4631 94924
rect 4665 94890 4681 94924
rect 4479 94870 4681 94890
rect -378 94752 -348 94796
rect -240 94752 -160 94760
rect -378 94740 -160 94752
rect -378 94700 -220 94740
rect -180 94700 -160 94740
rect -378 94690 -160 94700
rect -378 94666 -348 94690
rect -240 94680 -160 94690
rect -378 94340 -348 94366
rect -378 85516 -348 85542
rect 4479 85484 4681 85504
rect 4479 85450 4495 85484
rect 4529 85450 4563 85484
rect 4597 85450 4631 85484
rect 4665 85450 4681 85484
rect 4479 85434 4681 85450
rect 4522 85412 4552 85434
rect 4608 85412 4638 85434
rect 4522 85060 4552 85082
rect 4608 85060 4638 85082
rect 4479 85044 4681 85060
rect 4479 85010 4495 85044
rect 4529 85010 4563 85044
rect 4597 85010 4631 85044
rect 4665 85010 4681 85044
rect 4479 84990 4681 85010
rect 13679 85484 13881 85504
rect 13679 85450 13695 85484
rect 13729 85450 13763 85484
rect 13797 85450 13831 85484
rect 13865 85450 13881 85484
rect 13679 85434 13881 85450
rect 13722 85412 13752 85434
rect 13808 85412 13838 85434
rect 13722 85060 13752 85082
rect 13808 85060 13838 85082
rect 13679 85044 13881 85060
rect 13679 85010 13695 85044
rect 13729 85010 13763 85044
rect 13797 85010 13831 85044
rect 13865 85010 13881 85044
rect 13679 84990 13881 85010
rect -378 84872 -348 84916
rect -240 84872 -160 84880
rect -378 84860 -160 84872
rect -378 84820 -220 84860
rect -180 84820 -160 84860
rect -378 84810 -160 84820
rect -378 84786 -348 84810
rect -240 84800 -160 84810
rect -378 84460 -348 84486
rect -378 75636 -348 75662
rect 4479 75604 4681 75624
rect 4479 75570 4495 75604
rect 4529 75570 4563 75604
rect 4597 75570 4631 75604
rect 4665 75570 4681 75604
rect 4479 75554 4681 75570
rect 4522 75532 4552 75554
rect 4608 75532 4638 75554
rect 4522 75180 4552 75202
rect 4608 75180 4638 75202
rect 4479 75164 4681 75180
rect 4479 75130 4495 75164
rect 4529 75130 4563 75164
rect 4597 75130 4631 75164
rect 4665 75130 4681 75164
rect 4479 75110 4681 75130
rect 13679 75604 13881 75624
rect 13679 75570 13695 75604
rect 13729 75570 13763 75604
rect 13797 75570 13831 75604
rect 13865 75570 13881 75604
rect 13679 75554 13881 75570
rect 13722 75532 13752 75554
rect 13808 75532 13838 75554
rect 13722 75180 13752 75202
rect 13808 75180 13838 75202
rect 13679 75164 13881 75180
rect 13679 75130 13695 75164
rect 13729 75130 13763 75164
rect 13797 75130 13831 75164
rect 13865 75130 13881 75164
rect 13679 75110 13881 75130
rect 22879 75604 23081 75624
rect 22879 75570 22895 75604
rect 22929 75570 22963 75604
rect 22997 75570 23031 75604
rect 23065 75570 23081 75604
rect 22879 75554 23081 75570
rect 22922 75532 22952 75554
rect 23008 75532 23038 75554
rect 22922 75180 22952 75202
rect 23008 75180 23038 75202
rect 22879 75164 23081 75180
rect 22879 75130 22895 75164
rect 22929 75130 22963 75164
rect 22997 75130 23031 75164
rect 23065 75130 23081 75164
rect 22879 75110 23081 75130
rect 32079 75604 32281 75624
rect 32079 75570 32095 75604
rect 32129 75570 32163 75604
rect 32197 75570 32231 75604
rect 32265 75570 32281 75604
rect 32079 75554 32281 75570
rect 32122 75532 32152 75554
rect 32208 75532 32238 75554
rect 32122 75180 32152 75202
rect 32208 75180 32238 75202
rect 32079 75164 32281 75180
rect 32079 75130 32095 75164
rect 32129 75130 32163 75164
rect 32197 75130 32231 75164
rect 32265 75130 32281 75164
rect 32079 75110 32281 75130
rect -378 74992 -348 75036
rect -240 74992 -160 75000
rect -378 74980 -160 74992
rect -378 74940 -220 74980
rect -180 74940 -160 74980
rect -378 74930 -160 74940
rect -378 74906 -348 74930
rect -240 74920 -160 74930
rect -378 74580 -348 74606
rect -378 65756 -348 65782
rect 4479 65724 4681 65744
rect 4479 65690 4495 65724
rect 4529 65690 4563 65724
rect 4597 65690 4631 65724
rect 4665 65690 4681 65724
rect 4479 65674 4681 65690
rect 4522 65652 4552 65674
rect 4608 65652 4638 65674
rect 4522 65300 4552 65322
rect 4608 65300 4638 65322
rect 4479 65284 4681 65300
rect 4479 65250 4495 65284
rect 4529 65250 4563 65284
rect 4597 65250 4631 65284
rect 4665 65250 4681 65284
rect 4479 65230 4681 65250
rect 13679 65724 13881 65744
rect 13679 65690 13695 65724
rect 13729 65690 13763 65724
rect 13797 65690 13831 65724
rect 13865 65690 13881 65724
rect 13679 65674 13881 65690
rect 13722 65652 13752 65674
rect 13808 65652 13838 65674
rect 13722 65300 13752 65322
rect 13808 65300 13838 65322
rect 13679 65284 13881 65300
rect 13679 65250 13695 65284
rect 13729 65250 13763 65284
rect 13797 65250 13831 65284
rect 13865 65250 13881 65284
rect 13679 65230 13881 65250
rect 22879 65724 23081 65744
rect 22879 65690 22895 65724
rect 22929 65690 22963 65724
rect 22997 65690 23031 65724
rect 23065 65690 23081 65724
rect 22879 65674 23081 65690
rect 22922 65652 22952 65674
rect 23008 65652 23038 65674
rect 22922 65300 22952 65322
rect 23008 65300 23038 65322
rect 22879 65284 23081 65300
rect 22879 65250 22895 65284
rect 22929 65250 22963 65284
rect 22997 65250 23031 65284
rect 23065 65250 23081 65284
rect 22879 65230 23081 65250
rect 32079 65724 32281 65744
rect 32079 65690 32095 65724
rect 32129 65690 32163 65724
rect 32197 65690 32231 65724
rect 32265 65690 32281 65724
rect 32079 65674 32281 65690
rect 32122 65652 32152 65674
rect 32208 65652 32238 65674
rect 32122 65300 32152 65322
rect 32208 65300 32238 65322
rect 32079 65284 32281 65300
rect 32079 65250 32095 65284
rect 32129 65250 32163 65284
rect 32197 65250 32231 65284
rect 32265 65250 32281 65284
rect 32079 65230 32281 65250
rect 41279 65724 41481 65744
rect 41279 65690 41295 65724
rect 41329 65690 41363 65724
rect 41397 65690 41431 65724
rect 41465 65690 41481 65724
rect 41279 65674 41481 65690
rect 41322 65652 41352 65674
rect 41408 65652 41438 65674
rect 41322 65300 41352 65322
rect 41408 65300 41438 65322
rect 41279 65284 41481 65300
rect 41279 65250 41295 65284
rect 41329 65250 41363 65284
rect 41397 65250 41431 65284
rect 41465 65250 41481 65284
rect 41279 65230 41481 65250
rect 50479 65724 50681 65744
rect 50479 65690 50495 65724
rect 50529 65690 50563 65724
rect 50597 65690 50631 65724
rect 50665 65690 50681 65724
rect 50479 65674 50681 65690
rect 50522 65652 50552 65674
rect 50608 65652 50638 65674
rect 50522 65300 50552 65322
rect 50608 65300 50638 65322
rect 50479 65284 50681 65300
rect 50479 65250 50495 65284
rect 50529 65250 50563 65284
rect 50597 65250 50631 65284
rect 50665 65250 50681 65284
rect 50479 65230 50681 65250
rect 59679 65724 59881 65744
rect 59679 65690 59695 65724
rect 59729 65690 59763 65724
rect 59797 65690 59831 65724
rect 59865 65690 59881 65724
rect 59679 65674 59881 65690
rect 59722 65652 59752 65674
rect 59808 65652 59838 65674
rect 59722 65300 59752 65322
rect 59808 65300 59838 65322
rect 59679 65284 59881 65300
rect 59679 65250 59695 65284
rect 59729 65250 59763 65284
rect 59797 65250 59831 65284
rect 59865 65250 59881 65284
rect 59679 65230 59881 65250
rect 68879 65724 69081 65744
rect 68879 65690 68895 65724
rect 68929 65690 68963 65724
rect 68997 65690 69031 65724
rect 69065 65690 69081 65724
rect 68879 65674 69081 65690
rect 68922 65652 68952 65674
rect 69008 65652 69038 65674
rect 68922 65300 68952 65322
rect 69008 65300 69038 65322
rect 68879 65284 69081 65300
rect 68879 65250 68895 65284
rect 68929 65250 68963 65284
rect 68997 65250 69031 65284
rect 69065 65250 69081 65284
rect 68879 65230 69081 65250
rect -378 65112 -348 65156
rect -240 65112 -160 65120
rect -378 65100 -160 65112
rect -378 65060 -220 65100
rect -180 65060 -160 65100
rect -378 65050 -160 65060
rect -378 65026 -348 65050
rect -240 65040 -160 65050
rect -378 64700 -348 64726
rect 4479 55844 4681 55864
rect 4479 55810 4495 55844
rect 4529 55810 4563 55844
rect 4597 55810 4631 55844
rect 4665 55810 4681 55844
rect 4479 55794 4681 55810
rect 4522 55772 4552 55794
rect 4608 55772 4638 55794
rect 4522 55420 4552 55442
rect 4608 55420 4638 55442
rect 4479 55404 4681 55420
rect 4479 55370 4495 55404
rect 4529 55370 4563 55404
rect 4597 55370 4631 55404
rect 4665 55370 4681 55404
rect 4479 55350 4681 55370
rect 13679 55844 13881 55864
rect 13679 55810 13695 55844
rect 13729 55810 13763 55844
rect 13797 55810 13831 55844
rect 13865 55810 13881 55844
rect 13679 55794 13881 55810
rect 13722 55772 13752 55794
rect 13808 55772 13838 55794
rect 13722 55420 13752 55442
rect 13808 55420 13838 55442
rect 13679 55404 13881 55420
rect 13679 55370 13695 55404
rect 13729 55370 13763 55404
rect 13797 55370 13831 55404
rect 13865 55370 13881 55404
rect 13679 55350 13881 55370
rect 22879 55844 23081 55864
rect 22879 55810 22895 55844
rect 22929 55810 22963 55844
rect 22997 55810 23031 55844
rect 23065 55810 23081 55844
rect 22879 55794 23081 55810
rect 22922 55772 22952 55794
rect 23008 55772 23038 55794
rect 22922 55420 22952 55442
rect 23008 55420 23038 55442
rect 22879 55404 23081 55420
rect 22879 55370 22895 55404
rect 22929 55370 22963 55404
rect 22997 55370 23031 55404
rect 23065 55370 23081 55404
rect 22879 55350 23081 55370
rect 32079 55844 32281 55864
rect 32079 55810 32095 55844
rect 32129 55810 32163 55844
rect 32197 55810 32231 55844
rect 32265 55810 32281 55844
rect 32079 55794 32281 55810
rect 32122 55772 32152 55794
rect 32208 55772 32238 55794
rect 32122 55420 32152 55442
rect 32208 55420 32238 55442
rect 32079 55404 32281 55420
rect 32079 55370 32095 55404
rect 32129 55370 32163 55404
rect 32197 55370 32231 55404
rect 32265 55370 32281 55404
rect 32079 55350 32281 55370
rect 41279 55844 41481 55864
rect 41279 55810 41295 55844
rect 41329 55810 41363 55844
rect 41397 55810 41431 55844
rect 41465 55810 41481 55844
rect 41279 55794 41481 55810
rect 41322 55772 41352 55794
rect 41408 55772 41438 55794
rect 41322 55420 41352 55442
rect 41408 55420 41438 55442
rect 41279 55404 41481 55420
rect 41279 55370 41295 55404
rect 41329 55370 41363 55404
rect 41397 55370 41431 55404
rect 41465 55370 41481 55404
rect 41279 55350 41481 55370
rect 50479 55844 50681 55864
rect 50479 55810 50495 55844
rect 50529 55810 50563 55844
rect 50597 55810 50631 55844
rect 50665 55810 50681 55844
rect 50479 55794 50681 55810
rect 50522 55772 50552 55794
rect 50608 55772 50638 55794
rect 50522 55420 50552 55442
rect 50608 55420 50638 55442
rect 50479 55404 50681 55420
rect 50479 55370 50495 55404
rect 50529 55370 50563 55404
rect 50597 55370 50631 55404
rect 50665 55370 50681 55404
rect 50479 55350 50681 55370
rect 59679 55844 59881 55864
rect 59679 55810 59695 55844
rect 59729 55810 59763 55844
rect 59797 55810 59831 55844
rect 59865 55810 59881 55844
rect 59679 55794 59881 55810
rect 59722 55772 59752 55794
rect 59808 55772 59838 55794
rect 59722 55420 59752 55442
rect 59808 55420 59838 55442
rect 59679 55404 59881 55420
rect 59679 55370 59695 55404
rect 59729 55370 59763 55404
rect 59797 55370 59831 55404
rect 59865 55370 59881 55404
rect 59679 55350 59881 55370
rect 68879 55844 69081 55864
rect 68879 55810 68895 55844
rect 68929 55810 68963 55844
rect 68997 55810 69031 55844
rect 69065 55810 69081 55844
rect 68879 55794 69081 55810
rect 68922 55772 68952 55794
rect 69008 55772 69038 55794
rect 68922 55420 68952 55442
rect 69008 55420 69038 55442
rect 68879 55404 69081 55420
rect 68879 55370 68895 55404
rect 68929 55370 68963 55404
rect 68997 55370 69031 55404
rect 69065 55370 69081 55404
rect 68879 55350 69081 55370
rect -378 45996 -348 46022
rect 4479 45964 4681 45984
rect 4479 45930 4495 45964
rect 4529 45930 4563 45964
rect 4597 45930 4631 45964
rect 4665 45930 4681 45964
rect 4479 45914 4681 45930
rect 4522 45892 4552 45914
rect 4608 45892 4638 45914
rect 4522 45540 4552 45562
rect 4608 45540 4638 45562
rect 4479 45524 4681 45540
rect 4479 45490 4495 45524
rect 4529 45490 4563 45524
rect 4597 45490 4631 45524
rect 4665 45490 4681 45524
rect 4479 45470 4681 45490
rect 13679 45964 13881 45984
rect 13679 45930 13695 45964
rect 13729 45930 13763 45964
rect 13797 45930 13831 45964
rect 13865 45930 13881 45964
rect 13679 45914 13881 45930
rect 13722 45892 13752 45914
rect 13808 45892 13838 45914
rect 13722 45540 13752 45562
rect 13808 45540 13838 45562
rect 13679 45524 13881 45540
rect 13679 45490 13695 45524
rect 13729 45490 13763 45524
rect 13797 45490 13831 45524
rect 13865 45490 13881 45524
rect 13679 45470 13881 45490
rect 22879 45964 23081 45984
rect 22879 45930 22895 45964
rect 22929 45930 22963 45964
rect 22997 45930 23031 45964
rect 23065 45930 23081 45964
rect 22879 45914 23081 45930
rect 22922 45892 22952 45914
rect 23008 45892 23038 45914
rect 22922 45540 22952 45562
rect 23008 45540 23038 45562
rect 22879 45524 23081 45540
rect 22879 45490 22895 45524
rect 22929 45490 22963 45524
rect 22997 45490 23031 45524
rect 23065 45490 23081 45524
rect 22879 45470 23081 45490
rect 32079 45964 32281 45984
rect 32079 45930 32095 45964
rect 32129 45930 32163 45964
rect 32197 45930 32231 45964
rect 32265 45930 32281 45964
rect 32079 45914 32281 45930
rect 32122 45892 32152 45914
rect 32208 45892 32238 45914
rect 32122 45540 32152 45562
rect 32208 45540 32238 45562
rect 32079 45524 32281 45540
rect 32079 45490 32095 45524
rect 32129 45490 32163 45524
rect 32197 45490 32231 45524
rect 32265 45490 32281 45524
rect 32079 45470 32281 45490
rect 41279 45964 41481 45984
rect 41279 45930 41295 45964
rect 41329 45930 41363 45964
rect 41397 45930 41431 45964
rect 41465 45930 41481 45964
rect 41279 45914 41481 45930
rect 41322 45892 41352 45914
rect 41408 45892 41438 45914
rect 41322 45540 41352 45562
rect 41408 45540 41438 45562
rect 41279 45524 41481 45540
rect 41279 45490 41295 45524
rect 41329 45490 41363 45524
rect 41397 45490 41431 45524
rect 41465 45490 41481 45524
rect 41279 45470 41481 45490
rect 50479 45964 50681 45984
rect 50479 45930 50495 45964
rect 50529 45930 50563 45964
rect 50597 45930 50631 45964
rect 50665 45930 50681 45964
rect 50479 45914 50681 45930
rect 50522 45892 50552 45914
rect 50608 45892 50638 45914
rect 50522 45540 50552 45562
rect 50608 45540 50638 45562
rect 50479 45524 50681 45540
rect 50479 45490 50495 45524
rect 50529 45490 50563 45524
rect 50597 45490 50631 45524
rect 50665 45490 50681 45524
rect 50479 45470 50681 45490
rect 59679 45964 59881 45984
rect 59679 45930 59695 45964
rect 59729 45930 59763 45964
rect 59797 45930 59831 45964
rect 59865 45930 59881 45964
rect 59679 45914 59881 45930
rect 59722 45892 59752 45914
rect 59808 45892 59838 45914
rect 59722 45540 59752 45562
rect 59808 45540 59838 45562
rect 59679 45524 59881 45540
rect 59679 45490 59695 45524
rect 59729 45490 59763 45524
rect 59797 45490 59831 45524
rect 59865 45490 59881 45524
rect 59679 45470 59881 45490
rect 68879 45964 69081 45984
rect 68879 45930 68895 45964
rect 68929 45930 68963 45964
rect 68997 45930 69031 45964
rect 69065 45930 69081 45964
rect 68879 45914 69081 45930
rect 68922 45892 68952 45914
rect 69008 45892 69038 45914
rect 68922 45540 68952 45562
rect 69008 45540 69038 45562
rect 68879 45524 69081 45540
rect 68879 45490 68895 45524
rect 68929 45490 68963 45524
rect 68997 45490 69031 45524
rect 69065 45490 69081 45524
rect 68879 45470 69081 45490
rect -378 45352 -348 45396
rect -240 45352 -160 45360
rect -378 45340 -160 45352
rect -378 45300 -220 45340
rect -180 45300 -160 45340
rect -378 45290 -160 45300
rect -378 45266 -348 45290
rect -240 45280 -160 45290
rect -378 44940 -348 44966
rect 4479 36084 4681 36104
rect 4479 36050 4495 36084
rect 4529 36050 4563 36084
rect 4597 36050 4631 36084
rect 4665 36050 4681 36084
rect 4479 36034 4681 36050
rect 4522 36012 4552 36034
rect 4608 36012 4638 36034
rect 4522 35660 4552 35682
rect 4608 35660 4638 35682
rect 4479 35644 4681 35660
rect 4479 35610 4495 35644
rect 4529 35610 4563 35644
rect 4597 35610 4631 35644
rect 4665 35610 4681 35644
rect 4479 35590 4681 35610
rect 13679 36084 13881 36104
rect 13679 36050 13695 36084
rect 13729 36050 13763 36084
rect 13797 36050 13831 36084
rect 13865 36050 13881 36084
rect 13679 36034 13881 36050
rect 13722 36012 13752 36034
rect 13808 36012 13838 36034
rect 13722 35660 13752 35682
rect 13808 35660 13838 35682
rect 13679 35644 13881 35660
rect 13679 35610 13695 35644
rect 13729 35610 13763 35644
rect 13797 35610 13831 35644
rect 13865 35610 13881 35644
rect 13679 35590 13881 35610
rect 22879 36084 23081 36104
rect 22879 36050 22895 36084
rect 22929 36050 22963 36084
rect 22997 36050 23031 36084
rect 23065 36050 23081 36084
rect 22879 36034 23081 36050
rect 22922 36012 22952 36034
rect 23008 36012 23038 36034
rect 22922 35660 22952 35682
rect 23008 35660 23038 35682
rect 22879 35644 23081 35660
rect 22879 35610 22895 35644
rect 22929 35610 22963 35644
rect 22997 35610 23031 35644
rect 23065 35610 23081 35644
rect 22879 35590 23081 35610
rect 32079 36084 32281 36104
rect 32079 36050 32095 36084
rect 32129 36050 32163 36084
rect 32197 36050 32231 36084
rect 32265 36050 32281 36084
rect 32079 36034 32281 36050
rect 32122 36012 32152 36034
rect 32208 36012 32238 36034
rect 32122 35660 32152 35682
rect 32208 35660 32238 35682
rect 32079 35644 32281 35660
rect 32079 35610 32095 35644
rect 32129 35610 32163 35644
rect 32197 35610 32231 35644
rect 32265 35610 32281 35644
rect 32079 35590 32281 35610
rect 41279 36084 41481 36104
rect 41279 36050 41295 36084
rect 41329 36050 41363 36084
rect 41397 36050 41431 36084
rect 41465 36050 41481 36084
rect 41279 36034 41481 36050
rect 41322 36012 41352 36034
rect 41408 36012 41438 36034
rect 41322 35660 41352 35682
rect 41408 35660 41438 35682
rect 41279 35644 41481 35660
rect 41279 35610 41295 35644
rect 41329 35610 41363 35644
rect 41397 35610 41431 35644
rect 41465 35610 41481 35644
rect 41279 35590 41481 35610
rect 50479 36084 50681 36104
rect 50479 36050 50495 36084
rect 50529 36050 50563 36084
rect 50597 36050 50631 36084
rect 50665 36050 50681 36084
rect 50479 36034 50681 36050
rect 50522 36012 50552 36034
rect 50608 36012 50638 36034
rect 50522 35660 50552 35682
rect 50608 35660 50638 35682
rect 50479 35644 50681 35660
rect 50479 35610 50495 35644
rect 50529 35610 50563 35644
rect 50597 35610 50631 35644
rect 50665 35610 50681 35644
rect 50479 35590 50681 35610
rect 59679 36084 59881 36104
rect 59679 36050 59695 36084
rect 59729 36050 59763 36084
rect 59797 36050 59831 36084
rect 59865 36050 59881 36084
rect 59679 36034 59881 36050
rect 59722 36012 59752 36034
rect 59808 36012 59838 36034
rect 59722 35660 59752 35682
rect 59808 35660 59838 35682
rect 59679 35644 59881 35660
rect 59679 35610 59695 35644
rect 59729 35610 59763 35644
rect 59797 35610 59831 35644
rect 59865 35610 59881 35644
rect 59679 35590 59881 35610
rect 68879 36084 69081 36104
rect 68879 36050 68895 36084
rect 68929 36050 68963 36084
rect 68997 36050 69031 36084
rect 69065 36050 69081 36084
rect 68879 36034 69081 36050
rect 68922 36012 68952 36034
rect 69008 36012 69038 36034
rect 68922 35660 68952 35682
rect 69008 35660 69038 35682
rect 68879 35644 69081 35660
rect 68879 35610 68895 35644
rect 68929 35610 68963 35644
rect 68997 35610 69031 35644
rect 69065 35610 69081 35644
rect 68879 35590 69081 35610
rect 4479 26204 4681 26224
rect 4479 26170 4495 26204
rect 4529 26170 4563 26204
rect 4597 26170 4631 26204
rect 4665 26170 4681 26204
rect 4479 26154 4681 26170
rect 4522 26132 4552 26154
rect 4608 26132 4638 26154
rect 4522 25780 4552 25802
rect 4608 25780 4638 25802
rect 4479 25764 4681 25780
rect 4479 25730 4495 25764
rect 4529 25730 4563 25764
rect 4597 25730 4631 25764
rect 4665 25730 4681 25764
rect 4479 25710 4681 25730
rect 13679 26204 13881 26224
rect 13679 26170 13695 26204
rect 13729 26170 13763 26204
rect 13797 26170 13831 26204
rect 13865 26170 13881 26204
rect 13679 26154 13881 26170
rect 13722 26132 13752 26154
rect 13808 26132 13838 26154
rect 13722 25780 13752 25802
rect 13808 25780 13838 25802
rect 13679 25764 13881 25780
rect 13679 25730 13695 25764
rect 13729 25730 13763 25764
rect 13797 25730 13831 25764
rect 13865 25730 13881 25764
rect 13679 25710 13881 25730
rect 22879 26204 23081 26224
rect 22879 26170 22895 26204
rect 22929 26170 22963 26204
rect 22997 26170 23031 26204
rect 23065 26170 23081 26204
rect 22879 26154 23081 26170
rect 22922 26132 22952 26154
rect 23008 26132 23038 26154
rect 22922 25780 22952 25802
rect 23008 25780 23038 25802
rect 22879 25764 23081 25780
rect 22879 25730 22895 25764
rect 22929 25730 22963 25764
rect 22997 25730 23031 25764
rect 23065 25730 23081 25764
rect 22879 25710 23081 25730
rect 32079 26204 32281 26224
rect 32079 26170 32095 26204
rect 32129 26170 32163 26204
rect 32197 26170 32231 26204
rect 32265 26170 32281 26204
rect 32079 26154 32281 26170
rect 32122 26132 32152 26154
rect 32208 26132 32238 26154
rect 32122 25780 32152 25802
rect 32208 25780 32238 25802
rect 32079 25764 32281 25780
rect 32079 25730 32095 25764
rect 32129 25730 32163 25764
rect 32197 25730 32231 25764
rect 32265 25730 32281 25764
rect 32079 25710 32281 25730
rect 41279 26204 41481 26224
rect 41279 26170 41295 26204
rect 41329 26170 41363 26204
rect 41397 26170 41431 26204
rect 41465 26170 41481 26204
rect 41279 26154 41481 26170
rect 41322 26132 41352 26154
rect 41408 26132 41438 26154
rect 41322 25780 41352 25802
rect 41408 25780 41438 25802
rect 41279 25764 41481 25780
rect 41279 25730 41295 25764
rect 41329 25730 41363 25764
rect 41397 25730 41431 25764
rect 41465 25730 41481 25764
rect 41279 25710 41481 25730
rect 50479 26204 50681 26224
rect 50479 26170 50495 26204
rect 50529 26170 50563 26204
rect 50597 26170 50631 26204
rect 50665 26170 50681 26204
rect 50479 26154 50681 26170
rect 50522 26132 50552 26154
rect 50608 26132 50638 26154
rect 50522 25780 50552 25802
rect 50608 25780 50638 25802
rect 50479 25764 50681 25780
rect 50479 25730 50495 25764
rect 50529 25730 50563 25764
rect 50597 25730 50631 25764
rect 50665 25730 50681 25764
rect 50479 25710 50681 25730
rect 59679 26204 59881 26224
rect 59679 26170 59695 26204
rect 59729 26170 59763 26204
rect 59797 26170 59831 26204
rect 59865 26170 59881 26204
rect 59679 26154 59881 26170
rect 59722 26132 59752 26154
rect 59808 26132 59838 26154
rect 59722 25780 59752 25802
rect 59808 25780 59838 25802
rect 59679 25764 59881 25780
rect 59679 25730 59695 25764
rect 59729 25730 59763 25764
rect 59797 25730 59831 25764
rect 59865 25730 59881 25764
rect 59679 25710 59881 25730
rect 68879 26204 69081 26224
rect 68879 26170 68895 26204
rect 68929 26170 68963 26204
rect 68997 26170 69031 26204
rect 69065 26170 69081 26204
rect 68879 26154 69081 26170
rect 68922 26132 68952 26154
rect 69008 26132 69038 26154
rect 68922 25780 68952 25802
rect 69008 25780 69038 25802
rect 68879 25764 69081 25780
rect 68879 25730 68895 25764
rect 68929 25730 68963 25764
rect 68997 25730 69031 25764
rect 69065 25730 69081 25764
rect 68879 25710 69081 25730
rect 4479 16324 4681 16344
rect 4479 16290 4495 16324
rect 4529 16290 4563 16324
rect 4597 16290 4631 16324
rect 4665 16290 4681 16324
rect 4479 16274 4681 16290
rect 4522 16252 4552 16274
rect 4608 16252 4638 16274
rect 4522 15900 4552 15922
rect 4608 15900 4638 15922
rect 4479 15884 4681 15900
rect 4479 15850 4495 15884
rect 4529 15850 4563 15884
rect 4597 15850 4631 15884
rect 4665 15850 4681 15884
rect 4479 15830 4681 15850
rect 13679 16324 13881 16344
rect 13679 16290 13695 16324
rect 13729 16290 13763 16324
rect 13797 16290 13831 16324
rect 13865 16290 13881 16324
rect 13679 16274 13881 16290
rect 13722 16252 13752 16274
rect 13808 16252 13838 16274
rect 13722 15900 13752 15922
rect 13808 15900 13838 15922
rect 13679 15884 13881 15900
rect 13679 15850 13695 15884
rect 13729 15850 13763 15884
rect 13797 15850 13831 15884
rect 13865 15850 13881 15884
rect 13679 15830 13881 15850
rect 22879 16324 23081 16344
rect 22879 16290 22895 16324
rect 22929 16290 22963 16324
rect 22997 16290 23031 16324
rect 23065 16290 23081 16324
rect 22879 16274 23081 16290
rect 22922 16252 22952 16274
rect 23008 16252 23038 16274
rect 22922 15900 22952 15922
rect 23008 15900 23038 15922
rect 22879 15884 23081 15900
rect 22879 15850 22895 15884
rect 22929 15850 22963 15884
rect 22997 15850 23031 15884
rect 23065 15850 23081 15884
rect 22879 15830 23081 15850
rect 32079 16324 32281 16344
rect 32079 16290 32095 16324
rect 32129 16290 32163 16324
rect 32197 16290 32231 16324
rect 32265 16290 32281 16324
rect 32079 16274 32281 16290
rect 32122 16252 32152 16274
rect 32208 16252 32238 16274
rect 32122 15900 32152 15922
rect 32208 15900 32238 15922
rect 32079 15884 32281 15900
rect 32079 15850 32095 15884
rect 32129 15850 32163 15884
rect 32197 15850 32231 15884
rect 32265 15850 32281 15884
rect 32079 15830 32281 15850
rect 41279 16324 41481 16344
rect 41279 16290 41295 16324
rect 41329 16290 41363 16324
rect 41397 16290 41431 16324
rect 41465 16290 41481 16324
rect 41279 16274 41481 16290
rect 41322 16252 41352 16274
rect 41408 16252 41438 16274
rect 41322 15900 41352 15922
rect 41408 15900 41438 15922
rect 41279 15884 41481 15900
rect 41279 15850 41295 15884
rect 41329 15850 41363 15884
rect 41397 15850 41431 15884
rect 41465 15850 41481 15884
rect 41279 15830 41481 15850
rect 50479 16324 50681 16344
rect 50479 16290 50495 16324
rect 50529 16290 50563 16324
rect 50597 16290 50631 16324
rect 50665 16290 50681 16324
rect 50479 16274 50681 16290
rect 50522 16252 50552 16274
rect 50608 16252 50638 16274
rect 50522 15900 50552 15922
rect 50608 15900 50638 15922
rect 50479 15884 50681 15900
rect 50479 15850 50495 15884
rect 50529 15850 50563 15884
rect 50597 15850 50631 15884
rect 50665 15850 50681 15884
rect 50479 15830 50681 15850
rect 59679 16324 59881 16344
rect 59679 16290 59695 16324
rect 59729 16290 59763 16324
rect 59797 16290 59831 16324
rect 59865 16290 59881 16324
rect 59679 16274 59881 16290
rect 59722 16252 59752 16274
rect 59808 16252 59838 16274
rect 59722 15900 59752 15922
rect 59808 15900 59838 15922
rect 59679 15884 59881 15900
rect 59679 15850 59695 15884
rect 59729 15850 59763 15884
rect 59797 15850 59831 15884
rect 59865 15850 59881 15884
rect 59679 15830 59881 15850
rect 68879 16324 69081 16344
rect 68879 16290 68895 16324
rect 68929 16290 68963 16324
rect 68997 16290 69031 16324
rect 69065 16290 69081 16324
rect 68879 16274 69081 16290
rect 68922 16252 68952 16274
rect 69008 16252 69038 16274
rect 68922 15900 68952 15922
rect 69008 15900 69038 15922
rect 68879 15884 69081 15900
rect 68879 15850 68895 15884
rect 68929 15850 68963 15884
rect 68997 15850 69031 15884
rect 69065 15850 69081 15884
rect 68879 15830 69081 15850
rect -378 6476 -348 6502
rect 4479 6444 4681 6464
rect 4479 6410 4495 6444
rect 4529 6410 4563 6444
rect 4597 6410 4631 6444
rect 4665 6410 4681 6444
rect 4479 6394 4681 6410
rect 4522 6372 4552 6394
rect 4608 6372 4638 6394
rect 4522 6020 4552 6042
rect 4608 6020 4638 6042
rect 4479 6004 4681 6020
rect 4479 5970 4495 6004
rect 4529 5970 4563 6004
rect 4597 5970 4631 6004
rect 4665 5970 4681 6004
rect 4479 5950 4681 5970
rect 13679 6444 13881 6464
rect 13679 6410 13695 6444
rect 13729 6410 13763 6444
rect 13797 6410 13831 6444
rect 13865 6410 13881 6444
rect 13679 6394 13881 6410
rect 13722 6372 13752 6394
rect 13808 6372 13838 6394
rect 13722 6020 13752 6042
rect 13808 6020 13838 6042
rect 13679 6004 13881 6020
rect 13679 5970 13695 6004
rect 13729 5970 13763 6004
rect 13797 5970 13831 6004
rect 13865 5970 13881 6004
rect 13679 5950 13881 5970
rect 22879 6444 23081 6464
rect 22879 6410 22895 6444
rect 22929 6410 22963 6444
rect 22997 6410 23031 6444
rect 23065 6410 23081 6444
rect 22879 6394 23081 6410
rect 22922 6372 22952 6394
rect 23008 6372 23038 6394
rect 22922 6020 22952 6042
rect 23008 6020 23038 6042
rect 22879 6004 23081 6020
rect 22879 5970 22895 6004
rect 22929 5970 22963 6004
rect 22997 5970 23031 6004
rect 23065 5970 23081 6004
rect 22879 5950 23081 5970
rect 32079 6444 32281 6464
rect 32079 6410 32095 6444
rect 32129 6410 32163 6444
rect 32197 6410 32231 6444
rect 32265 6410 32281 6444
rect 32079 6394 32281 6410
rect 32122 6372 32152 6394
rect 32208 6372 32238 6394
rect 32122 6020 32152 6042
rect 32208 6020 32238 6042
rect 32079 6004 32281 6020
rect 32079 5970 32095 6004
rect 32129 5970 32163 6004
rect 32197 5970 32231 6004
rect 32265 5970 32281 6004
rect 32079 5950 32281 5970
rect 41279 6444 41481 6464
rect 41279 6410 41295 6444
rect 41329 6410 41363 6444
rect 41397 6410 41431 6444
rect 41465 6410 41481 6444
rect 41279 6394 41481 6410
rect 41322 6372 41352 6394
rect 41408 6372 41438 6394
rect 41322 6020 41352 6042
rect 41408 6020 41438 6042
rect 41279 6004 41481 6020
rect 41279 5970 41295 6004
rect 41329 5970 41363 6004
rect 41397 5970 41431 6004
rect 41465 5970 41481 6004
rect 41279 5950 41481 5970
rect 50479 6444 50681 6464
rect 50479 6410 50495 6444
rect 50529 6410 50563 6444
rect 50597 6410 50631 6444
rect 50665 6410 50681 6444
rect 50479 6394 50681 6410
rect 50522 6372 50552 6394
rect 50608 6372 50638 6394
rect 50522 6020 50552 6042
rect 50608 6020 50638 6042
rect 50479 6004 50681 6020
rect 50479 5970 50495 6004
rect 50529 5970 50563 6004
rect 50597 5970 50631 6004
rect 50665 5970 50681 6004
rect 50479 5950 50681 5970
rect 59679 6444 59881 6464
rect 59679 6410 59695 6444
rect 59729 6410 59763 6444
rect 59797 6410 59831 6444
rect 59865 6410 59881 6444
rect 59679 6394 59881 6410
rect 59722 6372 59752 6394
rect 59808 6372 59838 6394
rect 59722 6020 59752 6042
rect 59808 6020 59838 6042
rect 59679 6004 59881 6020
rect 59679 5970 59695 6004
rect 59729 5970 59763 6004
rect 59797 5970 59831 6004
rect 59865 5970 59881 6004
rect 59679 5950 59881 5970
rect 68879 6444 69081 6464
rect 68879 6410 68895 6444
rect 68929 6410 68963 6444
rect 68997 6410 69031 6444
rect 69065 6410 69081 6444
rect 68879 6394 69081 6410
rect 68922 6372 68952 6394
rect 69008 6372 69038 6394
rect 68922 6020 68952 6042
rect 69008 6020 69038 6042
rect 68879 6004 69081 6020
rect 68879 5970 68895 6004
rect 68929 5970 68963 6004
rect 68997 5970 69031 6004
rect 69065 5970 69081 6004
rect 68879 5950 69081 5970
rect -378 5832 -348 5876
rect -240 5832 -160 5840
rect -378 5820 -160 5832
rect -378 5780 -220 5820
rect -180 5780 -160 5820
rect -378 5770 -160 5780
rect -378 5746 -348 5770
rect -240 5760 -160 5770
rect -378 5420 -348 5446
<< polycont >>
rect 4495 95330 4529 95364
rect 4563 95330 4597 95364
rect 4631 95330 4665 95364
rect 4495 94890 4529 94924
rect 4563 94890 4597 94924
rect 4631 94890 4665 94924
rect -220 94700 -180 94740
rect 4495 85450 4529 85484
rect 4563 85450 4597 85484
rect 4631 85450 4665 85484
rect 4495 85010 4529 85044
rect 4563 85010 4597 85044
rect 4631 85010 4665 85044
rect 13695 85450 13729 85484
rect 13763 85450 13797 85484
rect 13831 85450 13865 85484
rect 13695 85010 13729 85044
rect 13763 85010 13797 85044
rect 13831 85010 13865 85044
rect -220 84820 -180 84860
rect 4495 75570 4529 75604
rect 4563 75570 4597 75604
rect 4631 75570 4665 75604
rect 4495 75130 4529 75164
rect 4563 75130 4597 75164
rect 4631 75130 4665 75164
rect 13695 75570 13729 75604
rect 13763 75570 13797 75604
rect 13831 75570 13865 75604
rect 13695 75130 13729 75164
rect 13763 75130 13797 75164
rect 13831 75130 13865 75164
rect 22895 75570 22929 75604
rect 22963 75570 22997 75604
rect 23031 75570 23065 75604
rect 22895 75130 22929 75164
rect 22963 75130 22997 75164
rect 23031 75130 23065 75164
rect 32095 75570 32129 75604
rect 32163 75570 32197 75604
rect 32231 75570 32265 75604
rect 32095 75130 32129 75164
rect 32163 75130 32197 75164
rect 32231 75130 32265 75164
rect -220 74940 -180 74980
rect 4495 65690 4529 65724
rect 4563 65690 4597 65724
rect 4631 65690 4665 65724
rect 4495 65250 4529 65284
rect 4563 65250 4597 65284
rect 4631 65250 4665 65284
rect 13695 65690 13729 65724
rect 13763 65690 13797 65724
rect 13831 65690 13865 65724
rect 13695 65250 13729 65284
rect 13763 65250 13797 65284
rect 13831 65250 13865 65284
rect 22895 65690 22929 65724
rect 22963 65690 22997 65724
rect 23031 65690 23065 65724
rect 22895 65250 22929 65284
rect 22963 65250 22997 65284
rect 23031 65250 23065 65284
rect 32095 65690 32129 65724
rect 32163 65690 32197 65724
rect 32231 65690 32265 65724
rect 32095 65250 32129 65284
rect 32163 65250 32197 65284
rect 32231 65250 32265 65284
rect 41295 65690 41329 65724
rect 41363 65690 41397 65724
rect 41431 65690 41465 65724
rect 41295 65250 41329 65284
rect 41363 65250 41397 65284
rect 41431 65250 41465 65284
rect 50495 65690 50529 65724
rect 50563 65690 50597 65724
rect 50631 65690 50665 65724
rect 50495 65250 50529 65284
rect 50563 65250 50597 65284
rect 50631 65250 50665 65284
rect 59695 65690 59729 65724
rect 59763 65690 59797 65724
rect 59831 65690 59865 65724
rect 59695 65250 59729 65284
rect 59763 65250 59797 65284
rect 59831 65250 59865 65284
rect 68895 65690 68929 65724
rect 68963 65690 68997 65724
rect 69031 65690 69065 65724
rect 68895 65250 68929 65284
rect 68963 65250 68997 65284
rect 69031 65250 69065 65284
rect -220 65060 -180 65100
rect 4495 55810 4529 55844
rect 4563 55810 4597 55844
rect 4631 55810 4665 55844
rect 4495 55370 4529 55404
rect 4563 55370 4597 55404
rect 4631 55370 4665 55404
rect 13695 55810 13729 55844
rect 13763 55810 13797 55844
rect 13831 55810 13865 55844
rect 13695 55370 13729 55404
rect 13763 55370 13797 55404
rect 13831 55370 13865 55404
rect 22895 55810 22929 55844
rect 22963 55810 22997 55844
rect 23031 55810 23065 55844
rect 22895 55370 22929 55404
rect 22963 55370 22997 55404
rect 23031 55370 23065 55404
rect 32095 55810 32129 55844
rect 32163 55810 32197 55844
rect 32231 55810 32265 55844
rect 32095 55370 32129 55404
rect 32163 55370 32197 55404
rect 32231 55370 32265 55404
rect 41295 55810 41329 55844
rect 41363 55810 41397 55844
rect 41431 55810 41465 55844
rect 41295 55370 41329 55404
rect 41363 55370 41397 55404
rect 41431 55370 41465 55404
rect 50495 55810 50529 55844
rect 50563 55810 50597 55844
rect 50631 55810 50665 55844
rect 50495 55370 50529 55404
rect 50563 55370 50597 55404
rect 50631 55370 50665 55404
rect 59695 55810 59729 55844
rect 59763 55810 59797 55844
rect 59831 55810 59865 55844
rect 59695 55370 59729 55404
rect 59763 55370 59797 55404
rect 59831 55370 59865 55404
rect 68895 55810 68929 55844
rect 68963 55810 68997 55844
rect 69031 55810 69065 55844
rect 68895 55370 68929 55404
rect 68963 55370 68997 55404
rect 69031 55370 69065 55404
rect 4495 45930 4529 45964
rect 4563 45930 4597 45964
rect 4631 45930 4665 45964
rect 4495 45490 4529 45524
rect 4563 45490 4597 45524
rect 4631 45490 4665 45524
rect 13695 45930 13729 45964
rect 13763 45930 13797 45964
rect 13831 45930 13865 45964
rect 13695 45490 13729 45524
rect 13763 45490 13797 45524
rect 13831 45490 13865 45524
rect 22895 45930 22929 45964
rect 22963 45930 22997 45964
rect 23031 45930 23065 45964
rect 22895 45490 22929 45524
rect 22963 45490 22997 45524
rect 23031 45490 23065 45524
rect 32095 45930 32129 45964
rect 32163 45930 32197 45964
rect 32231 45930 32265 45964
rect 32095 45490 32129 45524
rect 32163 45490 32197 45524
rect 32231 45490 32265 45524
rect 41295 45930 41329 45964
rect 41363 45930 41397 45964
rect 41431 45930 41465 45964
rect 41295 45490 41329 45524
rect 41363 45490 41397 45524
rect 41431 45490 41465 45524
rect 50495 45930 50529 45964
rect 50563 45930 50597 45964
rect 50631 45930 50665 45964
rect 50495 45490 50529 45524
rect 50563 45490 50597 45524
rect 50631 45490 50665 45524
rect 59695 45930 59729 45964
rect 59763 45930 59797 45964
rect 59831 45930 59865 45964
rect 59695 45490 59729 45524
rect 59763 45490 59797 45524
rect 59831 45490 59865 45524
rect 68895 45930 68929 45964
rect 68963 45930 68997 45964
rect 69031 45930 69065 45964
rect 68895 45490 68929 45524
rect 68963 45490 68997 45524
rect 69031 45490 69065 45524
rect -220 45300 -180 45340
rect 4495 36050 4529 36084
rect 4563 36050 4597 36084
rect 4631 36050 4665 36084
rect 4495 35610 4529 35644
rect 4563 35610 4597 35644
rect 4631 35610 4665 35644
rect 13695 36050 13729 36084
rect 13763 36050 13797 36084
rect 13831 36050 13865 36084
rect 13695 35610 13729 35644
rect 13763 35610 13797 35644
rect 13831 35610 13865 35644
rect 22895 36050 22929 36084
rect 22963 36050 22997 36084
rect 23031 36050 23065 36084
rect 22895 35610 22929 35644
rect 22963 35610 22997 35644
rect 23031 35610 23065 35644
rect 32095 36050 32129 36084
rect 32163 36050 32197 36084
rect 32231 36050 32265 36084
rect 32095 35610 32129 35644
rect 32163 35610 32197 35644
rect 32231 35610 32265 35644
rect 41295 36050 41329 36084
rect 41363 36050 41397 36084
rect 41431 36050 41465 36084
rect 41295 35610 41329 35644
rect 41363 35610 41397 35644
rect 41431 35610 41465 35644
rect 50495 36050 50529 36084
rect 50563 36050 50597 36084
rect 50631 36050 50665 36084
rect 50495 35610 50529 35644
rect 50563 35610 50597 35644
rect 50631 35610 50665 35644
rect 59695 36050 59729 36084
rect 59763 36050 59797 36084
rect 59831 36050 59865 36084
rect 59695 35610 59729 35644
rect 59763 35610 59797 35644
rect 59831 35610 59865 35644
rect 68895 36050 68929 36084
rect 68963 36050 68997 36084
rect 69031 36050 69065 36084
rect 68895 35610 68929 35644
rect 68963 35610 68997 35644
rect 69031 35610 69065 35644
rect 4495 26170 4529 26204
rect 4563 26170 4597 26204
rect 4631 26170 4665 26204
rect 4495 25730 4529 25764
rect 4563 25730 4597 25764
rect 4631 25730 4665 25764
rect 13695 26170 13729 26204
rect 13763 26170 13797 26204
rect 13831 26170 13865 26204
rect 13695 25730 13729 25764
rect 13763 25730 13797 25764
rect 13831 25730 13865 25764
rect 22895 26170 22929 26204
rect 22963 26170 22997 26204
rect 23031 26170 23065 26204
rect 22895 25730 22929 25764
rect 22963 25730 22997 25764
rect 23031 25730 23065 25764
rect 32095 26170 32129 26204
rect 32163 26170 32197 26204
rect 32231 26170 32265 26204
rect 32095 25730 32129 25764
rect 32163 25730 32197 25764
rect 32231 25730 32265 25764
rect 41295 26170 41329 26204
rect 41363 26170 41397 26204
rect 41431 26170 41465 26204
rect 41295 25730 41329 25764
rect 41363 25730 41397 25764
rect 41431 25730 41465 25764
rect 50495 26170 50529 26204
rect 50563 26170 50597 26204
rect 50631 26170 50665 26204
rect 50495 25730 50529 25764
rect 50563 25730 50597 25764
rect 50631 25730 50665 25764
rect 59695 26170 59729 26204
rect 59763 26170 59797 26204
rect 59831 26170 59865 26204
rect 59695 25730 59729 25764
rect 59763 25730 59797 25764
rect 59831 25730 59865 25764
rect 68895 26170 68929 26204
rect 68963 26170 68997 26204
rect 69031 26170 69065 26204
rect 68895 25730 68929 25764
rect 68963 25730 68997 25764
rect 69031 25730 69065 25764
rect 4495 16290 4529 16324
rect 4563 16290 4597 16324
rect 4631 16290 4665 16324
rect 4495 15850 4529 15884
rect 4563 15850 4597 15884
rect 4631 15850 4665 15884
rect 13695 16290 13729 16324
rect 13763 16290 13797 16324
rect 13831 16290 13865 16324
rect 13695 15850 13729 15884
rect 13763 15850 13797 15884
rect 13831 15850 13865 15884
rect 22895 16290 22929 16324
rect 22963 16290 22997 16324
rect 23031 16290 23065 16324
rect 22895 15850 22929 15884
rect 22963 15850 22997 15884
rect 23031 15850 23065 15884
rect 32095 16290 32129 16324
rect 32163 16290 32197 16324
rect 32231 16290 32265 16324
rect 32095 15850 32129 15884
rect 32163 15850 32197 15884
rect 32231 15850 32265 15884
rect 41295 16290 41329 16324
rect 41363 16290 41397 16324
rect 41431 16290 41465 16324
rect 41295 15850 41329 15884
rect 41363 15850 41397 15884
rect 41431 15850 41465 15884
rect 50495 16290 50529 16324
rect 50563 16290 50597 16324
rect 50631 16290 50665 16324
rect 50495 15850 50529 15884
rect 50563 15850 50597 15884
rect 50631 15850 50665 15884
rect 59695 16290 59729 16324
rect 59763 16290 59797 16324
rect 59831 16290 59865 16324
rect 59695 15850 59729 15884
rect 59763 15850 59797 15884
rect 59831 15850 59865 15884
rect 68895 16290 68929 16324
rect 68963 16290 68997 16324
rect 69031 16290 69065 16324
rect 68895 15850 68929 15884
rect 68963 15850 68997 15884
rect 69031 15850 69065 15884
rect 4495 6410 4529 6444
rect 4563 6410 4597 6444
rect 4631 6410 4665 6444
rect 4495 5970 4529 6004
rect 4563 5970 4597 6004
rect 4631 5970 4665 6004
rect 13695 6410 13729 6444
rect 13763 6410 13797 6444
rect 13831 6410 13865 6444
rect 13695 5970 13729 6004
rect 13763 5970 13797 6004
rect 13831 5970 13865 6004
rect 22895 6410 22929 6444
rect 22963 6410 22997 6444
rect 23031 6410 23065 6444
rect 22895 5970 22929 6004
rect 22963 5970 22997 6004
rect 23031 5970 23065 6004
rect 32095 6410 32129 6444
rect 32163 6410 32197 6444
rect 32231 6410 32265 6444
rect 32095 5970 32129 6004
rect 32163 5970 32197 6004
rect 32231 5970 32265 6004
rect 41295 6410 41329 6444
rect 41363 6410 41397 6444
rect 41431 6410 41465 6444
rect 41295 5970 41329 6004
rect 41363 5970 41397 6004
rect 41431 5970 41465 6004
rect 50495 6410 50529 6444
rect 50563 6410 50597 6444
rect 50631 6410 50665 6444
rect 50495 5970 50529 6004
rect 50563 5970 50597 6004
rect 50631 5970 50665 6004
rect 59695 6410 59729 6444
rect 59763 6410 59797 6444
rect 59831 6410 59865 6444
rect 59695 5970 59729 6004
rect 59763 5970 59797 6004
rect 59831 5970 59865 6004
rect 68895 6410 68929 6444
rect 68963 6410 68997 6444
rect 69031 6410 69065 6444
rect 68895 5970 68929 6004
rect 68963 5970 68997 6004
rect 69031 5970 69065 6004
rect -220 5780 -180 5820
<< xpolycontact >>
rect 4176 95518 4246 95950
rect 4914 95518 4984 95950
rect 4176 94886 4246 95318
rect 4914 94886 4984 95318
rect 4176 85638 4246 86070
rect 4914 85638 4984 86070
rect 4176 85006 4246 85438
rect 4914 85006 4984 85438
rect 13376 85638 13446 86070
rect 14114 85638 14184 86070
rect 13376 85006 13446 85438
rect 14114 85006 14184 85438
rect 4176 75758 4246 76190
rect 4914 75758 4984 76190
rect 4176 75126 4246 75558
rect 4914 75126 4984 75558
rect 13376 75758 13446 76190
rect 14114 75758 14184 76190
rect 13376 75126 13446 75558
rect 14114 75126 14184 75558
rect 22576 75758 22646 76190
rect 23314 75758 23384 76190
rect 22576 75126 22646 75558
rect 23314 75126 23384 75558
rect 31776 75758 31846 76190
rect 32514 75758 32584 76190
rect 31776 75126 31846 75558
rect 32514 75126 32584 75558
rect 4176 65878 4246 66310
rect 4914 65878 4984 66310
rect 4176 65246 4246 65678
rect 4914 65246 4984 65678
rect 13376 65878 13446 66310
rect 14114 65878 14184 66310
rect 13376 65246 13446 65678
rect 14114 65246 14184 65678
rect 22576 65878 22646 66310
rect 23314 65878 23384 66310
rect 22576 65246 22646 65678
rect 23314 65246 23384 65678
rect 31776 65878 31846 66310
rect 32514 65878 32584 66310
rect 31776 65246 31846 65678
rect 32514 65246 32584 65678
rect 40976 65878 41046 66310
rect 41714 65878 41784 66310
rect 40976 65246 41046 65678
rect 41714 65246 41784 65678
rect 50176 65878 50246 66310
rect 50914 65878 50984 66310
rect 50176 65246 50246 65678
rect 50914 65246 50984 65678
rect 59376 65878 59446 66310
rect 60114 65878 60184 66310
rect 59376 65246 59446 65678
rect 60114 65246 60184 65678
rect 68576 65878 68646 66310
rect 69314 65878 69384 66310
rect 68576 65246 68646 65678
rect 69314 65246 69384 65678
rect 4176 55998 4246 56430
rect 4914 55998 4984 56430
rect 4176 55366 4246 55798
rect 4914 55366 4984 55798
rect 13376 55998 13446 56430
rect 14114 55998 14184 56430
rect 13376 55366 13446 55798
rect 14114 55366 14184 55798
rect 22576 55998 22646 56430
rect 23314 55998 23384 56430
rect 22576 55366 22646 55798
rect 23314 55366 23384 55798
rect 31776 55998 31846 56430
rect 32514 55998 32584 56430
rect 31776 55366 31846 55798
rect 32514 55366 32584 55798
rect 40976 55998 41046 56430
rect 41714 55998 41784 56430
rect 40976 55366 41046 55798
rect 41714 55366 41784 55798
rect 50176 55998 50246 56430
rect 50914 55998 50984 56430
rect 50176 55366 50246 55798
rect 50914 55366 50984 55798
rect 59376 55998 59446 56430
rect 60114 55998 60184 56430
rect 59376 55366 59446 55798
rect 60114 55366 60184 55798
rect 68576 55998 68646 56430
rect 69314 55998 69384 56430
rect 68576 55366 68646 55798
rect 69314 55366 69384 55798
rect 4176 46118 4246 46550
rect 4914 46118 4984 46550
rect 4176 45486 4246 45918
rect 4914 45486 4984 45918
rect 13376 46118 13446 46550
rect 14114 46118 14184 46550
rect 13376 45486 13446 45918
rect 14114 45486 14184 45918
rect 22576 46118 22646 46550
rect 23314 46118 23384 46550
rect 22576 45486 22646 45918
rect 23314 45486 23384 45918
rect 31776 46118 31846 46550
rect 32514 46118 32584 46550
rect 31776 45486 31846 45918
rect 32514 45486 32584 45918
rect 40976 46118 41046 46550
rect 41714 46118 41784 46550
rect 40976 45486 41046 45918
rect 41714 45486 41784 45918
rect 50176 46118 50246 46550
rect 50914 46118 50984 46550
rect 50176 45486 50246 45918
rect 50914 45486 50984 45918
rect 59376 46118 59446 46550
rect 60114 46118 60184 46550
rect 59376 45486 59446 45918
rect 60114 45486 60184 45918
rect 68576 46118 68646 46550
rect 69314 46118 69384 46550
rect 68576 45486 68646 45918
rect 69314 45486 69384 45918
rect 4176 36238 4246 36670
rect 4914 36238 4984 36670
rect 4176 35606 4246 36038
rect 4914 35606 4984 36038
rect 13376 36238 13446 36670
rect 14114 36238 14184 36670
rect 13376 35606 13446 36038
rect 14114 35606 14184 36038
rect 22576 36238 22646 36670
rect 23314 36238 23384 36670
rect 22576 35606 22646 36038
rect 23314 35606 23384 36038
rect 31776 36238 31846 36670
rect 32514 36238 32584 36670
rect 31776 35606 31846 36038
rect 32514 35606 32584 36038
rect 40976 36238 41046 36670
rect 41714 36238 41784 36670
rect 40976 35606 41046 36038
rect 41714 35606 41784 36038
rect 50176 36238 50246 36670
rect 50914 36238 50984 36670
rect 50176 35606 50246 36038
rect 50914 35606 50984 36038
rect 59376 36238 59446 36670
rect 60114 36238 60184 36670
rect 59376 35606 59446 36038
rect 60114 35606 60184 36038
rect 68576 36238 68646 36670
rect 69314 36238 69384 36670
rect 68576 35606 68646 36038
rect 69314 35606 69384 36038
rect 4176 26358 4246 26790
rect 4914 26358 4984 26790
rect 4176 25726 4246 26158
rect 4914 25726 4984 26158
rect 13376 26358 13446 26790
rect 14114 26358 14184 26790
rect 13376 25726 13446 26158
rect 14114 25726 14184 26158
rect 22576 26358 22646 26790
rect 23314 26358 23384 26790
rect 22576 25726 22646 26158
rect 23314 25726 23384 26158
rect 31776 26358 31846 26790
rect 32514 26358 32584 26790
rect 31776 25726 31846 26158
rect 32514 25726 32584 26158
rect 40976 26358 41046 26790
rect 41714 26358 41784 26790
rect 40976 25726 41046 26158
rect 41714 25726 41784 26158
rect 50176 26358 50246 26790
rect 50914 26358 50984 26790
rect 50176 25726 50246 26158
rect 50914 25726 50984 26158
rect 59376 26358 59446 26790
rect 60114 26358 60184 26790
rect 59376 25726 59446 26158
rect 60114 25726 60184 26158
rect 68576 26358 68646 26790
rect 69314 26358 69384 26790
rect 68576 25726 68646 26158
rect 69314 25726 69384 26158
rect 4176 16478 4246 16910
rect 4914 16478 4984 16910
rect 4176 15846 4246 16278
rect 4914 15846 4984 16278
rect 13376 16478 13446 16910
rect 14114 16478 14184 16910
rect 13376 15846 13446 16278
rect 14114 15846 14184 16278
rect 22576 16478 22646 16910
rect 23314 16478 23384 16910
rect 22576 15846 22646 16278
rect 23314 15846 23384 16278
rect 31776 16478 31846 16910
rect 32514 16478 32584 16910
rect 31776 15846 31846 16278
rect 32514 15846 32584 16278
rect 40976 16478 41046 16910
rect 41714 16478 41784 16910
rect 40976 15846 41046 16278
rect 41714 15846 41784 16278
rect 50176 16478 50246 16910
rect 50914 16478 50984 16910
rect 50176 15846 50246 16278
rect 50914 15846 50984 16278
rect 59376 16478 59446 16910
rect 60114 16478 60184 16910
rect 59376 15846 59446 16278
rect 60114 15846 60184 16278
rect 68576 16478 68646 16910
rect 69314 16478 69384 16910
rect 68576 15846 68646 16278
rect 69314 15846 69384 16278
rect 4176 6598 4246 7030
rect 4914 6598 4984 7030
rect 4176 5966 4246 6398
rect 4914 5966 4984 6398
rect 13376 6598 13446 7030
rect 14114 6598 14184 7030
rect 13376 5966 13446 6398
rect 14114 5966 14184 6398
rect 22576 6598 22646 7030
rect 23314 6598 23384 7030
rect 22576 5966 22646 6398
rect 23314 5966 23384 6398
rect 31776 6598 31846 7030
rect 32514 6598 32584 7030
rect 31776 5966 31846 6398
rect 32514 5966 32584 6398
rect 40976 6598 41046 7030
rect 41714 6598 41784 7030
rect 40976 5966 41046 6398
rect 41714 5966 41784 6398
rect 50176 6598 50246 7030
rect 50914 6598 50984 7030
rect 50176 5966 50246 6398
rect 50914 5966 50984 6398
rect 59376 6598 59446 7030
rect 60114 6598 60184 7030
rect 59376 5966 59446 6398
rect 60114 5966 60184 6398
rect 68576 6598 68646 7030
rect 69314 6598 69384 7030
rect 68576 5966 68646 6398
rect 69314 5966 69384 6398
<< xpolyres >>
rect 4176 95318 4246 95518
rect 4914 95318 4984 95518
rect 4176 85438 4246 85638
rect 4914 85438 4984 85638
rect 13376 85438 13446 85638
rect 14114 85438 14184 85638
rect 4176 75558 4246 75758
rect 4914 75558 4984 75758
rect 13376 75558 13446 75758
rect 14114 75558 14184 75758
rect 22576 75558 22646 75758
rect 23314 75558 23384 75758
rect 31776 75558 31846 75758
rect 32514 75558 32584 75758
rect 4176 65678 4246 65878
rect 4914 65678 4984 65878
rect 13376 65678 13446 65878
rect 14114 65678 14184 65878
rect 22576 65678 22646 65878
rect 23314 65678 23384 65878
rect 31776 65678 31846 65878
rect 32514 65678 32584 65878
rect 40976 65678 41046 65878
rect 41714 65678 41784 65878
rect 50176 65678 50246 65878
rect 50914 65678 50984 65878
rect 59376 65678 59446 65878
rect 60114 65678 60184 65878
rect 68576 65678 68646 65878
rect 69314 65678 69384 65878
rect 4176 55798 4246 55998
rect 4914 55798 4984 55998
rect 13376 55798 13446 55998
rect 14114 55798 14184 55998
rect 22576 55798 22646 55998
rect 23314 55798 23384 55998
rect 31776 55798 31846 55998
rect 32514 55798 32584 55998
rect 40976 55798 41046 55998
rect 41714 55798 41784 55998
rect 50176 55798 50246 55998
rect 50914 55798 50984 55998
rect 59376 55798 59446 55998
rect 60114 55798 60184 55998
rect 68576 55798 68646 55998
rect 69314 55798 69384 55998
rect 4176 45918 4246 46118
rect 4914 45918 4984 46118
rect 13376 45918 13446 46118
rect 14114 45918 14184 46118
rect 22576 45918 22646 46118
rect 23314 45918 23384 46118
rect 31776 45918 31846 46118
rect 32514 45918 32584 46118
rect 40976 45918 41046 46118
rect 41714 45918 41784 46118
rect 50176 45918 50246 46118
rect 50914 45918 50984 46118
rect 59376 45918 59446 46118
rect 60114 45918 60184 46118
rect 68576 45918 68646 46118
rect 69314 45918 69384 46118
rect 4176 36038 4246 36238
rect 4914 36038 4984 36238
rect 13376 36038 13446 36238
rect 14114 36038 14184 36238
rect 22576 36038 22646 36238
rect 23314 36038 23384 36238
rect 31776 36038 31846 36238
rect 32514 36038 32584 36238
rect 40976 36038 41046 36238
rect 41714 36038 41784 36238
rect 50176 36038 50246 36238
rect 50914 36038 50984 36238
rect 59376 36038 59446 36238
rect 60114 36038 60184 36238
rect 68576 36038 68646 36238
rect 69314 36038 69384 36238
rect 4176 26158 4246 26358
rect 4914 26158 4984 26358
rect 13376 26158 13446 26358
rect 14114 26158 14184 26358
rect 22576 26158 22646 26358
rect 23314 26158 23384 26358
rect 31776 26158 31846 26358
rect 32514 26158 32584 26358
rect 40976 26158 41046 26358
rect 41714 26158 41784 26358
rect 50176 26158 50246 26358
rect 50914 26158 50984 26358
rect 59376 26158 59446 26358
rect 60114 26158 60184 26358
rect 68576 26158 68646 26358
rect 69314 26158 69384 26358
rect 4176 16278 4246 16478
rect 4914 16278 4984 16478
rect 13376 16278 13446 16478
rect 14114 16278 14184 16478
rect 22576 16278 22646 16478
rect 23314 16278 23384 16478
rect 31776 16278 31846 16478
rect 32514 16278 32584 16478
rect 40976 16278 41046 16478
rect 41714 16278 41784 16478
rect 50176 16278 50246 16478
rect 50914 16278 50984 16478
rect 59376 16278 59446 16478
rect 60114 16278 60184 16478
rect 68576 16278 68646 16478
rect 69314 16278 69384 16478
rect 4176 6398 4246 6598
rect 4914 6398 4984 6598
rect 13376 6398 13446 6598
rect 14114 6398 14184 6598
rect 22576 6398 22646 6598
rect 23314 6398 23384 6598
rect 31776 6398 31846 6598
rect 32514 6398 32584 6598
rect 40976 6398 41046 6598
rect 41714 6398 41784 6598
rect 50176 6398 50246 6598
rect 50914 6398 50984 6598
rect 59376 6398 59446 6598
rect 60114 6398 60184 6598
rect 68576 6398 68646 6598
rect 69314 6398 69384 6598
<< locali >>
rect -506 95532 -218 95560
rect -506 95530 -440 95532
rect -392 95530 -326 95532
rect -278 95530 -218 95532
rect -506 95490 -480 95530
rect -360 95494 -326 95530
rect -440 95490 -400 95494
rect -360 95490 -310 95494
rect -270 95490 -218 95530
rect -506 95458 -218 95490
rect -424 95384 -390 95400
rect -610 94760 -550 94770
rect -610 94720 -600 94760
rect -560 94750 -550 94760
rect -424 94752 -390 94808
rect -336 95384 -302 95458
rect 4479 95330 4491 95364
rect 4529 95330 4563 95364
rect 4597 95330 4631 95364
rect 4669 95330 4681 95364
rect 4477 95280 4511 95296
rect 4366 95252 4400 95262
rect 4366 95180 4400 95212
rect 4366 95110 4400 95144
rect 4366 95042 4400 95074
rect 4366 94992 4400 95002
rect 4477 95212 4511 95218
rect 4477 95144 4511 95146
rect 4477 95108 4511 95110
rect 4477 95036 4511 95042
rect 4477 94958 4511 94974
rect 4563 95280 4597 95296
rect 4563 95212 4597 95218
rect 4563 95144 4597 95146
rect 4563 95108 4597 95110
rect 4563 95036 4597 95042
rect 4563 94958 4597 94974
rect 4649 95280 4683 95296
rect 4649 95212 4683 95218
rect 4649 95144 4683 95146
rect 4649 95108 4683 95110
rect 4649 95036 4683 95042
rect 4760 95252 4794 95262
rect 4760 95180 4794 95212
rect 4760 95110 4794 95144
rect 4760 95042 4794 95074
rect 4760 94992 4794 95002
rect 4649 94958 4683 94974
rect 4479 94890 4491 94924
rect 4529 94890 4563 94924
rect 4597 94890 4631 94924
rect 4669 94890 4681 94924
rect -336 94792 -302 94808
rect -508 94750 -390 94752
rect -560 94720 -390 94750
rect -610 94712 -390 94720
rect -610 94710 -490 94712
rect -424 94654 -390 94712
rect -240 94740 -160 94760
rect -240 94700 -220 94740
rect -180 94700 -160 94740
rect -240 94680 -160 94700
rect -424 94362 -390 94378
rect -336 94654 -302 94670
rect -336 94298 -302 94378
rect -506 94290 -218 94298
rect -506 94240 -440 94290
rect -390 94276 -330 94290
rect -390 94240 -338 94276
rect -280 94240 -218 94290
rect -506 94220 -218 94240
rect -506 85652 -218 85680
rect -506 85650 -440 85652
rect -392 85650 -326 85652
rect -278 85650 -218 85652
rect -506 85610 -480 85650
rect -360 85614 -326 85650
rect -440 85610 -400 85614
rect -360 85610 -310 85614
rect -270 85610 -218 85650
rect -506 85578 -218 85610
rect -424 85504 -390 85520
rect -610 84880 -550 84890
rect -610 84840 -600 84880
rect -560 84870 -550 84880
rect -424 84872 -390 84928
rect -336 85504 -302 85578
rect 4479 85450 4491 85484
rect 4529 85450 4563 85484
rect 4597 85450 4631 85484
rect 4669 85450 4681 85484
rect 13679 85450 13691 85484
rect 13729 85450 13763 85484
rect 13797 85450 13831 85484
rect 13869 85450 13881 85484
rect 4477 85400 4511 85416
rect 4366 85372 4400 85382
rect 4366 85300 4400 85332
rect 4366 85230 4400 85264
rect 4366 85162 4400 85194
rect 4366 85112 4400 85122
rect 4477 85332 4511 85338
rect 4477 85264 4511 85266
rect 4477 85228 4511 85230
rect 4477 85156 4511 85162
rect 4477 85078 4511 85094
rect 4563 85400 4597 85416
rect 4563 85332 4597 85338
rect 4563 85264 4597 85266
rect 4563 85228 4597 85230
rect 4563 85156 4597 85162
rect 4563 85078 4597 85094
rect 4649 85400 4683 85416
rect 4649 85332 4683 85338
rect 4649 85264 4683 85266
rect 4649 85228 4683 85230
rect 4649 85156 4683 85162
rect 4760 85372 4794 85382
rect 4760 85300 4794 85332
rect 4760 85230 4794 85264
rect 4760 85162 4794 85194
rect 4760 85112 4794 85122
rect 4649 85078 4683 85094
rect 4479 85010 4491 85044
rect 4529 85010 4563 85044
rect 4597 85010 4631 85044
rect 4669 85010 4681 85044
rect 13677 85400 13711 85416
rect 13566 85372 13600 85382
rect 13566 85300 13600 85332
rect 13566 85230 13600 85264
rect 13566 85162 13600 85194
rect 13566 85112 13600 85122
rect 13677 85332 13711 85338
rect 13677 85264 13711 85266
rect 13677 85228 13711 85230
rect 13677 85156 13711 85162
rect 13677 85078 13711 85094
rect 13763 85400 13797 85416
rect 13763 85332 13797 85338
rect 13763 85264 13797 85266
rect 13763 85228 13797 85230
rect 13763 85156 13797 85162
rect 13763 85078 13797 85094
rect 13849 85400 13883 85416
rect 13849 85332 13883 85338
rect 13849 85264 13883 85266
rect 13849 85228 13883 85230
rect 13849 85156 13883 85162
rect 13960 85372 13994 85382
rect 13960 85300 13994 85332
rect 13960 85230 13994 85264
rect 13960 85162 13994 85194
rect 13960 85112 13994 85122
rect 13849 85078 13883 85094
rect 13679 85010 13691 85044
rect 13729 85010 13763 85044
rect 13797 85010 13831 85044
rect 13869 85010 13881 85044
rect -336 84912 -302 84928
rect -508 84870 -390 84872
rect -560 84840 -390 84870
rect -610 84832 -390 84840
rect -610 84830 -490 84832
rect -424 84774 -390 84832
rect -240 84860 -160 84880
rect -240 84820 -220 84860
rect -180 84820 -160 84860
rect -240 84800 -160 84820
rect -424 84482 -390 84498
rect -336 84774 -302 84790
rect -336 84418 -302 84498
rect -506 84410 -218 84418
rect -506 84360 -440 84410
rect -390 84396 -330 84410
rect -390 84360 -338 84396
rect -280 84360 -218 84410
rect -506 84340 -218 84360
rect -506 75772 -218 75800
rect -506 75770 -440 75772
rect -392 75770 -326 75772
rect -278 75770 -218 75772
rect -506 75730 -480 75770
rect -360 75734 -326 75770
rect -440 75730 -400 75734
rect -360 75730 -310 75734
rect -270 75730 -218 75770
rect -506 75698 -218 75730
rect -424 75624 -390 75640
rect -610 75000 -550 75010
rect -610 74960 -600 75000
rect -560 74990 -550 75000
rect -424 74992 -390 75048
rect -336 75624 -302 75698
rect 4479 75570 4491 75604
rect 4529 75570 4563 75604
rect 4597 75570 4631 75604
rect 4669 75570 4681 75604
rect 13679 75570 13691 75604
rect 13729 75570 13763 75604
rect 13797 75570 13831 75604
rect 13869 75570 13881 75604
rect 22879 75570 22891 75604
rect 22929 75570 22963 75604
rect 22997 75570 23031 75604
rect 23069 75570 23081 75604
rect 32079 75570 32091 75604
rect 32129 75570 32163 75604
rect 32197 75570 32231 75604
rect 32269 75570 32281 75604
rect 4477 75520 4511 75536
rect 4366 75492 4400 75502
rect 4366 75420 4400 75452
rect 4366 75350 4400 75384
rect 4366 75282 4400 75314
rect 4366 75232 4400 75242
rect 4477 75452 4511 75458
rect 4477 75384 4511 75386
rect 4477 75348 4511 75350
rect 4477 75276 4511 75282
rect 4477 75198 4511 75214
rect 4563 75520 4597 75536
rect 4563 75452 4597 75458
rect 4563 75384 4597 75386
rect 4563 75348 4597 75350
rect 4563 75276 4597 75282
rect 4563 75198 4597 75214
rect 4649 75520 4683 75536
rect 4649 75452 4683 75458
rect 4649 75384 4683 75386
rect 4649 75348 4683 75350
rect 4649 75276 4683 75282
rect 4760 75492 4794 75502
rect 4760 75420 4794 75452
rect 4760 75350 4794 75384
rect 4760 75282 4794 75314
rect 4760 75232 4794 75242
rect 4649 75198 4683 75214
rect 4479 75130 4491 75164
rect 4529 75130 4563 75164
rect 4597 75130 4631 75164
rect 4669 75130 4681 75164
rect 13677 75520 13711 75536
rect 13566 75492 13600 75502
rect 13566 75420 13600 75452
rect 13566 75350 13600 75384
rect 13566 75282 13600 75314
rect 13566 75232 13600 75242
rect 13677 75452 13711 75458
rect 13677 75384 13711 75386
rect 13677 75348 13711 75350
rect 13677 75276 13711 75282
rect 13677 75198 13711 75214
rect 13763 75520 13797 75536
rect 13763 75452 13797 75458
rect 13763 75384 13797 75386
rect 13763 75348 13797 75350
rect 13763 75276 13797 75282
rect 13763 75198 13797 75214
rect 13849 75520 13883 75536
rect 13849 75452 13883 75458
rect 13849 75384 13883 75386
rect 13849 75348 13883 75350
rect 13849 75276 13883 75282
rect 13960 75492 13994 75502
rect 13960 75420 13994 75452
rect 13960 75350 13994 75384
rect 13960 75282 13994 75314
rect 13960 75232 13994 75242
rect 13849 75198 13883 75214
rect 13679 75130 13691 75164
rect 13729 75130 13763 75164
rect 13797 75130 13831 75164
rect 13869 75130 13881 75164
rect 22877 75520 22911 75536
rect 22766 75492 22800 75502
rect 22766 75420 22800 75452
rect 22766 75350 22800 75384
rect 22766 75282 22800 75314
rect 22766 75232 22800 75242
rect 22877 75452 22911 75458
rect 22877 75384 22911 75386
rect 22877 75348 22911 75350
rect 22877 75276 22911 75282
rect 22877 75198 22911 75214
rect 22963 75520 22997 75536
rect 22963 75452 22997 75458
rect 22963 75384 22997 75386
rect 22963 75348 22997 75350
rect 22963 75276 22997 75282
rect 22963 75198 22997 75214
rect 23049 75520 23083 75536
rect 23049 75452 23083 75458
rect 23049 75384 23083 75386
rect 23049 75348 23083 75350
rect 23049 75276 23083 75282
rect 23160 75492 23194 75502
rect 23160 75420 23194 75452
rect 23160 75350 23194 75384
rect 23160 75282 23194 75314
rect 23160 75232 23194 75242
rect 23049 75198 23083 75214
rect 22879 75130 22891 75164
rect 22929 75130 22963 75164
rect 22997 75130 23031 75164
rect 23069 75130 23081 75164
rect 32077 75520 32111 75536
rect 31966 75492 32000 75502
rect 31966 75420 32000 75452
rect 31966 75350 32000 75384
rect 31966 75282 32000 75314
rect 31966 75232 32000 75242
rect 32077 75452 32111 75458
rect 32077 75384 32111 75386
rect 32077 75348 32111 75350
rect 32077 75276 32111 75282
rect 32077 75198 32111 75214
rect 32163 75520 32197 75536
rect 32163 75452 32197 75458
rect 32163 75384 32197 75386
rect 32163 75348 32197 75350
rect 32163 75276 32197 75282
rect 32163 75198 32197 75214
rect 32249 75520 32283 75536
rect 32249 75452 32283 75458
rect 32249 75384 32283 75386
rect 32249 75348 32283 75350
rect 32249 75276 32283 75282
rect 32360 75492 32394 75502
rect 32360 75420 32394 75452
rect 32360 75350 32394 75384
rect 32360 75282 32394 75314
rect 32360 75232 32394 75242
rect 32249 75198 32283 75214
rect 32079 75130 32091 75164
rect 32129 75130 32163 75164
rect 32197 75130 32231 75164
rect 32269 75130 32281 75164
rect -336 75032 -302 75048
rect -508 74990 -390 74992
rect -560 74960 -390 74990
rect -610 74952 -390 74960
rect -610 74950 -490 74952
rect -424 74894 -390 74952
rect -240 74980 -160 75000
rect -240 74940 -220 74980
rect -180 74940 -160 74980
rect -240 74920 -160 74940
rect -424 74602 -390 74618
rect -336 74894 -302 74910
rect -336 74538 -302 74618
rect -506 74530 -218 74538
rect -506 74480 -440 74530
rect -390 74516 -330 74530
rect -390 74480 -338 74516
rect -280 74480 -218 74530
rect -506 74460 -218 74480
rect -506 65892 -218 65920
rect -506 65890 -440 65892
rect -392 65890 -326 65892
rect -278 65890 -218 65892
rect -506 65850 -480 65890
rect -360 65854 -326 65890
rect -440 65850 -400 65854
rect -360 65850 -310 65854
rect -270 65850 -218 65890
rect -506 65818 -218 65850
rect -424 65744 -390 65760
rect -610 65120 -550 65130
rect -610 65080 -600 65120
rect -560 65110 -550 65120
rect -424 65112 -390 65168
rect -336 65744 -302 65818
rect 4479 65690 4491 65724
rect 4529 65690 4563 65724
rect 4597 65690 4631 65724
rect 4669 65690 4681 65724
rect 13679 65690 13691 65724
rect 13729 65690 13763 65724
rect 13797 65690 13831 65724
rect 13869 65690 13881 65724
rect 22879 65690 22891 65724
rect 22929 65690 22963 65724
rect 22997 65690 23031 65724
rect 23069 65690 23081 65724
rect 32079 65690 32091 65724
rect 32129 65690 32163 65724
rect 32197 65690 32231 65724
rect 32269 65690 32281 65724
rect 41279 65690 41291 65724
rect 41329 65690 41363 65724
rect 41397 65690 41431 65724
rect 41469 65690 41481 65724
rect 50479 65690 50491 65724
rect 50529 65690 50563 65724
rect 50597 65690 50631 65724
rect 50669 65690 50681 65724
rect 59679 65690 59691 65724
rect 59729 65690 59763 65724
rect 59797 65690 59831 65724
rect 59869 65690 59881 65724
rect 68879 65690 68891 65724
rect 68929 65690 68963 65724
rect 68997 65690 69031 65724
rect 69069 65690 69081 65724
rect 4477 65640 4511 65656
rect 4366 65612 4400 65622
rect 4366 65540 4400 65572
rect 4366 65470 4400 65504
rect 4366 65402 4400 65434
rect 4366 65352 4400 65362
rect 4477 65572 4511 65578
rect 4477 65504 4511 65506
rect 4477 65468 4511 65470
rect 4477 65396 4511 65402
rect 4477 65318 4511 65334
rect 4563 65640 4597 65656
rect 4563 65572 4597 65578
rect 4563 65504 4597 65506
rect 4563 65468 4597 65470
rect 4563 65396 4597 65402
rect 4563 65318 4597 65334
rect 4649 65640 4683 65656
rect 4649 65572 4683 65578
rect 4649 65504 4683 65506
rect 4649 65468 4683 65470
rect 4649 65396 4683 65402
rect 4760 65612 4794 65622
rect 4760 65540 4794 65572
rect 4760 65470 4794 65504
rect 4760 65402 4794 65434
rect 4760 65352 4794 65362
rect 4649 65318 4683 65334
rect 4479 65250 4491 65284
rect 4529 65250 4563 65284
rect 4597 65250 4631 65284
rect 4669 65250 4681 65284
rect 13677 65640 13711 65656
rect 13566 65612 13600 65622
rect 13566 65540 13600 65572
rect 13566 65470 13600 65504
rect 13566 65402 13600 65434
rect 13566 65352 13600 65362
rect 13677 65572 13711 65578
rect 13677 65504 13711 65506
rect 13677 65468 13711 65470
rect 13677 65396 13711 65402
rect 13677 65318 13711 65334
rect 13763 65640 13797 65656
rect 13763 65572 13797 65578
rect 13763 65504 13797 65506
rect 13763 65468 13797 65470
rect 13763 65396 13797 65402
rect 13763 65318 13797 65334
rect 13849 65640 13883 65656
rect 13849 65572 13883 65578
rect 13849 65504 13883 65506
rect 13849 65468 13883 65470
rect 13849 65396 13883 65402
rect 13960 65612 13994 65622
rect 13960 65540 13994 65572
rect 13960 65470 13994 65504
rect 13960 65402 13994 65434
rect 13960 65352 13994 65362
rect 13849 65318 13883 65334
rect 13679 65250 13691 65284
rect 13729 65250 13763 65284
rect 13797 65250 13831 65284
rect 13869 65250 13881 65284
rect 22877 65640 22911 65656
rect 22766 65612 22800 65622
rect 22766 65540 22800 65572
rect 22766 65470 22800 65504
rect 22766 65402 22800 65434
rect 22766 65352 22800 65362
rect 22877 65572 22911 65578
rect 22877 65504 22911 65506
rect 22877 65468 22911 65470
rect 22877 65396 22911 65402
rect 22877 65318 22911 65334
rect 22963 65640 22997 65656
rect 22963 65572 22997 65578
rect 22963 65504 22997 65506
rect 22963 65468 22997 65470
rect 22963 65396 22997 65402
rect 22963 65318 22997 65334
rect 23049 65640 23083 65656
rect 23049 65572 23083 65578
rect 23049 65504 23083 65506
rect 23049 65468 23083 65470
rect 23049 65396 23083 65402
rect 23160 65612 23194 65622
rect 23160 65540 23194 65572
rect 23160 65470 23194 65504
rect 23160 65402 23194 65434
rect 23160 65352 23194 65362
rect 23049 65318 23083 65334
rect 22879 65250 22891 65284
rect 22929 65250 22963 65284
rect 22997 65250 23031 65284
rect 23069 65250 23081 65284
rect 32077 65640 32111 65656
rect 31966 65612 32000 65622
rect 31966 65540 32000 65572
rect 31966 65470 32000 65504
rect 31966 65402 32000 65434
rect 31966 65352 32000 65362
rect 32077 65572 32111 65578
rect 32077 65504 32111 65506
rect 32077 65468 32111 65470
rect 32077 65396 32111 65402
rect 32077 65318 32111 65334
rect 32163 65640 32197 65656
rect 32163 65572 32197 65578
rect 32163 65504 32197 65506
rect 32163 65468 32197 65470
rect 32163 65396 32197 65402
rect 32163 65318 32197 65334
rect 32249 65640 32283 65656
rect 32249 65572 32283 65578
rect 32249 65504 32283 65506
rect 32249 65468 32283 65470
rect 32249 65396 32283 65402
rect 32360 65612 32394 65622
rect 32360 65540 32394 65572
rect 32360 65470 32394 65504
rect 32360 65402 32394 65434
rect 32360 65352 32394 65362
rect 32249 65318 32283 65334
rect 32079 65250 32091 65284
rect 32129 65250 32163 65284
rect 32197 65250 32231 65284
rect 32269 65250 32281 65284
rect 41277 65640 41311 65656
rect 41166 65612 41200 65622
rect 41166 65540 41200 65572
rect 41166 65470 41200 65504
rect 41166 65402 41200 65434
rect 41166 65352 41200 65362
rect 41277 65572 41311 65578
rect 41277 65504 41311 65506
rect 41277 65468 41311 65470
rect 41277 65396 41311 65402
rect 41277 65318 41311 65334
rect 41363 65640 41397 65656
rect 41363 65572 41397 65578
rect 41363 65504 41397 65506
rect 41363 65468 41397 65470
rect 41363 65396 41397 65402
rect 41363 65318 41397 65334
rect 41449 65640 41483 65656
rect 41449 65572 41483 65578
rect 41449 65504 41483 65506
rect 41449 65468 41483 65470
rect 41449 65396 41483 65402
rect 41560 65612 41594 65622
rect 41560 65540 41594 65572
rect 41560 65470 41594 65504
rect 41560 65402 41594 65434
rect 41560 65352 41594 65362
rect 41449 65318 41483 65334
rect 41279 65250 41291 65284
rect 41329 65250 41363 65284
rect 41397 65250 41431 65284
rect 41469 65250 41481 65284
rect 50477 65640 50511 65656
rect 50366 65612 50400 65622
rect 50366 65540 50400 65572
rect 50366 65470 50400 65504
rect 50366 65402 50400 65434
rect 50366 65352 50400 65362
rect 50477 65572 50511 65578
rect 50477 65504 50511 65506
rect 50477 65468 50511 65470
rect 50477 65396 50511 65402
rect 50477 65318 50511 65334
rect 50563 65640 50597 65656
rect 50563 65572 50597 65578
rect 50563 65504 50597 65506
rect 50563 65468 50597 65470
rect 50563 65396 50597 65402
rect 50563 65318 50597 65334
rect 50649 65640 50683 65656
rect 50649 65572 50683 65578
rect 50649 65504 50683 65506
rect 50649 65468 50683 65470
rect 50649 65396 50683 65402
rect 50760 65612 50794 65622
rect 50760 65540 50794 65572
rect 50760 65470 50794 65504
rect 50760 65402 50794 65434
rect 50760 65352 50794 65362
rect 50649 65318 50683 65334
rect 50479 65250 50491 65284
rect 50529 65250 50563 65284
rect 50597 65250 50631 65284
rect 50669 65250 50681 65284
rect 59677 65640 59711 65656
rect 59566 65612 59600 65622
rect 59566 65540 59600 65572
rect 59566 65470 59600 65504
rect 59566 65402 59600 65434
rect 59566 65352 59600 65362
rect 59677 65572 59711 65578
rect 59677 65504 59711 65506
rect 59677 65468 59711 65470
rect 59677 65396 59711 65402
rect 59677 65318 59711 65334
rect 59763 65640 59797 65656
rect 59763 65572 59797 65578
rect 59763 65504 59797 65506
rect 59763 65468 59797 65470
rect 59763 65396 59797 65402
rect 59763 65318 59797 65334
rect 59849 65640 59883 65656
rect 59849 65572 59883 65578
rect 59849 65504 59883 65506
rect 59849 65468 59883 65470
rect 59849 65396 59883 65402
rect 59960 65612 59994 65622
rect 59960 65540 59994 65572
rect 59960 65470 59994 65504
rect 59960 65402 59994 65434
rect 59960 65352 59994 65362
rect 59849 65318 59883 65334
rect 59679 65250 59691 65284
rect 59729 65250 59763 65284
rect 59797 65250 59831 65284
rect 59869 65250 59881 65284
rect 68877 65640 68911 65656
rect 68766 65612 68800 65622
rect 68766 65540 68800 65572
rect 68766 65470 68800 65504
rect 68766 65402 68800 65434
rect 68766 65352 68800 65362
rect 68877 65572 68911 65578
rect 68877 65504 68911 65506
rect 68877 65468 68911 65470
rect 68877 65396 68911 65402
rect 68877 65318 68911 65334
rect 68963 65640 68997 65656
rect 68963 65572 68997 65578
rect 68963 65504 68997 65506
rect 68963 65468 68997 65470
rect 68963 65396 68997 65402
rect 68963 65318 68997 65334
rect 69049 65640 69083 65656
rect 69049 65572 69083 65578
rect 69049 65504 69083 65506
rect 69049 65468 69083 65470
rect 69049 65396 69083 65402
rect 69160 65612 69194 65622
rect 69160 65540 69194 65572
rect 69160 65470 69194 65504
rect 69160 65402 69194 65434
rect 69160 65352 69194 65362
rect 69049 65318 69083 65334
rect 68879 65250 68891 65284
rect 68929 65250 68963 65284
rect 68997 65250 69031 65284
rect 69069 65250 69081 65284
rect -336 65152 -302 65168
rect -508 65110 -390 65112
rect -560 65080 -390 65110
rect -610 65072 -390 65080
rect -610 65070 -490 65072
rect -424 65014 -390 65072
rect -240 65100 -160 65120
rect -240 65060 -220 65100
rect -180 65060 -160 65100
rect -240 65040 -160 65060
rect -424 64722 -390 64738
rect -336 65014 -302 65030
rect -336 64658 -302 64738
rect -506 64650 -218 64658
rect -506 64600 -440 64650
rect -390 64636 -330 64650
rect -390 64600 -338 64636
rect -280 64600 -218 64650
rect -506 64580 -218 64600
rect 4479 55810 4491 55844
rect 4529 55810 4563 55844
rect 4597 55810 4631 55844
rect 4669 55810 4681 55844
rect 13679 55810 13691 55844
rect 13729 55810 13763 55844
rect 13797 55810 13831 55844
rect 13869 55810 13881 55844
rect 22879 55810 22891 55844
rect 22929 55810 22963 55844
rect 22997 55810 23031 55844
rect 23069 55810 23081 55844
rect 32079 55810 32091 55844
rect 32129 55810 32163 55844
rect 32197 55810 32231 55844
rect 32269 55810 32281 55844
rect 41279 55810 41291 55844
rect 41329 55810 41363 55844
rect 41397 55810 41431 55844
rect 41469 55810 41481 55844
rect 50479 55810 50491 55844
rect 50529 55810 50563 55844
rect 50597 55810 50631 55844
rect 50669 55810 50681 55844
rect 59679 55810 59691 55844
rect 59729 55810 59763 55844
rect 59797 55810 59831 55844
rect 59869 55810 59881 55844
rect 68879 55810 68891 55844
rect 68929 55810 68963 55844
rect 68997 55810 69031 55844
rect 69069 55810 69081 55844
rect 4477 55760 4511 55776
rect 4366 55732 4400 55742
rect 4366 55660 4400 55692
rect 4366 55590 4400 55624
rect 4366 55522 4400 55554
rect 4366 55472 4400 55482
rect 4477 55692 4511 55698
rect 4477 55624 4511 55626
rect 4477 55588 4511 55590
rect 4477 55516 4511 55522
rect 4477 55438 4511 55454
rect 4563 55760 4597 55776
rect 4563 55692 4597 55698
rect 4563 55624 4597 55626
rect 4563 55588 4597 55590
rect 4563 55516 4597 55522
rect 4563 55438 4597 55454
rect 4649 55760 4683 55776
rect 4649 55692 4683 55698
rect 4649 55624 4683 55626
rect 4649 55588 4683 55590
rect 4649 55516 4683 55522
rect 4760 55732 4794 55742
rect 4760 55660 4794 55692
rect 4760 55590 4794 55624
rect 4760 55522 4794 55554
rect 4760 55472 4794 55482
rect 4649 55438 4683 55454
rect 4479 55370 4491 55404
rect 4529 55370 4563 55404
rect 4597 55370 4631 55404
rect 4669 55370 4681 55404
rect 13677 55760 13711 55776
rect 13566 55732 13600 55742
rect 13566 55660 13600 55692
rect 13566 55590 13600 55624
rect 13566 55522 13600 55554
rect 13566 55472 13600 55482
rect 13677 55692 13711 55698
rect 13677 55624 13711 55626
rect 13677 55588 13711 55590
rect 13677 55516 13711 55522
rect 13677 55438 13711 55454
rect 13763 55760 13797 55776
rect 13763 55692 13797 55698
rect 13763 55624 13797 55626
rect 13763 55588 13797 55590
rect 13763 55516 13797 55522
rect 13763 55438 13797 55454
rect 13849 55760 13883 55776
rect 13849 55692 13883 55698
rect 13849 55624 13883 55626
rect 13849 55588 13883 55590
rect 13849 55516 13883 55522
rect 13960 55732 13994 55742
rect 13960 55660 13994 55692
rect 13960 55590 13994 55624
rect 13960 55522 13994 55554
rect 13960 55472 13994 55482
rect 13849 55438 13883 55454
rect 13679 55370 13691 55404
rect 13729 55370 13763 55404
rect 13797 55370 13831 55404
rect 13869 55370 13881 55404
rect 22877 55760 22911 55776
rect 22766 55732 22800 55742
rect 22766 55660 22800 55692
rect 22766 55590 22800 55624
rect 22766 55522 22800 55554
rect 22766 55472 22800 55482
rect 22877 55692 22911 55698
rect 22877 55624 22911 55626
rect 22877 55588 22911 55590
rect 22877 55516 22911 55522
rect 22877 55438 22911 55454
rect 22963 55760 22997 55776
rect 22963 55692 22997 55698
rect 22963 55624 22997 55626
rect 22963 55588 22997 55590
rect 22963 55516 22997 55522
rect 22963 55438 22997 55454
rect 23049 55760 23083 55776
rect 23049 55692 23083 55698
rect 23049 55624 23083 55626
rect 23049 55588 23083 55590
rect 23049 55516 23083 55522
rect 23160 55732 23194 55742
rect 23160 55660 23194 55692
rect 23160 55590 23194 55624
rect 23160 55522 23194 55554
rect 23160 55472 23194 55482
rect 23049 55438 23083 55454
rect 22879 55370 22891 55404
rect 22929 55370 22963 55404
rect 22997 55370 23031 55404
rect 23069 55370 23081 55404
rect 32077 55760 32111 55776
rect 31966 55732 32000 55742
rect 31966 55660 32000 55692
rect 31966 55590 32000 55624
rect 31966 55522 32000 55554
rect 31966 55472 32000 55482
rect 32077 55692 32111 55698
rect 32077 55624 32111 55626
rect 32077 55588 32111 55590
rect 32077 55516 32111 55522
rect 32077 55438 32111 55454
rect 32163 55760 32197 55776
rect 32163 55692 32197 55698
rect 32163 55624 32197 55626
rect 32163 55588 32197 55590
rect 32163 55516 32197 55522
rect 32163 55438 32197 55454
rect 32249 55760 32283 55776
rect 32249 55692 32283 55698
rect 32249 55624 32283 55626
rect 32249 55588 32283 55590
rect 32249 55516 32283 55522
rect 32360 55732 32394 55742
rect 32360 55660 32394 55692
rect 32360 55590 32394 55624
rect 32360 55522 32394 55554
rect 32360 55472 32394 55482
rect 32249 55438 32283 55454
rect 32079 55370 32091 55404
rect 32129 55370 32163 55404
rect 32197 55370 32231 55404
rect 32269 55370 32281 55404
rect 41277 55760 41311 55776
rect 41166 55732 41200 55742
rect 41166 55660 41200 55692
rect 41166 55590 41200 55624
rect 41166 55522 41200 55554
rect 41166 55472 41200 55482
rect 41277 55692 41311 55698
rect 41277 55624 41311 55626
rect 41277 55588 41311 55590
rect 41277 55516 41311 55522
rect 41277 55438 41311 55454
rect 41363 55760 41397 55776
rect 41363 55692 41397 55698
rect 41363 55624 41397 55626
rect 41363 55588 41397 55590
rect 41363 55516 41397 55522
rect 41363 55438 41397 55454
rect 41449 55760 41483 55776
rect 41449 55692 41483 55698
rect 41449 55624 41483 55626
rect 41449 55588 41483 55590
rect 41449 55516 41483 55522
rect 41560 55732 41594 55742
rect 41560 55660 41594 55692
rect 41560 55590 41594 55624
rect 41560 55522 41594 55554
rect 41560 55472 41594 55482
rect 41449 55438 41483 55454
rect 41279 55370 41291 55404
rect 41329 55370 41363 55404
rect 41397 55370 41431 55404
rect 41469 55370 41481 55404
rect 50477 55760 50511 55776
rect 50366 55732 50400 55742
rect 50366 55660 50400 55692
rect 50366 55590 50400 55624
rect 50366 55522 50400 55554
rect 50366 55472 50400 55482
rect 50477 55692 50511 55698
rect 50477 55624 50511 55626
rect 50477 55588 50511 55590
rect 50477 55516 50511 55522
rect 50477 55438 50511 55454
rect 50563 55760 50597 55776
rect 50563 55692 50597 55698
rect 50563 55624 50597 55626
rect 50563 55588 50597 55590
rect 50563 55516 50597 55522
rect 50563 55438 50597 55454
rect 50649 55760 50683 55776
rect 50649 55692 50683 55698
rect 50649 55624 50683 55626
rect 50649 55588 50683 55590
rect 50649 55516 50683 55522
rect 50760 55732 50794 55742
rect 50760 55660 50794 55692
rect 50760 55590 50794 55624
rect 50760 55522 50794 55554
rect 50760 55472 50794 55482
rect 50649 55438 50683 55454
rect 50479 55370 50491 55404
rect 50529 55370 50563 55404
rect 50597 55370 50631 55404
rect 50669 55370 50681 55404
rect 59677 55760 59711 55776
rect 59566 55732 59600 55742
rect 59566 55660 59600 55692
rect 59566 55590 59600 55624
rect 59566 55522 59600 55554
rect 59566 55472 59600 55482
rect 59677 55692 59711 55698
rect 59677 55624 59711 55626
rect 59677 55588 59711 55590
rect 59677 55516 59711 55522
rect 59677 55438 59711 55454
rect 59763 55760 59797 55776
rect 59763 55692 59797 55698
rect 59763 55624 59797 55626
rect 59763 55588 59797 55590
rect 59763 55516 59797 55522
rect 59763 55438 59797 55454
rect 59849 55760 59883 55776
rect 59849 55692 59883 55698
rect 59849 55624 59883 55626
rect 59849 55588 59883 55590
rect 59849 55516 59883 55522
rect 59960 55732 59994 55742
rect 59960 55660 59994 55692
rect 59960 55590 59994 55624
rect 59960 55522 59994 55554
rect 59960 55472 59994 55482
rect 59849 55438 59883 55454
rect 59679 55370 59691 55404
rect 59729 55370 59763 55404
rect 59797 55370 59831 55404
rect 59869 55370 59881 55404
rect 68877 55760 68911 55776
rect 68766 55732 68800 55742
rect 68766 55660 68800 55692
rect 68766 55590 68800 55624
rect 68766 55522 68800 55554
rect 68766 55472 68800 55482
rect 68877 55692 68911 55698
rect 68877 55624 68911 55626
rect 68877 55588 68911 55590
rect 68877 55516 68911 55522
rect 68877 55438 68911 55454
rect 68963 55760 68997 55776
rect 68963 55692 68997 55698
rect 68963 55624 68997 55626
rect 68963 55588 68997 55590
rect 68963 55516 68997 55522
rect 68963 55438 68997 55454
rect 69049 55760 69083 55776
rect 69049 55692 69083 55698
rect 69049 55624 69083 55626
rect 69049 55588 69083 55590
rect 69049 55516 69083 55522
rect 69160 55732 69194 55742
rect 69160 55660 69194 55692
rect 69160 55590 69194 55624
rect 69160 55522 69194 55554
rect 69160 55472 69194 55482
rect 69049 55438 69083 55454
rect 68879 55370 68891 55404
rect 68929 55370 68963 55404
rect 68997 55370 69031 55404
rect 69069 55370 69081 55404
rect -506 46132 -218 46160
rect -506 46130 -440 46132
rect -392 46130 -326 46132
rect -278 46130 -218 46132
rect -506 46090 -480 46130
rect -360 46094 -326 46130
rect -440 46090 -400 46094
rect -360 46090 -310 46094
rect -270 46090 -218 46130
rect -506 46058 -218 46090
rect -424 45984 -390 46000
rect -610 45360 -550 45370
rect -610 45320 -600 45360
rect -560 45350 -550 45360
rect -424 45352 -390 45408
rect -336 45984 -302 46058
rect 4479 45930 4491 45964
rect 4529 45930 4563 45964
rect 4597 45930 4631 45964
rect 4669 45930 4681 45964
rect 13679 45930 13691 45964
rect 13729 45930 13763 45964
rect 13797 45930 13831 45964
rect 13869 45930 13881 45964
rect 22879 45930 22891 45964
rect 22929 45930 22963 45964
rect 22997 45930 23031 45964
rect 23069 45930 23081 45964
rect 32079 45930 32091 45964
rect 32129 45930 32163 45964
rect 32197 45930 32231 45964
rect 32269 45930 32281 45964
rect 41279 45930 41291 45964
rect 41329 45930 41363 45964
rect 41397 45930 41431 45964
rect 41469 45930 41481 45964
rect 50479 45930 50491 45964
rect 50529 45930 50563 45964
rect 50597 45930 50631 45964
rect 50669 45930 50681 45964
rect 59679 45930 59691 45964
rect 59729 45930 59763 45964
rect 59797 45930 59831 45964
rect 59869 45930 59881 45964
rect 68879 45930 68891 45964
rect 68929 45930 68963 45964
rect 68997 45930 69031 45964
rect 69069 45930 69081 45964
rect 4477 45880 4511 45896
rect 4366 45852 4400 45862
rect 4366 45780 4400 45812
rect 4366 45710 4400 45744
rect 4366 45642 4400 45674
rect 4366 45592 4400 45602
rect 4477 45812 4511 45818
rect 4477 45744 4511 45746
rect 4477 45708 4511 45710
rect 4477 45636 4511 45642
rect 4477 45558 4511 45574
rect 4563 45880 4597 45896
rect 4563 45812 4597 45818
rect 4563 45744 4597 45746
rect 4563 45708 4597 45710
rect 4563 45636 4597 45642
rect 4563 45558 4597 45574
rect 4649 45880 4683 45896
rect 4649 45812 4683 45818
rect 4649 45744 4683 45746
rect 4649 45708 4683 45710
rect 4649 45636 4683 45642
rect 4760 45852 4794 45862
rect 4760 45780 4794 45812
rect 4760 45710 4794 45744
rect 4760 45642 4794 45674
rect 4760 45592 4794 45602
rect 4649 45558 4683 45574
rect 4479 45490 4491 45524
rect 4529 45490 4563 45524
rect 4597 45490 4631 45524
rect 4669 45490 4681 45524
rect 13677 45880 13711 45896
rect 13566 45852 13600 45862
rect 13566 45780 13600 45812
rect 13566 45710 13600 45744
rect 13566 45642 13600 45674
rect 13566 45592 13600 45602
rect 13677 45812 13711 45818
rect 13677 45744 13711 45746
rect 13677 45708 13711 45710
rect 13677 45636 13711 45642
rect 13677 45558 13711 45574
rect 13763 45880 13797 45896
rect 13763 45812 13797 45818
rect 13763 45744 13797 45746
rect 13763 45708 13797 45710
rect 13763 45636 13797 45642
rect 13763 45558 13797 45574
rect 13849 45880 13883 45896
rect 13849 45812 13883 45818
rect 13849 45744 13883 45746
rect 13849 45708 13883 45710
rect 13849 45636 13883 45642
rect 13960 45852 13994 45862
rect 13960 45780 13994 45812
rect 13960 45710 13994 45744
rect 13960 45642 13994 45674
rect 13960 45592 13994 45602
rect 13849 45558 13883 45574
rect 13679 45490 13691 45524
rect 13729 45490 13763 45524
rect 13797 45490 13831 45524
rect 13869 45490 13881 45524
rect 22877 45880 22911 45896
rect 22766 45852 22800 45862
rect 22766 45780 22800 45812
rect 22766 45710 22800 45744
rect 22766 45642 22800 45674
rect 22766 45592 22800 45602
rect 22877 45812 22911 45818
rect 22877 45744 22911 45746
rect 22877 45708 22911 45710
rect 22877 45636 22911 45642
rect 22877 45558 22911 45574
rect 22963 45880 22997 45896
rect 22963 45812 22997 45818
rect 22963 45744 22997 45746
rect 22963 45708 22997 45710
rect 22963 45636 22997 45642
rect 22963 45558 22997 45574
rect 23049 45880 23083 45896
rect 23049 45812 23083 45818
rect 23049 45744 23083 45746
rect 23049 45708 23083 45710
rect 23049 45636 23083 45642
rect 23160 45852 23194 45862
rect 23160 45780 23194 45812
rect 23160 45710 23194 45744
rect 23160 45642 23194 45674
rect 23160 45592 23194 45602
rect 23049 45558 23083 45574
rect 22879 45490 22891 45524
rect 22929 45490 22963 45524
rect 22997 45490 23031 45524
rect 23069 45490 23081 45524
rect 32077 45880 32111 45896
rect 31966 45852 32000 45862
rect 31966 45780 32000 45812
rect 31966 45710 32000 45744
rect 31966 45642 32000 45674
rect 31966 45592 32000 45602
rect 32077 45812 32111 45818
rect 32077 45744 32111 45746
rect 32077 45708 32111 45710
rect 32077 45636 32111 45642
rect 32077 45558 32111 45574
rect 32163 45880 32197 45896
rect 32163 45812 32197 45818
rect 32163 45744 32197 45746
rect 32163 45708 32197 45710
rect 32163 45636 32197 45642
rect 32163 45558 32197 45574
rect 32249 45880 32283 45896
rect 32249 45812 32283 45818
rect 32249 45744 32283 45746
rect 32249 45708 32283 45710
rect 32249 45636 32283 45642
rect 32360 45852 32394 45862
rect 32360 45780 32394 45812
rect 32360 45710 32394 45744
rect 32360 45642 32394 45674
rect 32360 45592 32394 45602
rect 32249 45558 32283 45574
rect 32079 45490 32091 45524
rect 32129 45490 32163 45524
rect 32197 45490 32231 45524
rect 32269 45490 32281 45524
rect 41277 45880 41311 45896
rect 41166 45852 41200 45862
rect 41166 45780 41200 45812
rect 41166 45710 41200 45744
rect 41166 45642 41200 45674
rect 41166 45592 41200 45602
rect 41277 45812 41311 45818
rect 41277 45744 41311 45746
rect 41277 45708 41311 45710
rect 41277 45636 41311 45642
rect 41277 45558 41311 45574
rect 41363 45880 41397 45896
rect 41363 45812 41397 45818
rect 41363 45744 41397 45746
rect 41363 45708 41397 45710
rect 41363 45636 41397 45642
rect 41363 45558 41397 45574
rect 41449 45880 41483 45896
rect 41449 45812 41483 45818
rect 41449 45744 41483 45746
rect 41449 45708 41483 45710
rect 41449 45636 41483 45642
rect 41560 45852 41594 45862
rect 41560 45780 41594 45812
rect 41560 45710 41594 45744
rect 41560 45642 41594 45674
rect 41560 45592 41594 45602
rect 41449 45558 41483 45574
rect 41279 45490 41291 45524
rect 41329 45490 41363 45524
rect 41397 45490 41431 45524
rect 41469 45490 41481 45524
rect 50477 45880 50511 45896
rect 50366 45852 50400 45862
rect 50366 45780 50400 45812
rect 50366 45710 50400 45744
rect 50366 45642 50400 45674
rect 50366 45592 50400 45602
rect 50477 45812 50511 45818
rect 50477 45744 50511 45746
rect 50477 45708 50511 45710
rect 50477 45636 50511 45642
rect 50477 45558 50511 45574
rect 50563 45880 50597 45896
rect 50563 45812 50597 45818
rect 50563 45744 50597 45746
rect 50563 45708 50597 45710
rect 50563 45636 50597 45642
rect 50563 45558 50597 45574
rect 50649 45880 50683 45896
rect 50649 45812 50683 45818
rect 50649 45744 50683 45746
rect 50649 45708 50683 45710
rect 50649 45636 50683 45642
rect 50760 45852 50794 45862
rect 50760 45780 50794 45812
rect 50760 45710 50794 45744
rect 50760 45642 50794 45674
rect 50760 45592 50794 45602
rect 50649 45558 50683 45574
rect 50479 45490 50491 45524
rect 50529 45490 50563 45524
rect 50597 45490 50631 45524
rect 50669 45490 50681 45524
rect 59677 45880 59711 45896
rect 59566 45852 59600 45862
rect 59566 45780 59600 45812
rect 59566 45710 59600 45744
rect 59566 45642 59600 45674
rect 59566 45592 59600 45602
rect 59677 45812 59711 45818
rect 59677 45744 59711 45746
rect 59677 45708 59711 45710
rect 59677 45636 59711 45642
rect 59677 45558 59711 45574
rect 59763 45880 59797 45896
rect 59763 45812 59797 45818
rect 59763 45744 59797 45746
rect 59763 45708 59797 45710
rect 59763 45636 59797 45642
rect 59763 45558 59797 45574
rect 59849 45880 59883 45896
rect 59849 45812 59883 45818
rect 59849 45744 59883 45746
rect 59849 45708 59883 45710
rect 59849 45636 59883 45642
rect 59960 45852 59994 45862
rect 59960 45780 59994 45812
rect 59960 45710 59994 45744
rect 59960 45642 59994 45674
rect 59960 45592 59994 45602
rect 59849 45558 59883 45574
rect 59679 45490 59691 45524
rect 59729 45490 59763 45524
rect 59797 45490 59831 45524
rect 59869 45490 59881 45524
rect 68877 45880 68911 45896
rect 68766 45852 68800 45862
rect 68766 45780 68800 45812
rect 68766 45710 68800 45744
rect 68766 45642 68800 45674
rect 68766 45592 68800 45602
rect 68877 45812 68911 45818
rect 68877 45744 68911 45746
rect 68877 45708 68911 45710
rect 68877 45636 68911 45642
rect 68877 45558 68911 45574
rect 68963 45880 68997 45896
rect 68963 45812 68997 45818
rect 68963 45744 68997 45746
rect 68963 45708 68997 45710
rect 68963 45636 68997 45642
rect 68963 45558 68997 45574
rect 69049 45880 69083 45896
rect 69049 45812 69083 45818
rect 69049 45744 69083 45746
rect 69049 45708 69083 45710
rect 69049 45636 69083 45642
rect 69160 45852 69194 45862
rect 69160 45780 69194 45812
rect 69160 45710 69194 45744
rect 69160 45642 69194 45674
rect 69160 45592 69194 45602
rect 69049 45558 69083 45574
rect 68879 45490 68891 45524
rect 68929 45490 68963 45524
rect 68997 45490 69031 45524
rect 69069 45490 69081 45524
rect -336 45392 -302 45408
rect -508 45350 -390 45352
rect -560 45320 -390 45350
rect -610 45312 -390 45320
rect -610 45310 -490 45312
rect -424 45254 -390 45312
rect -240 45340 -160 45360
rect -240 45300 -220 45340
rect -180 45300 -160 45340
rect -240 45280 -160 45300
rect -424 44962 -390 44978
rect -336 45254 -302 45270
rect -336 44898 -302 44978
rect -506 44890 -218 44898
rect -506 44840 -440 44890
rect -390 44876 -330 44890
rect -390 44840 -338 44876
rect -280 44840 -218 44890
rect -506 44820 -218 44840
rect 4479 36050 4491 36084
rect 4529 36050 4563 36084
rect 4597 36050 4631 36084
rect 4669 36050 4681 36084
rect 13679 36050 13691 36084
rect 13729 36050 13763 36084
rect 13797 36050 13831 36084
rect 13869 36050 13881 36084
rect 22879 36050 22891 36084
rect 22929 36050 22963 36084
rect 22997 36050 23031 36084
rect 23069 36050 23081 36084
rect 32079 36050 32091 36084
rect 32129 36050 32163 36084
rect 32197 36050 32231 36084
rect 32269 36050 32281 36084
rect 41279 36050 41291 36084
rect 41329 36050 41363 36084
rect 41397 36050 41431 36084
rect 41469 36050 41481 36084
rect 50479 36050 50491 36084
rect 50529 36050 50563 36084
rect 50597 36050 50631 36084
rect 50669 36050 50681 36084
rect 59679 36050 59691 36084
rect 59729 36050 59763 36084
rect 59797 36050 59831 36084
rect 59869 36050 59881 36084
rect 68879 36050 68891 36084
rect 68929 36050 68963 36084
rect 68997 36050 69031 36084
rect 69069 36050 69081 36084
rect 4477 36000 4511 36016
rect 4366 35972 4400 35982
rect 4366 35900 4400 35932
rect 4366 35830 4400 35864
rect 4366 35762 4400 35794
rect 4366 35712 4400 35722
rect 4477 35932 4511 35938
rect 4477 35864 4511 35866
rect 4477 35828 4511 35830
rect 4477 35756 4511 35762
rect 4477 35678 4511 35694
rect 4563 36000 4597 36016
rect 4563 35932 4597 35938
rect 4563 35864 4597 35866
rect 4563 35828 4597 35830
rect 4563 35756 4597 35762
rect 4563 35678 4597 35694
rect 4649 36000 4683 36016
rect 4649 35932 4683 35938
rect 4649 35864 4683 35866
rect 4649 35828 4683 35830
rect 4649 35756 4683 35762
rect 4760 35972 4794 35982
rect 4760 35900 4794 35932
rect 4760 35830 4794 35864
rect 4760 35762 4794 35794
rect 4760 35712 4794 35722
rect 4649 35678 4683 35694
rect 4479 35610 4491 35644
rect 4529 35610 4563 35644
rect 4597 35610 4631 35644
rect 4669 35610 4681 35644
rect 13677 36000 13711 36016
rect 13566 35972 13600 35982
rect 13566 35900 13600 35932
rect 13566 35830 13600 35864
rect 13566 35762 13600 35794
rect 13566 35712 13600 35722
rect 13677 35932 13711 35938
rect 13677 35864 13711 35866
rect 13677 35828 13711 35830
rect 13677 35756 13711 35762
rect 13677 35678 13711 35694
rect 13763 36000 13797 36016
rect 13763 35932 13797 35938
rect 13763 35864 13797 35866
rect 13763 35828 13797 35830
rect 13763 35756 13797 35762
rect 13763 35678 13797 35694
rect 13849 36000 13883 36016
rect 13849 35932 13883 35938
rect 13849 35864 13883 35866
rect 13849 35828 13883 35830
rect 13849 35756 13883 35762
rect 13960 35972 13994 35982
rect 13960 35900 13994 35932
rect 13960 35830 13994 35864
rect 13960 35762 13994 35794
rect 13960 35712 13994 35722
rect 13849 35678 13883 35694
rect 13679 35610 13691 35644
rect 13729 35610 13763 35644
rect 13797 35610 13831 35644
rect 13869 35610 13881 35644
rect 22877 36000 22911 36016
rect 22766 35972 22800 35982
rect 22766 35900 22800 35932
rect 22766 35830 22800 35864
rect 22766 35762 22800 35794
rect 22766 35712 22800 35722
rect 22877 35932 22911 35938
rect 22877 35864 22911 35866
rect 22877 35828 22911 35830
rect 22877 35756 22911 35762
rect 22877 35678 22911 35694
rect 22963 36000 22997 36016
rect 22963 35932 22997 35938
rect 22963 35864 22997 35866
rect 22963 35828 22997 35830
rect 22963 35756 22997 35762
rect 22963 35678 22997 35694
rect 23049 36000 23083 36016
rect 23049 35932 23083 35938
rect 23049 35864 23083 35866
rect 23049 35828 23083 35830
rect 23049 35756 23083 35762
rect 23160 35972 23194 35982
rect 23160 35900 23194 35932
rect 23160 35830 23194 35864
rect 23160 35762 23194 35794
rect 23160 35712 23194 35722
rect 23049 35678 23083 35694
rect 22879 35610 22891 35644
rect 22929 35610 22963 35644
rect 22997 35610 23031 35644
rect 23069 35610 23081 35644
rect 32077 36000 32111 36016
rect 31966 35972 32000 35982
rect 31966 35900 32000 35932
rect 31966 35830 32000 35864
rect 31966 35762 32000 35794
rect 31966 35712 32000 35722
rect 32077 35932 32111 35938
rect 32077 35864 32111 35866
rect 32077 35828 32111 35830
rect 32077 35756 32111 35762
rect 32077 35678 32111 35694
rect 32163 36000 32197 36016
rect 32163 35932 32197 35938
rect 32163 35864 32197 35866
rect 32163 35828 32197 35830
rect 32163 35756 32197 35762
rect 32163 35678 32197 35694
rect 32249 36000 32283 36016
rect 32249 35932 32283 35938
rect 32249 35864 32283 35866
rect 32249 35828 32283 35830
rect 32249 35756 32283 35762
rect 32360 35972 32394 35982
rect 32360 35900 32394 35932
rect 32360 35830 32394 35864
rect 32360 35762 32394 35794
rect 32360 35712 32394 35722
rect 32249 35678 32283 35694
rect 32079 35610 32091 35644
rect 32129 35610 32163 35644
rect 32197 35610 32231 35644
rect 32269 35610 32281 35644
rect 41277 36000 41311 36016
rect 41166 35972 41200 35982
rect 41166 35900 41200 35932
rect 41166 35830 41200 35864
rect 41166 35762 41200 35794
rect 41166 35712 41200 35722
rect 41277 35932 41311 35938
rect 41277 35864 41311 35866
rect 41277 35828 41311 35830
rect 41277 35756 41311 35762
rect 41277 35678 41311 35694
rect 41363 36000 41397 36016
rect 41363 35932 41397 35938
rect 41363 35864 41397 35866
rect 41363 35828 41397 35830
rect 41363 35756 41397 35762
rect 41363 35678 41397 35694
rect 41449 36000 41483 36016
rect 41449 35932 41483 35938
rect 41449 35864 41483 35866
rect 41449 35828 41483 35830
rect 41449 35756 41483 35762
rect 41560 35972 41594 35982
rect 41560 35900 41594 35932
rect 41560 35830 41594 35864
rect 41560 35762 41594 35794
rect 41560 35712 41594 35722
rect 41449 35678 41483 35694
rect 41279 35610 41291 35644
rect 41329 35610 41363 35644
rect 41397 35610 41431 35644
rect 41469 35610 41481 35644
rect 50477 36000 50511 36016
rect 50366 35972 50400 35982
rect 50366 35900 50400 35932
rect 50366 35830 50400 35864
rect 50366 35762 50400 35794
rect 50366 35712 50400 35722
rect 50477 35932 50511 35938
rect 50477 35864 50511 35866
rect 50477 35828 50511 35830
rect 50477 35756 50511 35762
rect 50477 35678 50511 35694
rect 50563 36000 50597 36016
rect 50563 35932 50597 35938
rect 50563 35864 50597 35866
rect 50563 35828 50597 35830
rect 50563 35756 50597 35762
rect 50563 35678 50597 35694
rect 50649 36000 50683 36016
rect 50649 35932 50683 35938
rect 50649 35864 50683 35866
rect 50649 35828 50683 35830
rect 50649 35756 50683 35762
rect 50760 35972 50794 35982
rect 50760 35900 50794 35932
rect 50760 35830 50794 35864
rect 50760 35762 50794 35794
rect 50760 35712 50794 35722
rect 50649 35678 50683 35694
rect 50479 35610 50491 35644
rect 50529 35610 50563 35644
rect 50597 35610 50631 35644
rect 50669 35610 50681 35644
rect 59677 36000 59711 36016
rect 59566 35972 59600 35982
rect 59566 35900 59600 35932
rect 59566 35830 59600 35864
rect 59566 35762 59600 35794
rect 59566 35712 59600 35722
rect 59677 35932 59711 35938
rect 59677 35864 59711 35866
rect 59677 35828 59711 35830
rect 59677 35756 59711 35762
rect 59677 35678 59711 35694
rect 59763 36000 59797 36016
rect 59763 35932 59797 35938
rect 59763 35864 59797 35866
rect 59763 35828 59797 35830
rect 59763 35756 59797 35762
rect 59763 35678 59797 35694
rect 59849 36000 59883 36016
rect 59849 35932 59883 35938
rect 59849 35864 59883 35866
rect 59849 35828 59883 35830
rect 59849 35756 59883 35762
rect 59960 35972 59994 35982
rect 59960 35900 59994 35932
rect 59960 35830 59994 35864
rect 59960 35762 59994 35794
rect 59960 35712 59994 35722
rect 59849 35678 59883 35694
rect 59679 35610 59691 35644
rect 59729 35610 59763 35644
rect 59797 35610 59831 35644
rect 59869 35610 59881 35644
rect 68877 36000 68911 36016
rect 68766 35972 68800 35982
rect 68766 35900 68800 35932
rect 68766 35830 68800 35864
rect 68766 35762 68800 35794
rect 68766 35712 68800 35722
rect 68877 35932 68911 35938
rect 68877 35864 68911 35866
rect 68877 35828 68911 35830
rect 68877 35756 68911 35762
rect 68877 35678 68911 35694
rect 68963 36000 68997 36016
rect 68963 35932 68997 35938
rect 68963 35864 68997 35866
rect 68963 35828 68997 35830
rect 68963 35756 68997 35762
rect 68963 35678 68997 35694
rect 69049 36000 69083 36016
rect 69049 35932 69083 35938
rect 69049 35864 69083 35866
rect 69049 35828 69083 35830
rect 69049 35756 69083 35762
rect 69160 35972 69194 35982
rect 69160 35900 69194 35932
rect 69160 35830 69194 35864
rect 69160 35762 69194 35794
rect 69160 35712 69194 35722
rect 69049 35678 69083 35694
rect 68879 35610 68891 35644
rect 68929 35610 68963 35644
rect 68997 35610 69031 35644
rect 69069 35610 69081 35644
rect 4479 26170 4491 26204
rect 4529 26170 4563 26204
rect 4597 26170 4631 26204
rect 4669 26170 4681 26204
rect 13679 26170 13691 26204
rect 13729 26170 13763 26204
rect 13797 26170 13831 26204
rect 13869 26170 13881 26204
rect 22879 26170 22891 26204
rect 22929 26170 22963 26204
rect 22997 26170 23031 26204
rect 23069 26170 23081 26204
rect 32079 26170 32091 26204
rect 32129 26170 32163 26204
rect 32197 26170 32231 26204
rect 32269 26170 32281 26204
rect 41279 26170 41291 26204
rect 41329 26170 41363 26204
rect 41397 26170 41431 26204
rect 41469 26170 41481 26204
rect 50479 26170 50491 26204
rect 50529 26170 50563 26204
rect 50597 26170 50631 26204
rect 50669 26170 50681 26204
rect 59679 26170 59691 26204
rect 59729 26170 59763 26204
rect 59797 26170 59831 26204
rect 59869 26170 59881 26204
rect 68879 26170 68891 26204
rect 68929 26170 68963 26204
rect 68997 26170 69031 26204
rect 69069 26170 69081 26204
rect 4477 26120 4511 26136
rect 4366 26092 4400 26102
rect 4366 26020 4400 26052
rect 4366 25950 4400 25984
rect 4366 25882 4400 25914
rect 4366 25832 4400 25842
rect 4477 26052 4511 26058
rect 4477 25984 4511 25986
rect 4477 25948 4511 25950
rect 4477 25876 4511 25882
rect 4477 25798 4511 25814
rect 4563 26120 4597 26136
rect 4563 26052 4597 26058
rect 4563 25984 4597 25986
rect 4563 25948 4597 25950
rect 4563 25876 4597 25882
rect 4563 25798 4597 25814
rect 4649 26120 4683 26136
rect 4649 26052 4683 26058
rect 4649 25984 4683 25986
rect 4649 25948 4683 25950
rect 4649 25876 4683 25882
rect 4760 26092 4794 26102
rect 4760 26020 4794 26052
rect 4760 25950 4794 25984
rect 4760 25882 4794 25914
rect 4760 25832 4794 25842
rect 4649 25798 4683 25814
rect 4479 25730 4491 25764
rect 4529 25730 4563 25764
rect 4597 25730 4631 25764
rect 4669 25730 4681 25764
rect 13677 26120 13711 26136
rect 13566 26092 13600 26102
rect 13566 26020 13600 26052
rect 13566 25950 13600 25984
rect 13566 25882 13600 25914
rect 13566 25832 13600 25842
rect 13677 26052 13711 26058
rect 13677 25984 13711 25986
rect 13677 25948 13711 25950
rect 13677 25876 13711 25882
rect 13677 25798 13711 25814
rect 13763 26120 13797 26136
rect 13763 26052 13797 26058
rect 13763 25984 13797 25986
rect 13763 25948 13797 25950
rect 13763 25876 13797 25882
rect 13763 25798 13797 25814
rect 13849 26120 13883 26136
rect 13849 26052 13883 26058
rect 13849 25984 13883 25986
rect 13849 25948 13883 25950
rect 13849 25876 13883 25882
rect 13960 26092 13994 26102
rect 13960 26020 13994 26052
rect 13960 25950 13994 25984
rect 13960 25882 13994 25914
rect 13960 25832 13994 25842
rect 13849 25798 13883 25814
rect 13679 25730 13691 25764
rect 13729 25730 13763 25764
rect 13797 25730 13831 25764
rect 13869 25730 13881 25764
rect 22877 26120 22911 26136
rect 22766 26092 22800 26102
rect 22766 26020 22800 26052
rect 22766 25950 22800 25984
rect 22766 25882 22800 25914
rect 22766 25832 22800 25842
rect 22877 26052 22911 26058
rect 22877 25984 22911 25986
rect 22877 25948 22911 25950
rect 22877 25876 22911 25882
rect 22877 25798 22911 25814
rect 22963 26120 22997 26136
rect 22963 26052 22997 26058
rect 22963 25984 22997 25986
rect 22963 25948 22997 25950
rect 22963 25876 22997 25882
rect 22963 25798 22997 25814
rect 23049 26120 23083 26136
rect 23049 26052 23083 26058
rect 23049 25984 23083 25986
rect 23049 25948 23083 25950
rect 23049 25876 23083 25882
rect 23160 26092 23194 26102
rect 23160 26020 23194 26052
rect 23160 25950 23194 25984
rect 23160 25882 23194 25914
rect 23160 25832 23194 25842
rect 23049 25798 23083 25814
rect 22879 25730 22891 25764
rect 22929 25730 22963 25764
rect 22997 25730 23031 25764
rect 23069 25730 23081 25764
rect 32077 26120 32111 26136
rect 31966 26092 32000 26102
rect 31966 26020 32000 26052
rect 31966 25950 32000 25984
rect 31966 25882 32000 25914
rect 31966 25832 32000 25842
rect 32077 26052 32111 26058
rect 32077 25984 32111 25986
rect 32077 25948 32111 25950
rect 32077 25876 32111 25882
rect 32077 25798 32111 25814
rect 32163 26120 32197 26136
rect 32163 26052 32197 26058
rect 32163 25984 32197 25986
rect 32163 25948 32197 25950
rect 32163 25876 32197 25882
rect 32163 25798 32197 25814
rect 32249 26120 32283 26136
rect 32249 26052 32283 26058
rect 32249 25984 32283 25986
rect 32249 25948 32283 25950
rect 32249 25876 32283 25882
rect 32360 26092 32394 26102
rect 32360 26020 32394 26052
rect 32360 25950 32394 25984
rect 32360 25882 32394 25914
rect 32360 25832 32394 25842
rect 32249 25798 32283 25814
rect 32079 25730 32091 25764
rect 32129 25730 32163 25764
rect 32197 25730 32231 25764
rect 32269 25730 32281 25764
rect 41277 26120 41311 26136
rect 41166 26092 41200 26102
rect 41166 26020 41200 26052
rect 41166 25950 41200 25984
rect 41166 25882 41200 25914
rect 41166 25832 41200 25842
rect 41277 26052 41311 26058
rect 41277 25984 41311 25986
rect 41277 25948 41311 25950
rect 41277 25876 41311 25882
rect 41277 25798 41311 25814
rect 41363 26120 41397 26136
rect 41363 26052 41397 26058
rect 41363 25984 41397 25986
rect 41363 25948 41397 25950
rect 41363 25876 41397 25882
rect 41363 25798 41397 25814
rect 41449 26120 41483 26136
rect 41449 26052 41483 26058
rect 41449 25984 41483 25986
rect 41449 25948 41483 25950
rect 41449 25876 41483 25882
rect 41560 26092 41594 26102
rect 41560 26020 41594 26052
rect 41560 25950 41594 25984
rect 41560 25882 41594 25914
rect 41560 25832 41594 25842
rect 41449 25798 41483 25814
rect 41279 25730 41291 25764
rect 41329 25730 41363 25764
rect 41397 25730 41431 25764
rect 41469 25730 41481 25764
rect 50477 26120 50511 26136
rect 50366 26092 50400 26102
rect 50366 26020 50400 26052
rect 50366 25950 50400 25984
rect 50366 25882 50400 25914
rect 50366 25832 50400 25842
rect 50477 26052 50511 26058
rect 50477 25984 50511 25986
rect 50477 25948 50511 25950
rect 50477 25876 50511 25882
rect 50477 25798 50511 25814
rect 50563 26120 50597 26136
rect 50563 26052 50597 26058
rect 50563 25984 50597 25986
rect 50563 25948 50597 25950
rect 50563 25876 50597 25882
rect 50563 25798 50597 25814
rect 50649 26120 50683 26136
rect 50649 26052 50683 26058
rect 50649 25984 50683 25986
rect 50649 25948 50683 25950
rect 50649 25876 50683 25882
rect 50760 26092 50794 26102
rect 50760 26020 50794 26052
rect 50760 25950 50794 25984
rect 50760 25882 50794 25914
rect 50760 25832 50794 25842
rect 50649 25798 50683 25814
rect 50479 25730 50491 25764
rect 50529 25730 50563 25764
rect 50597 25730 50631 25764
rect 50669 25730 50681 25764
rect 59677 26120 59711 26136
rect 59566 26092 59600 26102
rect 59566 26020 59600 26052
rect 59566 25950 59600 25984
rect 59566 25882 59600 25914
rect 59566 25832 59600 25842
rect 59677 26052 59711 26058
rect 59677 25984 59711 25986
rect 59677 25948 59711 25950
rect 59677 25876 59711 25882
rect 59677 25798 59711 25814
rect 59763 26120 59797 26136
rect 59763 26052 59797 26058
rect 59763 25984 59797 25986
rect 59763 25948 59797 25950
rect 59763 25876 59797 25882
rect 59763 25798 59797 25814
rect 59849 26120 59883 26136
rect 59849 26052 59883 26058
rect 59849 25984 59883 25986
rect 59849 25948 59883 25950
rect 59849 25876 59883 25882
rect 59960 26092 59994 26102
rect 59960 26020 59994 26052
rect 59960 25950 59994 25984
rect 59960 25882 59994 25914
rect 59960 25832 59994 25842
rect 59849 25798 59883 25814
rect 59679 25730 59691 25764
rect 59729 25730 59763 25764
rect 59797 25730 59831 25764
rect 59869 25730 59881 25764
rect 68877 26120 68911 26136
rect 68766 26092 68800 26102
rect 68766 26020 68800 26052
rect 68766 25950 68800 25984
rect 68766 25882 68800 25914
rect 68766 25832 68800 25842
rect 68877 26052 68911 26058
rect 68877 25984 68911 25986
rect 68877 25948 68911 25950
rect 68877 25876 68911 25882
rect 68877 25798 68911 25814
rect 68963 26120 68997 26136
rect 68963 26052 68997 26058
rect 68963 25984 68997 25986
rect 68963 25948 68997 25950
rect 68963 25876 68997 25882
rect 68963 25798 68997 25814
rect 69049 26120 69083 26136
rect 69049 26052 69083 26058
rect 69049 25984 69083 25986
rect 69049 25948 69083 25950
rect 69049 25876 69083 25882
rect 69160 26092 69194 26102
rect 69160 26020 69194 26052
rect 69160 25950 69194 25984
rect 69160 25882 69194 25914
rect 69160 25832 69194 25842
rect 69049 25798 69083 25814
rect 68879 25730 68891 25764
rect 68929 25730 68963 25764
rect 68997 25730 69031 25764
rect 69069 25730 69081 25764
rect 4479 16290 4491 16324
rect 4529 16290 4563 16324
rect 4597 16290 4631 16324
rect 4669 16290 4681 16324
rect 13679 16290 13691 16324
rect 13729 16290 13763 16324
rect 13797 16290 13831 16324
rect 13869 16290 13881 16324
rect 22879 16290 22891 16324
rect 22929 16290 22963 16324
rect 22997 16290 23031 16324
rect 23069 16290 23081 16324
rect 32079 16290 32091 16324
rect 32129 16290 32163 16324
rect 32197 16290 32231 16324
rect 32269 16290 32281 16324
rect 41279 16290 41291 16324
rect 41329 16290 41363 16324
rect 41397 16290 41431 16324
rect 41469 16290 41481 16324
rect 50479 16290 50491 16324
rect 50529 16290 50563 16324
rect 50597 16290 50631 16324
rect 50669 16290 50681 16324
rect 59679 16290 59691 16324
rect 59729 16290 59763 16324
rect 59797 16290 59831 16324
rect 59869 16290 59881 16324
rect 68879 16290 68891 16324
rect 68929 16290 68963 16324
rect 68997 16290 69031 16324
rect 69069 16290 69081 16324
rect 4477 16240 4511 16256
rect 4366 16212 4400 16222
rect 4366 16140 4400 16172
rect 4366 16070 4400 16104
rect 4366 16002 4400 16034
rect 4366 15952 4400 15962
rect 4477 16172 4511 16178
rect 4477 16104 4511 16106
rect 4477 16068 4511 16070
rect 4477 15996 4511 16002
rect 4477 15918 4511 15934
rect 4563 16240 4597 16256
rect 4563 16172 4597 16178
rect 4563 16104 4597 16106
rect 4563 16068 4597 16070
rect 4563 15996 4597 16002
rect 4563 15918 4597 15934
rect 4649 16240 4683 16256
rect 4649 16172 4683 16178
rect 4649 16104 4683 16106
rect 4649 16068 4683 16070
rect 4649 15996 4683 16002
rect 4760 16212 4794 16222
rect 4760 16140 4794 16172
rect 4760 16070 4794 16104
rect 4760 16002 4794 16034
rect 4760 15952 4794 15962
rect 4649 15918 4683 15934
rect 4479 15850 4491 15884
rect 4529 15850 4563 15884
rect 4597 15850 4631 15884
rect 4669 15850 4681 15884
rect 13677 16240 13711 16256
rect 13566 16212 13600 16222
rect 13566 16140 13600 16172
rect 13566 16070 13600 16104
rect 13566 16002 13600 16034
rect 13566 15952 13600 15962
rect 13677 16172 13711 16178
rect 13677 16104 13711 16106
rect 13677 16068 13711 16070
rect 13677 15996 13711 16002
rect 13677 15918 13711 15934
rect 13763 16240 13797 16256
rect 13763 16172 13797 16178
rect 13763 16104 13797 16106
rect 13763 16068 13797 16070
rect 13763 15996 13797 16002
rect 13763 15918 13797 15934
rect 13849 16240 13883 16256
rect 13849 16172 13883 16178
rect 13849 16104 13883 16106
rect 13849 16068 13883 16070
rect 13849 15996 13883 16002
rect 13960 16212 13994 16222
rect 13960 16140 13994 16172
rect 13960 16070 13994 16104
rect 13960 16002 13994 16034
rect 13960 15952 13994 15962
rect 13849 15918 13883 15934
rect 13679 15850 13691 15884
rect 13729 15850 13763 15884
rect 13797 15850 13831 15884
rect 13869 15850 13881 15884
rect 22877 16240 22911 16256
rect 22766 16212 22800 16222
rect 22766 16140 22800 16172
rect 22766 16070 22800 16104
rect 22766 16002 22800 16034
rect 22766 15952 22800 15962
rect 22877 16172 22911 16178
rect 22877 16104 22911 16106
rect 22877 16068 22911 16070
rect 22877 15996 22911 16002
rect 22877 15918 22911 15934
rect 22963 16240 22997 16256
rect 22963 16172 22997 16178
rect 22963 16104 22997 16106
rect 22963 16068 22997 16070
rect 22963 15996 22997 16002
rect 22963 15918 22997 15934
rect 23049 16240 23083 16256
rect 23049 16172 23083 16178
rect 23049 16104 23083 16106
rect 23049 16068 23083 16070
rect 23049 15996 23083 16002
rect 23160 16212 23194 16222
rect 23160 16140 23194 16172
rect 23160 16070 23194 16104
rect 23160 16002 23194 16034
rect 23160 15952 23194 15962
rect 23049 15918 23083 15934
rect 22879 15850 22891 15884
rect 22929 15850 22963 15884
rect 22997 15850 23031 15884
rect 23069 15850 23081 15884
rect 32077 16240 32111 16256
rect 31966 16212 32000 16222
rect 31966 16140 32000 16172
rect 31966 16070 32000 16104
rect 31966 16002 32000 16034
rect 31966 15952 32000 15962
rect 32077 16172 32111 16178
rect 32077 16104 32111 16106
rect 32077 16068 32111 16070
rect 32077 15996 32111 16002
rect 32077 15918 32111 15934
rect 32163 16240 32197 16256
rect 32163 16172 32197 16178
rect 32163 16104 32197 16106
rect 32163 16068 32197 16070
rect 32163 15996 32197 16002
rect 32163 15918 32197 15934
rect 32249 16240 32283 16256
rect 32249 16172 32283 16178
rect 32249 16104 32283 16106
rect 32249 16068 32283 16070
rect 32249 15996 32283 16002
rect 32360 16212 32394 16222
rect 32360 16140 32394 16172
rect 32360 16070 32394 16104
rect 32360 16002 32394 16034
rect 32360 15952 32394 15962
rect 32249 15918 32283 15934
rect 32079 15850 32091 15884
rect 32129 15850 32163 15884
rect 32197 15850 32231 15884
rect 32269 15850 32281 15884
rect 41277 16240 41311 16256
rect 41166 16212 41200 16222
rect 41166 16140 41200 16172
rect 41166 16070 41200 16104
rect 41166 16002 41200 16034
rect 41166 15952 41200 15962
rect 41277 16172 41311 16178
rect 41277 16104 41311 16106
rect 41277 16068 41311 16070
rect 41277 15996 41311 16002
rect 41277 15918 41311 15934
rect 41363 16240 41397 16256
rect 41363 16172 41397 16178
rect 41363 16104 41397 16106
rect 41363 16068 41397 16070
rect 41363 15996 41397 16002
rect 41363 15918 41397 15934
rect 41449 16240 41483 16256
rect 41449 16172 41483 16178
rect 41449 16104 41483 16106
rect 41449 16068 41483 16070
rect 41449 15996 41483 16002
rect 41560 16212 41594 16222
rect 41560 16140 41594 16172
rect 41560 16070 41594 16104
rect 41560 16002 41594 16034
rect 41560 15952 41594 15962
rect 41449 15918 41483 15934
rect 41279 15850 41291 15884
rect 41329 15850 41363 15884
rect 41397 15850 41431 15884
rect 41469 15850 41481 15884
rect 50477 16240 50511 16256
rect 50366 16212 50400 16222
rect 50366 16140 50400 16172
rect 50366 16070 50400 16104
rect 50366 16002 50400 16034
rect 50366 15952 50400 15962
rect 50477 16172 50511 16178
rect 50477 16104 50511 16106
rect 50477 16068 50511 16070
rect 50477 15996 50511 16002
rect 50477 15918 50511 15934
rect 50563 16240 50597 16256
rect 50563 16172 50597 16178
rect 50563 16104 50597 16106
rect 50563 16068 50597 16070
rect 50563 15996 50597 16002
rect 50563 15918 50597 15934
rect 50649 16240 50683 16256
rect 50649 16172 50683 16178
rect 50649 16104 50683 16106
rect 50649 16068 50683 16070
rect 50649 15996 50683 16002
rect 50760 16212 50794 16222
rect 50760 16140 50794 16172
rect 50760 16070 50794 16104
rect 50760 16002 50794 16034
rect 50760 15952 50794 15962
rect 50649 15918 50683 15934
rect 50479 15850 50491 15884
rect 50529 15850 50563 15884
rect 50597 15850 50631 15884
rect 50669 15850 50681 15884
rect 59677 16240 59711 16256
rect 59566 16212 59600 16222
rect 59566 16140 59600 16172
rect 59566 16070 59600 16104
rect 59566 16002 59600 16034
rect 59566 15952 59600 15962
rect 59677 16172 59711 16178
rect 59677 16104 59711 16106
rect 59677 16068 59711 16070
rect 59677 15996 59711 16002
rect 59677 15918 59711 15934
rect 59763 16240 59797 16256
rect 59763 16172 59797 16178
rect 59763 16104 59797 16106
rect 59763 16068 59797 16070
rect 59763 15996 59797 16002
rect 59763 15918 59797 15934
rect 59849 16240 59883 16256
rect 59849 16172 59883 16178
rect 59849 16104 59883 16106
rect 59849 16068 59883 16070
rect 59849 15996 59883 16002
rect 59960 16212 59994 16222
rect 59960 16140 59994 16172
rect 59960 16070 59994 16104
rect 59960 16002 59994 16034
rect 59960 15952 59994 15962
rect 59849 15918 59883 15934
rect 59679 15850 59691 15884
rect 59729 15850 59763 15884
rect 59797 15850 59831 15884
rect 59869 15850 59881 15884
rect 68877 16240 68911 16256
rect 68766 16212 68800 16222
rect 68766 16140 68800 16172
rect 68766 16070 68800 16104
rect 68766 16002 68800 16034
rect 68766 15952 68800 15962
rect 68877 16172 68911 16178
rect 68877 16104 68911 16106
rect 68877 16068 68911 16070
rect 68877 15996 68911 16002
rect 68877 15918 68911 15934
rect 68963 16240 68997 16256
rect 68963 16172 68997 16178
rect 68963 16104 68997 16106
rect 68963 16068 68997 16070
rect 68963 15996 68997 16002
rect 68963 15918 68997 15934
rect 69049 16240 69083 16256
rect 69049 16172 69083 16178
rect 69049 16104 69083 16106
rect 69049 16068 69083 16070
rect 69049 15996 69083 16002
rect 69160 16212 69194 16222
rect 69160 16140 69194 16172
rect 69160 16070 69194 16104
rect 69160 16002 69194 16034
rect 69160 15952 69194 15962
rect 69049 15918 69083 15934
rect 68879 15850 68891 15884
rect 68929 15850 68963 15884
rect 68997 15850 69031 15884
rect 69069 15850 69081 15884
rect -506 6612 -218 6640
rect -506 6610 -440 6612
rect -392 6610 -326 6612
rect -278 6610 -218 6612
rect -506 6570 -480 6610
rect -360 6574 -326 6610
rect -440 6570 -400 6574
rect -360 6570 -310 6574
rect -270 6570 -218 6610
rect -506 6538 -218 6570
rect -424 6464 -390 6480
rect -610 5840 -550 5850
rect -610 5800 -600 5840
rect -560 5830 -550 5840
rect -424 5832 -390 5888
rect -336 6464 -302 6538
rect 4479 6410 4491 6444
rect 4529 6410 4563 6444
rect 4597 6410 4631 6444
rect 4669 6410 4681 6444
rect 13679 6410 13691 6444
rect 13729 6410 13763 6444
rect 13797 6410 13831 6444
rect 13869 6410 13881 6444
rect 22879 6410 22891 6444
rect 22929 6410 22963 6444
rect 22997 6410 23031 6444
rect 23069 6410 23081 6444
rect 32079 6410 32091 6444
rect 32129 6410 32163 6444
rect 32197 6410 32231 6444
rect 32269 6410 32281 6444
rect 41279 6410 41291 6444
rect 41329 6410 41363 6444
rect 41397 6410 41431 6444
rect 41469 6410 41481 6444
rect 50479 6410 50491 6444
rect 50529 6410 50563 6444
rect 50597 6410 50631 6444
rect 50669 6410 50681 6444
rect 59679 6410 59691 6444
rect 59729 6410 59763 6444
rect 59797 6410 59831 6444
rect 59869 6410 59881 6444
rect 68879 6410 68891 6444
rect 68929 6410 68963 6444
rect 68997 6410 69031 6444
rect 69069 6410 69081 6444
rect 4477 6360 4511 6376
rect 4366 6332 4400 6342
rect 4366 6260 4400 6292
rect 4366 6190 4400 6224
rect 4366 6122 4400 6154
rect 4366 6072 4400 6082
rect 4477 6292 4511 6298
rect 4477 6224 4511 6226
rect 4477 6188 4511 6190
rect 4477 6116 4511 6122
rect 4477 6038 4511 6054
rect 4563 6360 4597 6376
rect 4563 6292 4597 6298
rect 4563 6224 4597 6226
rect 4563 6188 4597 6190
rect 4563 6116 4597 6122
rect 4563 6038 4597 6054
rect 4649 6360 4683 6376
rect 4649 6292 4683 6298
rect 4649 6224 4683 6226
rect 4649 6188 4683 6190
rect 4649 6116 4683 6122
rect 4760 6332 4794 6342
rect 4760 6260 4794 6292
rect 4760 6190 4794 6224
rect 4760 6122 4794 6154
rect 4760 6072 4794 6082
rect 4649 6038 4683 6054
rect 4479 5970 4491 6004
rect 4529 5970 4563 6004
rect 4597 5970 4631 6004
rect 4669 5970 4681 6004
rect 13677 6360 13711 6376
rect 13566 6332 13600 6342
rect 13566 6260 13600 6292
rect 13566 6190 13600 6224
rect 13566 6122 13600 6154
rect 13566 6072 13600 6082
rect 13677 6292 13711 6298
rect 13677 6224 13711 6226
rect 13677 6188 13711 6190
rect 13677 6116 13711 6122
rect 13677 6038 13711 6054
rect 13763 6360 13797 6376
rect 13763 6292 13797 6298
rect 13763 6224 13797 6226
rect 13763 6188 13797 6190
rect 13763 6116 13797 6122
rect 13763 6038 13797 6054
rect 13849 6360 13883 6376
rect 13849 6292 13883 6298
rect 13849 6224 13883 6226
rect 13849 6188 13883 6190
rect 13849 6116 13883 6122
rect 13960 6332 13994 6342
rect 13960 6260 13994 6292
rect 13960 6190 13994 6224
rect 13960 6122 13994 6154
rect 13960 6072 13994 6082
rect 13849 6038 13883 6054
rect 13679 5970 13691 6004
rect 13729 5970 13763 6004
rect 13797 5970 13831 6004
rect 13869 5970 13881 6004
rect 22877 6360 22911 6376
rect 22766 6332 22800 6342
rect 22766 6260 22800 6292
rect 22766 6190 22800 6224
rect 22766 6122 22800 6154
rect 22766 6072 22800 6082
rect 22877 6292 22911 6298
rect 22877 6224 22911 6226
rect 22877 6188 22911 6190
rect 22877 6116 22911 6122
rect 22877 6038 22911 6054
rect 22963 6360 22997 6376
rect 22963 6292 22997 6298
rect 22963 6224 22997 6226
rect 22963 6188 22997 6190
rect 22963 6116 22997 6122
rect 22963 6038 22997 6054
rect 23049 6360 23083 6376
rect 23049 6292 23083 6298
rect 23049 6224 23083 6226
rect 23049 6188 23083 6190
rect 23049 6116 23083 6122
rect 23160 6332 23194 6342
rect 23160 6260 23194 6292
rect 23160 6190 23194 6224
rect 23160 6122 23194 6154
rect 23160 6072 23194 6082
rect 23049 6038 23083 6054
rect 22879 5970 22891 6004
rect 22929 5970 22963 6004
rect 22997 5970 23031 6004
rect 23069 5970 23081 6004
rect 32077 6360 32111 6376
rect 31966 6332 32000 6342
rect 31966 6260 32000 6292
rect 31966 6190 32000 6224
rect 31966 6122 32000 6154
rect 31966 6072 32000 6082
rect 32077 6292 32111 6298
rect 32077 6224 32111 6226
rect 32077 6188 32111 6190
rect 32077 6116 32111 6122
rect 32077 6038 32111 6054
rect 32163 6360 32197 6376
rect 32163 6292 32197 6298
rect 32163 6224 32197 6226
rect 32163 6188 32197 6190
rect 32163 6116 32197 6122
rect 32163 6038 32197 6054
rect 32249 6360 32283 6376
rect 32249 6292 32283 6298
rect 32249 6224 32283 6226
rect 32249 6188 32283 6190
rect 32249 6116 32283 6122
rect 32360 6332 32394 6342
rect 32360 6260 32394 6292
rect 32360 6190 32394 6224
rect 32360 6122 32394 6154
rect 32360 6072 32394 6082
rect 32249 6038 32283 6054
rect 32079 5970 32091 6004
rect 32129 5970 32163 6004
rect 32197 5970 32231 6004
rect 32269 5970 32281 6004
rect 41277 6360 41311 6376
rect 41166 6332 41200 6342
rect 41166 6260 41200 6292
rect 41166 6190 41200 6224
rect 41166 6122 41200 6154
rect 41166 6072 41200 6082
rect 41277 6292 41311 6298
rect 41277 6224 41311 6226
rect 41277 6188 41311 6190
rect 41277 6116 41311 6122
rect 41277 6038 41311 6054
rect 41363 6360 41397 6376
rect 41363 6292 41397 6298
rect 41363 6224 41397 6226
rect 41363 6188 41397 6190
rect 41363 6116 41397 6122
rect 41363 6038 41397 6054
rect 41449 6360 41483 6376
rect 41449 6292 41483 6298
rect 41449 6224 41483 6226
rect 41449 6188 41483 6190
rect 41449 6116 41483 6122
rect 41560 6332 41594 6342
rect 41560 6260 41594 6292
rect 41560 6190 41594 6224
rect 41560 6122 41594 6154
rect 41560 6072 41594 6082
rect 41449 6038 41483 6054
rect 41279 5970 41291 6004
rect 41329 5970 41363 6004
rect 41397 5970 41431 6004
rect 41469 5970 41481 6004
rect 50477 6360 50511 6376
rect 50366 6332 50400 6342
rect 50366 6260 50400 6292
rect 50366 6190 50400 6224
rect 50366 6122 50400 6154
rect 50366 6072 50400 6082
rect 50477 6292 50511 6298
rect 50477 6224 50511 6226
rect 50477 6188 50511 6190
rect 50477 6116 50511 6122
rect 50477 6038 50511 6054
rect 50563 6360 50597 6376
rect 50563 6292 50597 6298
rect 50563 6224 50597 6226
rect 50563 6188 50597 6190
rect 50563 6116 50597 6122
rect 50563 6038 50597 6054
rect 50649 6360 50683 6376
rect 50649 6292 50683 6298
rect 50649 6224 50683 6226
rect 50649 6188 50683 6190
rect 50649 6116 50683 6122
rect 50760 6332 50794 6342
rect 50760 6260 50794 6292
rect 50760 6190 50794 6224
rect 50760 6122 50794 6154
rect 50760 6072 50794 6082
rect 50649 6038 50683 6054
rect 50479 5970 50491 6004
rect 50529 5970 50563 6004
rect 50597 5970 50631 6004
rect 50669 5970 50681 6004
rect 59677 6360 59711 6376
rect 59566 6332 59600 6342
rect 59566 6260 59600 6292
rect 59566 6190 59600 6224
rect 59566 6122 59600 6154
rect 59566 6072 59600 6082
rect 59677 6292 59711 6298
rect 59677 6224 59711 6226
rect 59677 6188 59711 6190
rect 59677 6116 59711 6122
rect 59677 6038 59711 6054
rect 59763 6360 59797 6376
rect 59763 6292 59797 6298
rect 59763 6224 59797 6226
rect 59763 6188 59797 6190
rect 59763 6116 59797 6122
rect 59763 6038 59797 6054
rect 59849 6360 59883 6376
rect 59849 6292 59883 6298
rect 59849 6224 59883 6226
rect 59849 6188 59883 6190
rect 59849 6116 59883 6122
rect 59960 6332 59994 6342
rect 59960 6260 59994 6292
rect 59960 6190 59994 6224
rect 59960 6122 59994 6154
rect 59960 6072 59994 6082
rect 59849 6038 59883 6054
rect 59679 5970 59691 6004
rect 59729 5970 59763 6004
rect 59797 5970 59831 6004
rect 59869 5970 59881 6004
rect 68877 6360 68911 6376
rect 68766 6332 68800 6342
rect 68766 6260 68800 6292
rect 68766 6190 68800 6224
rect 68766 6122 68800 6154
rect 68766 6072 68800 6082
rect 68877 6292 68911 6298
rect 68877 6224 68911 6226
rect 68877 6188 68911 6190
rect 68877 6116 68911 6122
rect 68877 6038 68911 6054
rect 68963 6360 68997 6376
rect 68963 6292 68997 6298
rect 68963 6224 68997 6226
rect 68963 6188 68997 6190
rect 68963 6116 68997 6122
rect 68963 6038 68997 6054
rect 69049 6360 69083 6376
rect 69049 6292 69083 6298
rect 69049 6224 69083 6226
rect 69049 6188 69083 6190
rect 69049 6116 69083 6122
rect 69160 6332 69194 6342
rect 69160 6260 69194 6292
rect 69160 6190 69194 6224
rect 69160 6122 69194 6154
rect 69160 6072 69194 6082
rect 69049 6038 69083 6054
rect 68879 5970 68891 6004
rect 68929 5970 68963 6004
rect 68997 5970 69031 6004
rect 69069 5970 69081 6004
rect -336 5872 -302 5888
rect -508 5830 -390 5832
rect -560 5800 -390 5830
rect -610 5792 -390 5800
rect -610 5790 -490 5792
rect -424 5734 -390 5792
rect -240 5820 -160 5840
rect -240 5780 -220 5820
rect -180 5780 -160 5820
rect -240 5760 -160 5780
rect -424 5442 -390 5458
rect -336 5734 -302 5750
rect -336 5378 -302 5458
rect -506 5370 -218 5378
rect -506 5320 -440 5370
rect -390 5356 -330 5370
rect -390 5320 -338 5356
rect -280 5320 -218 5370
rect -506 5300 -218 5320
<< viali >>
rect -480 95490 -440 95530
rect -400 95494 -392 95530
rect -392 95494 -360 95530
rect -310 95494 -278 95530
rect -278 95494 -270 95530
rect -400 95490 -360 95494
rect -310 95490 -270 95494
rect 4192 95535 4230 95932
rect 4930 95535 4968 95932
rect -424 94808 -390 95384
rect -600 94720 -560 94760
rect -336 94808 -302 95384
rect 4491 95330 4495 95364
rect 4495 95330 4525 95364
rect 4563 95330 4597 95364
rect 4635 95330 4665 95364
rect 4665 95330 4669 95364
rect 4192 94904 4230 95301
rect 4366 95246 4400 95252
rect 4366 95218 4400 95246
rect 4366 95178 4400 95180
rect 4366 95146 4400 95178
rect 4366 95076 4400 95108
rect 4366 95074 4400 95076
rect 4366 95008 4400 95036
rect 4366 95002 4400 95008
rect 4477 95246 4511 95252
rect 4477 95218 4511 95246
rect 4477 95178 4511 95180
rect 4477 95146 4511 95178
rect 4477 95076 4511 95108
rect 4477 95074 4511 95076
rect 4477 95008 4511 95036
rect 4477 95002 4511 95008
rect 4563 95246 4597 95252
rect 4563 95218 4597 95246
rect 4563 95178 4597 95180
rect 4563 95146 4597 95178
rect 4563 95076 4597 95108
rect 4563 95074 4597 95076
rect 4563 95008 4597 95036
rect 4563 95002 4597 95008
rect 4649 95246 4683 95252
rect 4649 95218 4683 95246
rect 4649 95178 4683 95180
rect 4649 95146 4683 95178
rect 4649 95076 4683 95108
rect 4649 95074 4683 95076
rect 4649 95008 4683 95036
rect 4649 95002 4683 95008
rect 4760 95246 4794 95252
rect 4760 95218 4794 95246
rect 4760 95178 4794 95180
rect 4760 95146 4794 95178
rect 4760 95076 4794 95108
rect 4760 95074 4794 95076
rect 4760 95008 4794 95036
rect 4760 95002 4794 95008
rect 4491 94890 4495 94924
rect 4495 94890 4525 94924
rect 4563 94890 4597 94924
rect 4635 94890 4665 94924
rect 4665 94890 4669 94924
rect 4930 94904 4968 95301
rect -220 94700 -180 94740
rect -424 94378 -390 94654
rect -336 94378 -302 94654
rect -440 94276 -390 94290
rect -330 94276 -280 94290
rect -440 94240 -434 94276
rect -434 94240 -398 94276
rect -398 94240 -390 94276
rect -330 94240 -300 94276
rect -300 94240 -280 94276
rect -480 85610 -440 85650
rect -400 85614 -392 85650
rect -392 85614 -360 85650
rect -310 85614 -278 85650
rect -278 85614 -270 85650
rect -400 85610 -360 85614
rect -310 85610 -270 85614
rect 4192 85655 4230 86052
rect 4930 85655 4968 86052
rect 13392 85655 13430 86052
rect 14130 85655 14168 86052
rect -424 84928 -390 85504
rect -600 84840 -560 84880
rect -336 84928 -302 85504
rect 4491 85450 4495 85484
rect 4495 85450 4525 85484
rect 4563 85450 4597 85484
rect 4635 85450 4665 85484
rect 4665 85450 4669 85484
rect 13691 85450 13695 85484
rect 13695 85450 13725 85484
rect 13763 85450 13797 85484
rect 13835 85450 13865 85484
rect 13865 85450 13869 85484
rect 4192 85024 4230 85421
rect 4366 85366 4400 85372
rect 4366 85338 4400 85366
rect 4366 85298 4400 85300
rect 4366 85266 4400 85298
rect 4366 85196 4400 85228
rect 4366 85194 4400 85196
rect 4366 85128 4400 85156
rect 4366 85122 4400 85128
rect 4477 85366 4511 85372
rect 4477 85338 4511 85366
rect 4477 85298 4511 85300
rect 4477 85266 4511 85298
rect 4477 85196 4511 85228
rect 4477 85194 4511 85196
rect 4477 85128 4511 85156
rect 4477 85122 4511 85128
rect 4563 85366 4597 85372
rect 4563 85338 4597 85366
rect 4563 85298 4597 85300
rect 4563 85266 4597 85298
rect 4563 85196 4597 85228
rect 4563 85194 4597 85196
rect 4563 85128 4597 85156
rect 4563 85122 4597 85128
rect 4649 85366 4683 85372
rect 4649 85338 4683 85366
rect 4649 85298 4683 85300
rect 4649 85266 4683 85298
rect 4649 85196 4683 85228
rect 4649 85194 4683 85196
rect 4649 85128 4683 85156
rect 4649 85122 4683 85128
rect 4760 85366 4794 85372
rect 4760 85338 4794 85366
rect 4760 85298 4794 85300
rect 4760 85266 4794 85298
rect 4760 85196 4794 85228
rect 4760 85194 4794 85196
rect 4760 85128 4794 85156
rect 4760 85122 4794 85128
rect 4491 85010 4495 85044
rect 4495 85010 4525 85044
rect 4563 85010 4597 85044
rect 4635 85010 4665 85044
rect 4665 85010 4669 85044
rect 4930 85024 4968 85421
rect 13392 85024 13430 85421
rect 13566 85366 13600 85372
rect 13566 85338 13600 85366
rect 13566 85298 13600 85300
rect 13566 85266 13600 85298
rect 13566 85196 13600 85228
rect 13566 85194 13600 85196
rect 13566 85128 13600 85156
rect 13566 85122 13600 85128
rect 13677 85366 13711 85372
rect 13677 85338 13711 85366
rect 13677 85298 13711 85300
rect 13677 85266 13711 85298
rect 13677 85196 13711 85228
rect 13677 85194 13711 85196
rect 13677 85128 13711 85156
rect 13677 85122 13711 85128
rect 13763 85366 13797 85372
rect 13763 85338 13797 85366
rect 13763 85298 13797 85300
rect 13763 85266 13797 85298
rect 13763 85196 13797 85228
rect 13763 85194 13797 85196
rect 13763 85128 13797 85156
rect 13763 85122 13797 85128
rect 13849 85366 13883 85372
rect 13849 85338 13883 85366
rect 13849 85298 13883 85300
rect 13849 85266 13883 85298
rect 13849 85196 13883 85228
rect 13849 85194 13883 85196
rect 13849 85128 13883 85156
rect 13849 85122 13883 85128
rect 13960 85366 13994 85372
rect 13960 85338 13994 85366
rect 13960 85298 13994 85300
rect 13960 85266 13994 85298
rect 13960 85196 13994 85228
rect 13960 85194 13994 85196
rect 13960 85128 13994 85156
rect 13960 85122 13994 85128
rect 13691 85010 13695 85044
rect 13695 85010 13725 85044
rect 13763 85010 13797 85044
rect 13835 85010 13865 85044
rect 13865 85010 13869 85044
rect 14130 85024 14168 85421
rect -220 84820 -180 84860
rect -424 84498 -390 84774
rect -336 84498 -302 84774
rect -440 84396 -390 84410
rect -330 84396 -280 84410
rect -440 84360 -434 84396
rect -434 84360 -398 84396
rect -398 84360 -390 84396
rect -330 84360 -300 84396
rect -300 84360 -280 84396
rect -480 75730 -440 75770
rect -400 75734 -392 75770
rect -392 75734 -360 75770
rect -310 75734 -278 75770
rect -278 75734 -270 75770
rect -400 75730 -360 75734
rect -310 75730 -270 75734
rect 4192 75775 4230 76172
rect 4930 75775 4968 76172
rect 13392 75775 13430 76172
rect 14130 75775 14168 76172
rect 22592 75775 22630 76172
rect 23330 75775 23368 76172
rect 31792 75775 31830 76172
rect 32530 75775 32568 76172
rect -424 75048 -390 75624
rect -600 74960 -560 75000
rect -336 75048 -302 75624
rect 4491 75570 4495 75604
rect 4495 75570 4525 75604
rect 4563 75570 4597 75604
rect 4635 75570 4665 75604
rect 4665 75570 4669 75604
rect 13691 75570 13695 75604
rect 13695 75570 13725 75604
rect 13763 75570 13797 75604
rect 13835 75570 13865 75604
rect 13865 75570 13869 75604
rect 22891 75570 22895 75604
rect 22895 75570 22925 75604
rect 22963 75570 22997 75604
rect 23035 75570 23065 75604
rect 23065 75570 23069 75604
rect 32091 75570 32095 75604
rect 32095 75570 32125 75604
rect 32163 75570 32197 75604
rect 32235 75570 32265 75604
rect 32265 75570 32269 75604
rect 4192 75144 4230 75541
rect 4366 75486 4400 75492
rect 4366 75458 4400 75486
rect 4366 75418 4400 75420
rect 4366 75386 4400 75418
rect 4366 75316 4400 75348
rect 4366 75314 4400 75316
rect 4366 75248 4400 75276
rect 4366 75242 4400 75248
rect 4477 75486 4511 75492
rect 4477 75458 4511 75486
rect 4477 75418 4511 75420
rect 4477 75386 4511 75418
rect 4477 75316 4511 75348
rect 4477 75314 4511 75316
rect 4477 75248 4511 75276
rect 4477 75242 4511 75248
rect 4563 75486 4597 75492
rect 4563 75458 4597 75486
rect 4563 75418 4597 75420
rect 4563 75386 4597 75418
rect 4563 75316 4597 75348
rect 4563 75314 4597 75316
rect 4563 75248 4597 75276
rect 4563 75242 4597 75248
rect 4649 75486 4683 75492
rect 4649 75458 4683 75486
rect 4649 75418 4683 75420
rect 4649 75386 4683 75418
rect 4649 75316 4683 75348
rect 4649 75314 4683 75316
rect 4649 75248 4683 75276
rect 4649 75242 4683 75248
rect 4760 75486 4794 75492
rect 4760 75458 4794 75486
rect 4760 75418 4794 75420
rect 4760 75386 4794 75418
rect 4760 75316 4794 75348
rect 4760 75314 4794 75316
rect 4760 75248 4794 75276
rect 4760 75242 4794 75248
rect 4491 75130 4495 75164
rect 4495 75130 4525 75164
rect 4563 75130 4597 75164
rect 4635 75130 4665 75164
rect 4665 75130 4669 75164
rect 4930 75144 4968 75541
rect 13392 75144 13430 75541
rect 13566 75486 13600 75492
rect 13566 75458 13600 75486
rect 13566 75418 13600 75420
rect 13566 75386 13600 75418
rect 13566 75316 13600 75348
rect 13566 75314 13600 75316
rect 13566 75248 13600 75276
rect 13566 75242 13600 75248
rect 13677 75486 13711 75492
rect 13677 75458 13711 75486
rect 13677 75418 13711 75420
rect 13677 75386 13711 75418
rect 13677 75316 13711 75348
rect 13677 75314 13711 75316
rect 13677 75248 13711 75276
rect 13677 75242 13711 75248
rect 13763 75486 13797 75492
rect 13763 75458 13797 75486
rect 13763 75418 13797 75420
rect 13763 75386 13797 75418
rect 13763 75316 13797 75348
rect 13763 75314 13797 75316
rect 13763 75248 13797 75276
rect 13763 75242 13797 75248
rect 13849 75486 13883 75492
rect 13849 75458 13883 75486
rect 13849 75418 13883 75420
rect 13849 75386 13883 75418
rect 13849 75316 13883 75348
rect 13849 75314 13883 75316
rect 13849 75248 13883 75276
rect 13849 75242 13883 75248
rect 13960 75486 13994 75492
rect 13960 75458 13994 75486
rect 13960 75418 13994 75420
rect 13960 75386 13994 75418
rect 13960 75316 13994 75348
rect 13960 75314 13994 75316
rect 13960 75248 13994 75276
rect 13960 75242 13994 75248
rect 13691 75130 13695 75164
rect 13695 75130 13725 75164
rect 13763 75130 13797 75164
rect 13835 75130 13865 75164
rect 13865 75130 13869 75164
rect 14130 75144 14168 75541
rect 22592 75144 22630 75541
rect 22766 75486 22800 75492
rect 22766 75458 22800 75486
rect 22766 75418 22800 75420
rect 22766 75386 22800 75418
rect 22766 75316 22800 75348
rect 22766 75314 22800 75316
rect 22766 75248 22800 75276
rect 22766 75242 22800 75248
rect 22877 75486 22911 75492
rect 22877 75458 22911 75486
rect 22877 75418 22911 75420
rect 22877 75386 22911 75418
rect 22877 75316 22911 75348
rect 22877 75314 22911 75316
rect 22877 75248 22911 75276
rect 22877 75242 22911 75248
rect 22963 75486 22997 75492
rect 22963 75458 22997 75486
rect 22963 75418 22997 75420
rect 22963 75386 22997 75418
rect 22963 75316 22997 75348
rect 22963 75314 22997 75316
rect 22963 75248 22997 75276
rect 22963 75242 22997 75248
rect 23049 75486 23083 75492
rect 23049 75458 23083 75486
rect 23049 75418 23083 75420
rect 23049 75386 23083 75418
rect 23049 75316 23083 75348
rect 23049 75314 23083 75316
rect 23049 75248 23083 75276
rect 23049 75242 23083 75248
rect 23160 75486 23194 75492
rect 23160 75458 23194 75486
rect 23160 75418 23194 75420
rect 23160 75386 23194 75418
rect 23160 75316 23194 75348
rect 23160 75314 23194 75316
rect 23160 75248 23194 75276
rect 23160 75242 23194 75248
rect 22891 75130 22895 75164
rect 22895 75130 22925 75164
rect 22963 75130 22997 75164
rect 23035 75130 23065 75164
rect 23065 75130 23069 75164
rect 23330 75144 23368 75541
rect 31792 75144 31830 75541
rect 31966 75486 32000 75492
rect 31966 75458 32000 75486
rect 31966 75418 32000 75420
rect 31966 75386 32000 75418
rect 31966 75316 32000 75348
rect 31966 75314 32000 75316
rect 31966 75248 32000 75276
rect 31966 75242 32000 75248
rect 32077 75486 32111 75492
rect 32077 75458 32111 75486
rect 32077 75418 32111 75420
rect 32077 75386 32111 75418
rect 32077 75316 32111 75348
rect 32077 75314 32111 75316
rect 32077 75248 32111 75276
rect 32077 75242 32111 75248
rect 32163 75486 32197 75492
rect 32163 75458 32197 75486
rect 32163 75418 32197 75420
rect 32163 75386 32197 75418
rect 32163 75316 32197 75348
rect 32163 75314 32197 75316
rect 32163 75248 32197 75276
rect 32163 75242 32197 75248
rect 32249 75486 32283 75492
rect 32249 75458 32283 75486
rect 32249 75418 32283 75420
rect 32249 75386 32283 75418
rect 32249 75316 32283 75348
rect 32249 75314 32283 75316
rect 32249 75248 32283 75276
rect 32249 75242 32283 75248
rect 32360 75486 32394 75492
rect 32360 75458 32394 75486
rect 32360 75418 32394 75420
rect 32360 75386 32394 75418
rect 32360 75316 32394 75348
rect 32360 75314 32394 75316
rect 32360 75248 32394 75276
rect 32360 75242 32394 75248
rect 32091 75130 32095 75164
rect 32095 75130 32125 75164
rect 32163 75130 32197 75164
rect 32235 75130 32265 75164
rect 32265 75130 32269 75164
rect 32530 75144 32568 75541
rect -220 74940 -180 74980
rect -424 74618 -390 74894
rect -336 74618 -302 74894
rect -440 74516 -390 74530
rect -330 74516 -280 74530
rect -440 74480 -434 74516
rect -434 74480 -398 74516
rect -398 74480 -390 74516
rect -330 74480 -300 74516
rect -300 74480 -280 74516
rect -480 65850 -440 65890
rect -400 65854 -392 65890
rect -392 65854 -360 65890
rect -310 65854 -278 65890
rect -278 65854 -270 65890
rect -400 65850 -360 65854
rect -310 65850 -270 65854
rect 4192 65895 4230 66292
rect 4930 65895 4968 66292
rect 13392 65895 13430 66292
rect 14130 65895 14168 66292
rect 22592 65895 22630 66292
rect 23330 65895 23368 66292
rect 31792 65895 31830 66292
rect 32530 65895 32568 66292
rect 40992 65895 41030 66292
rect 41730 65895 41768 66292
rect 50192 65895 50230 66292
rect 50930 65895 50968 66292
rect 59392 65895 59430 66292
rect 60130 65895 60168 66292
rect 68592 65895 68630 66292
rect 69330 65895 69368 66292
rect -424 65168 -390 65744
rect -600 65080 -560 65120
rect -336 65168 -302 65744
rect 4491 65690 4495 65724
rect 4495 65690 4525 65724
rect 4563 65690 4597 65724
rect 4635 65690 4665 65724
rect 4665 65690 4669 65724
rect 13691 65690 13695 65724
rect 13695 65690 13725 65724
rect 13763 65690 13797 65724
rect 13835 65690 13865 65724
rect 13865 65690 13869 65724
rect 22891 65690 22895 65724
rect 22895 65690 22925 65724
rect 22963 65690 22997 65724
rect 23035 65690 23065 65724
rect 23065 65690 23069 65724
rect 32091 65690 32095 65724
rect 32095 65690 32125 65724
rect 32163 65690 32197 65724
rect 32235 65690 32265 65724
rect 32265 65690 32269 65724
rect 41291 65690 41295 65724
rect 41295 65690 41325 65724
rect 41363 65690 41397 65724
rect 41435 65690 41465 65724
rect 41465 65690 41469 65724
rect 50491 65690 50495 65724
rect 50495 65690 50525 65724
rect 50563 65690 50597 65724
rect 50635 65690 50665 65724
rect 50665 65690 50669 65724
rect 59691 65690 59695 65724
rect 59695 65690 59725 65724
rect 59763 65690 59797 65724
rect 59835 65690 59865 65724
rect 59865 65690 59869 65724
rect 68891 65690 68895 65724
rect 68895 65690 68925 65724
rect 68963 65690 68997 65724
rect 69035 65690 69065 65724
rect 69065 65690 69069 65724
rect 4192 65264 4230 65661
rect 4366 65606 4400 65612
rect 4366 65578 4400 65606
rect 4366 65538 4400 65540
rect 4366 65506 4400 65538
rect 4366 65436 4400 65468
rect 4366 65434 4400 65436
rect 4366 65368 4400 65396
rect 4366 65362 4400 65368
rect 4477 65606 4511 65612
rect 4477 65578 4511 65606
rect 4477 65538 4511 65540
rect 4477 65506 4511 65538
rect 4477 65436 4511 65468
rect 4477 65434 4511 65436
rect 4477 65368 4511 65396
rect 4477 65362 4511 65368
rect 4563 65606 4597 65612
rect 4563 65578 4597 65606
rect 4563 65538 4597 65540
rect 4563 65506 4597 65538
rect 4563 65436 4597 65468
rect 4563 65434 4597 65436
rect 4563 65368 4597 65396
rect 4563 65362 4597 65368
rect 4649 65606 4683 65612
rect 4649 65578 4683 65606
rect 4649 65538 4683 65540
rect 4649 65506 4683 65538
rect 4649 65436 4683 65468
rect 4649 65434 4683 65436
rect 4649 65368 4683 65396
rect 4649 65362 4683 65368
rect 4760 65606 4794 65612
rect 4760 65578 4794 65606
rect 4760 65538 4794 65540
rect 4760 65506 4794 65538
rect 4760 65436 4794 65468
rect 4760 65434 4794 65436
rect 4760 65368 4794 65396
rect 4760 65362 4794 65368
rect 4491 65250 4495 65284
rect 4495 65250 4525 65284
rect 4563 65250 4597 65284
rect 4635 65250 4665 65284
rect 4665 65250 4669 65284
rect 4930 65264 4968 65661
rect 13392 65264 13430 65661
rect 13566 65606 13600 65612
rect 13566 65578 13600 65606
rect 13566 65538 13600 65540
rect 13566 65506 13600 65538
rect 13566 65436 13600 65468
rect 13566 65434 13600 65436
rect 13566 65368 13600 65396
rect 13566 65362 13600 65368
rect 13677 65606 13711 65612
rect 13677 65578 13711 65606
rect 13677 65538 13711 65540
rect 13677 65506 13711 65538
rect 13677 65436 13711 65468
rect 13677 65434 13711 65436
rect 13677 65368 13711 65396
rect 13677 65362 13711 65368
rect 13763 65606 13797 65612
rect 13763 65578 13797 65606
rect 13763 65538 13797 65540
rect 13763 65506 13797 65538
rect 13763 65436 13797 65468
rect 13763 65434 13797 65436
rect 13763 65368 13797 65396
rect 13763 65362 13797 65368
rect 13849 65606 13883 65612
rect 13849 65578 13883 65606
rect 13849 65538 13883 65540
rect 13849 65506 13883 65538
rect 13849 65436 13883 65468
rect 13849 65434 13883 65436
rect 13849 65368 13883 65396
rect 13849 65362 13883 65368
rect 13960 65606 13994 65612
rect 13960 65578 13994 65606
rect 13960 65538 13994 65540
rect 13960 65506 13994 65538
rect 13960 65436 13994 65468
rect 13960 65434 13994 65436
rect 13960 65368 13994 65396
rect 13960 65362 13994 65368
rect 13691 65250 13695 65284
rect 13695 65250 13725 65284
rect 13763 65250 13797 65284
rect 13835 65250 13865 65284
rect 13865 65250 13869 65284
rect 14130 65264 14168 65661
rect 22592 65264 22630 65661
rect 22766 65606 22800 65612
rect 22766 65578 22800 65606
rect 22766 65538 22800 65540
rect 22766 65506 22800 65538
rect 22766 65436 22800 65468
rect 22766 65434 22800 65436
rect 22766 65368 22800 65396
rect 22766 65362 22800 65368
rect 22877 65606 22911 65612
rect 22877 65578 22911 65606
rect 22877 65538 22911 65540
rect 22877 65506 22911 65538
rect 22877 65436 22911 65468
rect 22877 65434 22911 65436
rect 22877 65368 22911 65396
rect 22877 65362 22911 65368
rect 22963 65606 22997 65612
rect 22963 65578 22997 65606
rect 22963 65538 22997 65540
rect 22963 65506 22997 65538
rect 22963 65436 22997 65468
rect 22963 65434 22997 65436
rect 22963 65368 22997 65396
rect 22963 65362 22997 65368
rect 23049 65606 23083 65612
rect 23049 65578 23083 65606
rect 23049 65538 23083 65540
rect 23049 65506 23083 65538
rect 23049 65436 23083 65468
rect 23049 65434 23083 65436
rect 23049 65368 23083 65396
rect 23049 65362 23083 65368
rect 23160 65606 23194 65612
rect 23160 65578 23194 65606
rect 23160 65538 23194 65540
rect 23160 65506 23194 65538
rect 23160 65436 23194 65468
rect 23160 65434 23194 65436
rect 23160 65368 23194 65396
rect 23160 65362 23194 65368
rect 22891 65250 22895 65284
rect 22895 65250 22925 65284
rect 22963 65250 22997 65284
rect 23035 65250 23065 65284
rect 23065 65250 23069 65284
rect 23330 65264 23368 65661
rect 31792 65264 31830 65661
rect 31966 65606 32000 65612
rect 31966 65578 32000 65606
rect 31966 65538 32000 65540
rect 31966 65506 32000 65538
rect 31966 65436 32000 65468
rect 31966 65434 32000 65436
rect 31966 65368 32000 65396
rect 31966 65362 32000 65368
rect 32077 65606 32111 65612
rect 32077 65578 32111 65606
rect 32077 65538 32111 65540
rect 32077 65506 32111 65538
rect 32077 65436 32111 65468
rect 32077 65434 32111 65436
rect 32077 65368 32111 65396
rect 32077 65362 32111 65368
rect 32163 65606 32197 65612
rect 32163 65578 32197 65606
rect 32163 65538 32197 65540
rect 32163 65506 32197 65538
rect 32163 65436 32197 65468
rect 32163 65434 32197 65436
rect 32163 65368 32197 65396
rect 32163 65362 32197 65368
rect 32249 65606 32283 65612
rect 32249 65578 32283 65606
rect 32249 65538 32283 65540
rect 32249 65506 32283 65538
rect 32249 65436 32283 65468
rect 32249 65434 32283 65436
rect 32249 65368 32283 65396
rect 32249 65362 32283 65368
rect 32360 65606 32394 65612
rect 32360 65578 32394 65606
rect 32360 65538 32394 65540
rect 32360 65506 32394 65538
rect 32360 65436 32394 65468
rect 32360 65434 32394 65436
rect 32360 65368 32394 65396
rect 32360 65362 32394 65368
rect 32091 65250 32095 65284
rect 32095 65250 32125 65284
rect 32163 65250 32197 65284
rect 32235 65250 32265 65284
rect 32265 65250 32269 65284
rect 32530 65264 32568 65661
rect 40992 65264 41030 65661
rect 41166 65606 41200 65612
rect 41166 65578 41200 65606
rect 41166 65538 41200 65540
rect 41166 65506 41200 65538
rect 41166 65436 41200 65468
rect 41166 65434 41200 65436
rect 41166 65368 41200 65396
rect 41166 65362 41200 65368
rect 41277 65606 41311 65612
rect 41277 65578 41311 65606
rect 41277 65538 41311 65540
rect 41277 65506 41311 65538
rect 41277 65436 41311 65468
rect 41277 65434 41311 65436
rect 41277 65368 41311 65396
rect 41277 65362 41311 65368
rect 41363 65606 41397 65612
rect 41363 65578 41397 65606
rect 41363 65538 41397 65540
rect 41363 65506 41397 65538
rect 41363 65436 41397 65468
rect 41363 65434 41397 65436
rect 41363 65368 41397 65396
rect 41363 65362 41397 65368
rect 41449 65606 41483 65612
rect 41449 65578 41483 65606
rect 41449 65538 41483 65540
rect 41449 65506 41483 65538
rect 41449 65436 41483 65468
rect 41449 65434 41483 65436
rect 41449 65368 41483 65396
rect 41449 65362 41483 65368
rect 41560 65606 41594 65612
rect 41560 65578 41594 65606
rect 41560 65538 41594 65540
rect 41560 65506 41594 65538
rect 41560 65436 41594 65468
rect 41560 65434 41594 65436
rect 41560 65368 41594 65396
rect 41560 65362 41594 65368
rect 41291 65250 41295 65284
rect 41295 65250 41325 65284
rect 41363 65250 41397 65284
rect 41435 65250 41465 65284
rect 41465 65250 41469 65284
rect 41730 65264 41768 65661
rect 50192 65264 50230 65661
rect 50366 65606 50400 65612
rect 50366 65578 50400 65606
rect 50366 65538 50400 65540
rect 50366 65506 50400 65538
rect 50366 65436 50400 65468
rect 50366 65434 50400 65436
rect 50366 65368 50400 65396
rect 50366 65362 50400 65368
rect 50477 65606 50511 65612
rect 50477 65578 50511 65606
rect 50477 65538 50511 65540
rect 50477 65506 50511 65538
rect 50477 65436 50511 65468
rect 50477 65434 50511 65436
rect 50477 65368 50511 65396
rect 50477 65362 50511 65368
rect 50563 65606 50597 65612
rect 50563 65578 50597 65606
rect 50563 65538 50597 65540
rect 50563 65506 50597 65538
rect 50563 65436 50597 65468
rect 50563 65434 50597 65436
rect 50563 65368 50597 65396
rect 50563 65362 50597 65368
rect 50649 65606 50683 65612
rect 50649 65578 50683 65606
rect 50649 65538 50683 65540
rect 50649 65506 50683 65538
rect 50649 65436 50683 65468
rect 50649 65434 50683 65436
rect 50649 65368 50683 65396
rect 50649 65362 50683 65368
rect 50760 65606 50794 65612
rect 50760 65578 50794 65606
rect 50760 65538 50794 65540
rect 50760 65506 50794 65538
rect 50760 65436 50794 65468
rect 50760 65434 50794 65436
rect 50760 65368 50794 65396
rect 50760 65362 50794 65368
rect 50491 65250 50495 65284
rect 50495 65250 50525 65284
rect 50563 65250 50597 65284
rect 50635 65250 50665 65284
rect 50665 65250 50669 65284
rect 50930 65264 50968 65661
rect 59392 65264 59430 65661
rect 59566 65606 59600 65612
rect 59566 65578 59600 65606
rect 59566 65538 59600 65540
rect 59566 65506 59600 65538
rect 59566 65436 59600 65468
rect 59566 65434 59600 65436
rect 59566 65368 59600 65396
rect 59566 65362 59600 65368
rect 59677 65606 59711 65612
rect 59677 65578 59711 65606
rect 59677 65538 59711 65540
rect 59677 65506 59711 65538
rect 59677 65436 59711 65468
rect 59677 65434 59711 65436
rect 59677 65368 59711 65396
rect 59677 65362 59711 65368
rect 59763 65606 59797 65612
rect 59763 65578 59797 65606
rect 59763 65538 59797 65540
rect 59763 65506 59797 65538
rect 59763 65436 59797 65468
rect 59763 65434 59797 65436
rect 59763 65368 59797 65396
rect 59763 65362 59797 65368
rect 59849 65606 59883 65612
rect 59849 65578 59883 65606
rect 59849 65538 59883 65540
rect 59849 65506 59883 65538
rect 59849 65436 59883 65468
rect 59849 65434 59883 65436
rect 59849 65368 59883 65396
rect 59849 65362 59883 65368
rect 59960 65606 59994 65612
rect 59960 65578 59994 65606
rect 59960 65538 59994 65540
rect 59960 65506 59994 65538
rect 59960 65436 59994 65468
rect 59960 65434 59994 65436
rect 59960 65368 59994 65396
rect 59960 65362 59994 65368
rect 59691 65250 59695 65284
rect 59695 65250 59725 65284
rect 59763 65250 59797 65284
rect 59835 65250 59865 65284
rect 59865 65250 59869 65284
rect 60130 65264 60168 65661
rect 68592 65264 68630 65661
rect 68766 65606 68800 65612
rect 68766 65578 68800 65606
rect 68766 65538 68800 65540
rect 68766 65506 68800 65538
rect 68766 65436 68800 65468
rect 68766 65434 68800 65436
rect 68766 65368 68800 65396
rect 68766 65362 68800 65368
rect 68877 65606 68911 65612
rect 68877 65578 68911 65606
rect 68877 65538 68911 65540
rect 68877 65506 68911 65538
rect 68877 65436 68911 65468
rect 68877 65434 68911 65436
rect 68877 65368 68911 65396
rect 68877 65362 68911 65368
rect 68963 65606 68997 65612
rect 68963 65578 68997 65606
rect 68963 65538 68997 65540
rect 68963 65506 68997 65538
rect 68963 65436 68997 65468
rect 68963 65434 68997 65436
rect 68963 65368 68997 65396
rect 68963 65362 68997 65368
rect 69049 65606 69083 65612
rect 69049 65578 69083 65606
rect 69049 65538 69083 65540
rect 69049 65506 69083 65538
rect 69049 65436 69083 65468
rect 69049 65434 69083 65436
rect 69049 65368 69083 65396
rect 69049 65362 69083 65368
rect 69160 65606 69194 65612
rect 69160 65578 69194 65606
rect 69160 65538 69194 65540
rect 69160 65506 69194 65538
rect 69160 65436 69194 65468
rect 69160 65434 69194 65436
rect 69160 65368 69194 65396
rect 69160 65362 69194 65368
rect 68891 65250 68895 65284
rect 68895 65250 68925 65284
rect 68963 65250 68997 65284
rect 69035 65250 69065 65284
rect 69065 65250 69069 65284
rect 69330 65264 69368 65661
rect -220 65060 -180 65100
rect -424 64738 -390 65014
rect -336 64738 -302 65014
rect -440 64636 -390 64650
rect -330 64636 -280 64650
rect -440 64600 -434 64636
rect -434 64600 -398 64636
rect -398 64600 -390 64636
rect -330 64600 -300 64636
rect -300 64600 -280 64636
rect 4192 56015 4230 56412
rect 4930 56015 4968 56412
rect 13392 56015 13430 56412
rect 14130 56015 14168 56412
rect 22592 56015 22630 56412
rect 23330 56015 23368 56412
rect 31792 56015 31830 56412
rect 32530 56015 32568 56412
rect 40992 56015 41030 56412
rect 41730 56015 41768 56412
rect 50192 56015 50230 56412
rect 50930 56015 50968 56412
rect 59392 56015 59430 56412
rect 60130 56015 60168 56412
rect 68592 56015 68630 56412
rect 69330 56015 69368 56412
rect 4491 55810 4495 55844
rect 4495 55810 4525 55844
rect 4563 55810 4597 55844
rect 4635 55810 4665 55844
rect 4665 55810 4669 55844
rect 13691 55810 13695 55844
rect 13695 55810 13725 55844
rect 13763 55810 13797 55844
rect 13835 55810 13865 55844
rect 13865 55810 13869 55844
rect 22891 55810 22895 55844
rect 22895 55810 22925 55844
rect 22963 55810 22997 55844
rect 23035 55810 23065 55844
rect 23065 55810 23069 55844
rect 32091 55810 32095 55844
rect 32095 55810 32125 55844
rect 32163 55810 32197 55844
rect 32235 55810 32265 55844
rect 32265 55810 32269 55844
rect 41291 55810 41295 55844
rect 41295 55810 41325 55844
rect 41363 55810 41397 55844
rect 41435 55810 41465 55844
rect 41465 55810 41469 55844
rect 50491 55810 50495 55844
rect 50495 55810 50525 55844
rect 50563 55810 50597 55844
rect 50635 55810 50665 55844
rect 50665 55810 50669 55844
rect 59691 55810 59695 55844
rect 59695 55810 59725 55844
rect 59763 55810 59797 55844
rect 59835 55810 59865 55844
rect 59865 55810 59869 55844
rect 68891 55810 68895 55844
rect 68895 55810 68925 55844
rect 68963 55810 68997 55844
rect 69035 55810 69065 55844
rect 69065 55810 69069 55844
rect 4192 55384 4230 55781
rect 4366 55726 4400 55732
rect 4366 55698 4400 55726
rect 4366 55658 4400 55660
rect 4366 55626 4400 55658
rect 4366 55556 4400 55588
rect 4366 55554 4400 55556
rect 4366 55488 4400 55516
rect 4366 55482 4400 55488
rect 4477 55726 4511 55732
rect 4477 55698 4511 55726
rect 4477 55658 4511 55660
rect 4477 55626 4511 55658
rect 4477 55556 4511 55588
rect 4477 55554 4511 55556
rect 4477 55488 4511 55516
rect 4477 55482 4511 55488
rect 4563 55726 4597 55732
rect 4563 55698 4597 55726
rect 4563 55658 4597 55660
rect 4563 55626 4597 55658
rect 4563 55556 4597 55588
rect 4563 55554 4597 55556
rect 4563 55488 4597 55516
rect 4563 55482 4597 55488
rect 4649 55726 4683 55732
rect 4649 55698 4683 55726
rect 4649 55658 4683 55660
rect 4649 55626 4683 55658
rect 4649 55556 4683 55588
rect 4649 55554 4683 55556
rect 4649 55488 4683 55516
rect 4649 55482 4683 55488
rect 4760 55726 4794 55732
rect 4760 55698 4794 55726
rect 4760 55658 4794 55660
rect 4760 55626 4794 55658
rect 4760 55556 4794 55588
rect 4760 55554 4794 55556
rect 4760 55488 4794 55516
rect 4760 55482 4794 55488
rect 4491 55370 4495 55404
rect 4495 55370 4525 55404
rect 4563 55370 4597 55404
rect 4635 55370 4665 55404
rect 4665 55370 4669 55404
rect 4930 55384 4968 55781
rect 13392 55384 13430 55781
rect 13566 55726 13600 55732
rect 13566 55698 13600 55726
rect 13566 55658 13600 55660
rect 13566 55626 13600 55658
rect 13566 55556 13600 55588
rect 13566 55554 13600 55556
rect 13566 55488 13600 55516
rect 13566 55482 13600 55488
rect 13677 55726 13711 55732
rect 13677 55698 13711 55726
rect 13677 55658 13711 55660
rect 13677 55626 13711 55658
rect 13677 55556 13711 55588
rect 13677 55554 13711 55556
rect 13677 55488 13711 55516
rect 13677 55482 13711 55488
rect 13763 55726 13797 55732
rect 13763 55698 13797 55726
rect 13763 55658 13797 55660
rect 13763 55626 13797 55658
rect 13763 55556 13797 55588
rect 13763 55554 13797 55556
rect 13763 55488 13797 55516
rect 13763 55482 13797 55488
rect 13849 55726 13883 55732
rect 13849 55698 13883 55726
rect 13849 55658 13883 55660
rect 13849 55626 13883 55658
rect 13849 55556 13883 55588
rect 13849 55554 13883 55556
rect 13849 55488 13883 55516
rect 13849 55482 13883 55488
rect 13960 55726 13994 55732
rect 13960 55698 13994 55726
rect 13960 55658 13994 55660
rect 13960 55626 13994 55658
rect 13960 55556 13994 55588
rect 13960 55554 13994 55556
rect 13960 55488 13994 55516
rect 13960 55482 13994 55488
rect 13691 55370 13695 55404
rect 13695 55370 13725 55404
rect 13763 55370 13797 55404
rect 13835 55370 13865 55404
rect 13865 55370 13869 55404
rect 14130 55384 14168 55781
rect 22592 55384 22630 55781
rect 22766 55726 22800 55732
rect 22766 55698 22800 55726
rect 22766 55658 22800 55660
rect 22766 55626 22800 55658
rect 22766 55556 22800 55588
rect 22766 55554 22800 55556
rect 22766 55488 22800 55516
rect 22766 55482 22800 55488
rect 22877 55726 22911 55732
rect 22877 55698 22911 55726
rect 22877 55658 22911 55660
rect 22877 55626 22911 55658
rect 22877 55556 22911 55588
rect 22877 55554 22911 55556
rect 22877 55488 22911 55516
rect 22877 55482 22911 55488
rect 22963 55726 22997 55732
rect 22963 55698 22997 55726
rect 22963 55658 22997 55660
rect 22963 55626 22997 55658
rect 22963 55556 22997 55588
rect 22963 55554 22997 55556
rect 22963 55488 22997 55516
rect 22963 55482 22997 55488
rect 23049 55726 23083 55732
rect 23049 55698 23083 55726
rect 23049 55658 23083 55660
rect 23049 55626 23083 55658
rect 23049 55556 23083 55588
rect 23049 55554 23083 55556
rect 23049 55488 23083 55516
rect 23049 55482 23083 55488
rect 23160 55726 23194 55732
rect 23160 55698 23194 55726
rect 23160 55658 23194 55660
rect 23160 55626 23194 55658
rect 23160 55556 23194 55588
rect 23160 55554 23194 55556
rect 23160 55488 23194 55516
rect 23160 55482 23194 55488
rect 22891 55370 22895 55404
rect 22895 55370 22925 55404
rect 22963 55370 22997 55404
rect 23035 55370 23065 55404
rect 23065 55370 23069 55404
rect 23330 55384 23368 55781
rect 31792 55384 31830 55781
rect 31966 55726 32000 55732
rect 31966 55698 32000 55726
rect 31966 55658 32000 55660
rect 31966 55626 32000 55658
rect 31966 55556 32000 55588
rect 31966 55554 32000 55556
rect 31966 55488 32000 55516
rect 31966 55482 32000 55488
rect 32077 55726 32111 55732
rect 32077 55698 32111 55726
rect 32077 55658 32111 55660
rect 32077 55626 32111 55658
rect 32077 55556 32111 55588
rect 32077 55554 32111 55556
rect 32077 55488 32111 55516
rect 32077 55482 32111 55488
rect 32163 55726 32197 55732
rect 32163 55698 32197 55726
rect 32163 55658 32197 55660
rect 32163 55626 32197 55658
rect 32163 55556 32197 55588
rect 32163 55554 32197 55556
rect 32163 55488 32197 55516
rect 32163 55482 32197 55488
rect 32249 55726 32283 55732
rect 32249 55698 32283 55726
rect 32249 55658 32283 55660
rect 32249 55626 32283 55658
rect 32249 55556 32283 55588
rect 32249 55554 32283 55556
rect 32249 55488 32283 55516
rect 32249 55482 32283 55488
rect 32360 55726 32394 55732
rect 32360 55698 32394 55726
rect 32360 55658 32394 55660
rect 32360 55626 32394 55658
rect 32360 55556 32394 55588
rect 32360 55554 32394 55556
rect 32360 55488 32394 55516
rect 32360 55482 32394 55488
rect 32091 55370 32095 55404
rect 32095 55370 32125 55404
rect 32163 55370 32197 55404
rect 32235 55370 32265 55404
rect 32265 55370 32269 55404
rect 32530 55384 32568 55781
rect 40992 55384 41030 55781
rect 41166 55726 41200 55732
rect 41166 55698 41200 55726
rect 41166 55658 41200 55660
rect 41166 55626 41200 55658
rect 41166 55556 41200 55588
rect 41166 55554 41200 55556
rect 41166 55488 41200 55516
rect 41166 55482 41200 55488
rect 41277 55726 41311 55732
rect 41277 55698 41311 55726
rect 41277 55658 41311 55660
rect 41277 55626 41311 55658
rect 41277 55556 41311 55588
rect 41277 55554 41311 55556
rect 41277 55488 41311 55516
rect 41277 55482 41311 55488
rect 41363 55726 41397 55732
rect 41363 55698 41397 55726
rect 41363 55658 41397 55660
rect 41363 55626 41397 55658
rect 41363 55556 41397 55588
rect 41363 55554 41397 55556
rect 41363 55488 41397 55516
rect 41363 55482 41397 55488
rect 41449 55726 41483 55732
rect 41449 55698 41483 55726
rect 41449 55658 41483 55660
rect 41449 55626 41483 55658
rect 41449 55556 41483 55588
rect 41449 55554 41483 55556
rect 41449 55488 41483 55516
rect 41449 55482 41483 55488
rect 41560 55726 41594 55732
rect 41560 55698 41594 55726
rect 41560 55658 41594 55660
rect 41560 55626 41594 55658
rect 41560 55556 41594 55588
rect 41560 55554 41594 55556
rect 41560 55488 41594 55516
rect 41560 55482 41594 55488
rect 41291 55370 41295 55404
rect 41295 55370 41325 55404
rect 41363 55370 41397 55404
rect 41435 55370 41465 55404
rect 41465 55370 41469 55404
rect 41730 55384 41768 55781
rect 50192 55384 50230 55781
rect 50366 55726 50400 55732
rect 50366 55698 50400 55726
rect 50366 55658 50400 55660
rect 50366 55626 50400 55658
rect 50366 55556 50400 55588
rect 50366 55554 50400 55556
rect 50366 55488 50400 55516
rect 50366 55482 50400 55488
rect 50477 55726 50511 55732
rect 50477 55698 50511 55726
rect 50477 55658 50511 55660
rect 50477 55626 50511 55658
rect 50477 55556 50511 55588
rect 50477 55554 50511 55556
rect 50477 55488 50511 55516
rect 50477 55482 50511 55488
rect 50563 55726 50597 55732
rect 50563 55698 50597 55726
rect 50563 55658 50597 55660
rect 50563 55626 50597 55658
rect 50563 55556 50597 55588
rect 50563 55554 50597 55556
rect 50563 55488 50597 55516
rect 50563 55482 50597 55488
rect 50649 55726 50683 55732
rect 50649 55698 50683 55726
rect 50649 55658 50683 55660
rect 50649 55626 50683 55658
rect 50649 55556 50683 55588
rect 50649 55554 50683 55556
rect 50649 55488 50683 55516
rect 50649 55482 50683 55488
rect 50760 55726 50794 55732
rect 50760 55698 50794 55726
rect 50760 55658 50794 55660
rect 50760 55626 50794 55658
rect 50760 55556 50794 55588
rect 50760 55554 50794 55556
rect 50760 55488 50794 55516
rect 50760 55482 50794 55488
rect 50491 55370 50495 55404
rect 50495 55370 50525 55404
rect 50563 55370 50597 55404
rect 50635 55370 50665 55404
rect 50665 55370 50669 55404
rect 50930 55384 50968 55781
rect 59392 55384 59430 55781
rect 59566 55726 59600 55732
rect 59566 55698 59600 55726
rect 59566 55658 59600 55660
rect 59566 55626 59600 55658
rect 59566 55556 59600 55588
rect 59566 55554 59600 55556
rect 59566 55488 59600 55516
rect 59566 55482 59600 55488
rect 59677 55726 59711 55732
rect 59677 55698 59711 55726
rect 59677 55658 59711 55660
rect 59677 55626 59711 55658
rect 59677 55556 59711 55588
rect 59677 55554 59711 55556
rect 59677 55488 59711 55516
rect 59677 55482 59711 55488
rect 59763 55726 59797 55732
rect 59763 55698 59797 55726
rect 59763 55658 59797 55660
rect 59763 55626 59797 55658
rect 59763 55556 59797 55588
rect 59763 55554 59797 55556
rect 59763 55488 59797 55516
rect 59763 55482 59797 55488
rect 59849 55726 59883 55732
rect 59849 55698 59883 55726
rect 59849 55658 59883 55660
rect 59849 55626 59883 55658
rect 59849 55556 59883 55588
rect 59849 55554 59883 55556
rect 59849 55488 59883 55516
rect 59849 55482 59883 55488
rect 59960 55726 59994 55732
rect 59960 55698 59994 55726
rect 59960 55658 59994 55660
rect 59960 55626 59994 55658
rect 59960 55556 59994 55588
rect 59960 55554 59994 55556
rect 59960 55488 59994 55516
rect 59960 55482 59994 55488
rect 59691 55370 59695 55404
rect 59695 55370 59725 55404
rect 59763 55370 59797 55404
rect 59835 55370 59865 55404
rect 59865 55370 59869 55404
rect 60130 55384 60168 55781
rect 68592 55384 68630 55781
rect 68766 55726 68800 55732
rect 68766 55698 68800 55726
rect 68766 55658 68800 55660
rect 68766 55626 68800 55658
rect 68766 55556 68800 55588
rect 68766 55554 68800 55556
rect 68766 55488 68800 55516
rect 68766 55482 68800 55488
rect 68877 55726 68911 55732
rect 68877 55698 68911 55726
rect 68877 55658 68911 55660
rect 68877 55626 68911 55658
rect 68877 55556 68911 55588
rect 68877 55554 68911 55556
rect 68877 55488 68911 55516
rect 68877 55482 68911 55488
rect 68963 55726 68997 55732
rect 68963 55698 68997 55726
rect 68963 55658 68997 55660
rect 68963 55626 68997 55658
rect 68963 55556 68997 55588
rect 68963 55554 68997 55556
rect 68963 55488 68997 55516
rect 68963 55482 68997 55488
rect 69049 55726 69083 55732
rect 69049 55698 69083 55726
rect 69049 55658 69083 55660
rect 69049 55626 69083 55658
rect 69049 55556 69083 55588
rect 69049 55554 69083 55556
rect 69049 55488 69083 55516
rect 69049 55482 69083 55488
rect 69160 55726 69194 55732
rect 69160 55698 69194 55726
rect 69160 55658 69194 55660
rect 69160 55626 69194 55658
rect 69160 55556 69194 55588
rect 69160 55554 69194 55556
rect 69160 55488 69194 55516
rect 69160 55482 69194 55488
rect 68891 55370 68895 55404
rect 68895 55370 68925 55404
rect 68963 55370 68997 55404
rect 69035 55370 69065 55404
rect 69065 55370 69069 55404
rect 69330 55384 69368 55781
rect -480 46090 -440 46130
rect -400 46094 -392 46130
rect -392 46094 -360 46130
rect -310 46094 -278 46130
rect -278 46094 -270 46130
rect -400 46090 -360 46094
rect -310 46090 -270 46094
rect 4192 46135 4230 46532
rect 4930 46135 4968 46532
rect 13392 46135 13430 46532
rect 14130 46135 14168 46532
rect 22592 46135 22630 46532
rect 23330 46135 23368 46532
rect 31792 46135 31830 46532
rect 32530 46135 32568 46532
rect 40992 46135 41030 46532
rect 41730 46135 41768 46532
rect 50192 46135 50230 46532
rect 50930 46135 50968 46532
rect 59392 46135 59430 46532
rect 60130 46135 60168 46532
rect 68592 46135 68630 46532
rect 69330 46135 69368 46532
rect -424 45408 -390 45984
rect -600 45320 -560 45360
rect -336 45408 -302 45984
rect 4491 45930 4495 45964
rect 4495 45930 4525 45964
rect 4563 45930 4597 45964
rect 4635 45930 4665 45964
rect 4665 45930 4669 45964
rect 13691 45930 13695 45964
rect 13695 45930 13725 45964
rect 13763 45930 13797 45964
rect 13835 45930 13865 45964
rect 13865 45930 13869 45964
rect 22891 45930 22895 45964
rect 22895 45930 22925 45964
rect 22963 45930 22997 45964
rect 23035 45930 23065 45964
rect 23065 45930 23069 45964
rect 32091 45930 32095 45964
rect 32095 45930 32125 45964
rect 32163 45930 32197 45964
rect 32235 45930 32265 45964
rect 32265 45930 32269 45964
rect 41291 45930 41295 45964
rect 41295 45930 41325 45964
rect 41363 45930 41397 45964
rect 41435 45930 41465 45964
rect 41465 45930 41469 45964
rect 50491 45930 50495 45964
rect 50495 45930 50525 45964
rect 50563 45930 50597 45964
rect 50635 45930 50665 45964
rect 50665 45930 50669 45964
rect 59691 45930 59695 45964
rect 59695 45930 59725 45964
rect 59763 45930 59797 45964
rect 59835 45930 59865 45964
rect 59865 45930 59869 45964
rect 68891 45930 68895 45964
rect 68895 45930 68925 45964
rect 68963 45930 68997 45964
rect 69035 45930 69065 45964
rect 69065 45930 69069 45964
rect 4192 45504 4230 45901
rect 4366 45846 4400 45852
rect 4366 45818 4400 45846
rect 4366 45778 4400 45780
rect 4366 45746 4400 45778
rect 4366 45676 4400 45708
rect 4366 45674 4400 45676
rect 4366 45608 4400 45636
rect 4366 45602 4400 45608
rect 4477 45846 4511 45852
rect 4477 45818 4511 45846
rect 4477 45778 4511 45780
rect 4477 45746 4511 45778
rect 4477 45676 4511 45708
rect 4477 45674 4511 45676
rect 4477 45608 4511 45636
rect 4477 45602 4511 45608
rect 4563 45846 4597 45852
rect 4563 45818 4597 45846
rect 4563 45778 4597 45780
rect 4563 45746 4597 45778
rect 4563 45676 4597 45708
rect 4563 45674 4597 45676
rect 4563 45608 4597 45636
rect 4563 45602 4597 45608
rect 4649 45846 4683 45852
rect 4649 45818 4683 45846
rect 4649 45778 4683 45780
rect 4649 45746 4683 45778
rect 4649 45676 4683 45708
rect 4649 45674 4683 45676
rect 4649 45608 4683 45636
rect 4649 45602 4683 45608
rect 4760 45846 4794 45852
rect 4760 45818 4794 45846
rect 4760 45778 4794 45780
rect 4760 45746 4794 45778
rect 4760 45676 4794 45708
rect 4760 45674 4794 45676
rect 4760 45608 4794 45636
rect 4760 45602 4794 45608
rect 4491 45490 4495 45524
rect 4495 45490 4525 45524
rect 4563 45490 4597 45524
rect 4635 45490 4665 45524
rect 4665 45490 4669 45524
rect 4930 45504 4968 45901
rect 13392 45504 13430 45901
rect 13566 45846 13600 45852
rect 13566 45818 13600 45846
rect 13566 45778 13600 45780
rect 13566 45746 13600 45778
rect 13566 45676 13600 45708
rect 13566 45674 13600 45676
rect 13566 45608 13600 45636
rect 13566 45602 13600 45608
rect 13677 45846 13711 45852
rect 13677 45818 13711 45846
rect 13677 45778 13711 45780
rect 13677 45746 13711 45778
rect 13677 45676 13711 45708
rect 13677 45674 13711 45676
rect 13677 45608 13711 45636
rect 13677 45602 13711 45608
rect 13763 45846 13797 45852
rect 13763 45818 13797 45846
rect 13763 45778 13797 45780
rect 13763 45746 13797 45778
rect 13763 45676 13797 45708
rect 13763 45674 13797 45676
rect 13763 45608 13797 45636
rect 13763 45602 13797 45608
rect 13849 45846 13883 45852
rect 13849 45818 13883 45846
rect 13849 45778 13883 45780
rect 13849 45746 13883 45778
rect 13849 45676 13883 45708
rect 13849 45674 13883 45676
rect 13849 45608 13883 45636
rect 13849 45602 13883 45608
rect 13960 45846 13994 45852
rect 13960 45818 13994 45846
rect 13960 45778 13994 45780
rect 13960 45746 13994 45778
rect 13960 45676 13994 45708
rect 13960 45674 13994 45676
rect 13960 45608 13994 45636
rect 13960 45602 13994 45608
rect 13691 45490 13695 45524
rect 13695 45490 13725 45524
rect 13763 45490 13797 45524
rect 13835 45490 13865 45524
rect 13865 45490 13869 45524
rect 14130 45504 14168 45901
rect 22592 45504 22630 45901
rect 22766 45846 22800 45852
rect 22766 45818 22800 45846
rect 22766 45778 22800 45780
rect 22766 45746 22800 45778
rect 22766 45676 22800 45708
rect 22766 45674 22800 45676
rect 22766 45608 22800 45636
rect 22766 45602 22800 45608
rect 22877 45846 22911 45852
rect 22877 45818 22911 45846
rect 22877 45778 22911 45780
rect 22877 45746 22911 45778
rect 22877 45676 22911 45708
rect 22877 45674 22911 45676
rect 22877 45608 22911 45636
rect 22877 45602 22911 45608
rect 22963 45846 22997 45852
rect 22963 45818 22997 45846
rect 22963 45778 22997 45780
rect 22963 45746 22997 45778
rect 22963 45676 22997 45708
rect 22963 45674 22997 45676
rect 22963 45608 22997 45636
rect 22963 45602 22997 45608
rect 23049 45846 23083 45852
rect 23049 45818 23083 45846
rect 23049 45778 23083 45780
rect 23049 45746 23083 45778
rect 23049 45676 23083 45708
rect 23049 45674 23083 45676
rect 23049 45608 23083 45636
rect 23049 45602 23083 45608
rect 23160 45846 23194 45852
rect 23160 45818 23194 45846
rect 23160 45778 23194 45780
rect 23160 45746 23194 45778
rect 23160 45676 23194 45708
rect 23160 45674 23194 45676
rect 23160 45608 23194 45636
rect 23160 45602 23194 45608
rect 22891 45490 22895 45524
rect 22895 45490 22925 45524
rect 22963 45490 22997 45524
rect 23035 45490 23065 45524
rect 23065 45490 23069 45524
rect 23330 45504 23368 45901
rect 31792 45504 31830 45901
rect 31966 45846 32000 45852
rect 31966 45818 32000 45846
rect 31966 45778 32000 45780
rect 31966 45746 32000 45778
rect 31966 45676 32000 45708
rect 31966 45674 32000 45676
rect 31966 45608 32000 45636
rect 31966 45602 32000 45608
rect 32077 45846 32111 45852
rect 32077 45818 32111 45846
rect 32077 45778 32111 45780
rect 32077 45746 32111 45778
rect 32077 45676 32111 45708
rect 32077 45674 32111 45676
rect 32077 45608 32111 45636
rect 32077 45602 32111 45608
rect 32163 45846 32197 45852
rect 32163 45818 32197 45846
rect 32163 45778 32197 45780
rect 32163 45746 32197 45778
rect 32163 45676 32197 45708
rect 32163 45674 32197 45676
rect 32163 45608 32197 45636
rect 32163 45602 32197 45608
rect 32249 45846 32283 45852
rect 32249 45818 32283 45846
rect 32249 45778 32283 45780
rect 32249 45746 32283 45778
rect 32249 45676 32283 45708
rect 32249 45674 32283 45676
rect 32249 45608 32283 45636
rect 32249 45602 32283 45608
rect 32360 45846 32394 45852
rect 32360 45818 32394 45846
rect 32360 45778 32394 45780
rect 32360 45746 32394 45778
rect 32360 45676 32394 45708
rect 32360 45674 32394 45676
rect 32360 45608 32394 45636
rect 32360 45602 32394 45608
rect 32091 45490 32095 45524
rect 32095 45490 32125 45524
rect 32163 45490 32197 45524
rect 32235 45490 32265 45524
rect 32265 45490 32269 45524
rect 32530 45504 32568 45901
rect 40992 45504 41030 45901
rect 41166 45846 41200 45852
rect 41166 45818 41200 45846
rect 41166 45778 41200 45780
rect 41166 45746 41200 45778
rect 41166 45676 41200 45708
rect 41166 45674 41200 45676
rect 41166 45608 41200 45636
rect 41166 45602 41200 45608
rect 41277 45846 41311 45852
rect 41277 45818 41311 45846
rect 41277 45778 41311 45780
rect 41277 45746 41311 45778
rect 41277 45676 41311 45708
rect 41277 45674 41311 45676
rect 41277 45608 41311 45636
rect 41277 45602 41311 45608
rect 41363 45846 41397 45852
rect 41363 45818 41397 45846
rect 41363 45778 41397 45780
rect 41363 45746 41397 45778
rect 41363 45676 41397 45708
rect 41363 45674 41397 45676
rect 41363 45608 41397 45636
rect 41363 45602 41397 45608
rect 41449 45846 41483 45852
rect 41449 45818 41483 45846
rect 41449 45778 41483 45780
rect 41449 45746 41483 45778
rect 41449 45676 41483 45708
rect 41449 45674 41483 45676
rect 41449 45608 41483 45636
rect 41449 45602 41483 45608
rect 41560 45846 41594 45852
rect 41560 45818 41594 45846
rect 41560 45778 41594 45780
rect 41560 45746 41594 45778
rect 41560 45676 41594 45708
rect 41560 45674 41594 45676
rect 41560 45608 41594 45636
rect 41560 45602 41594 45608
rect 41291 45490 41295 45524
rect 41295 45490 41325 45524
rect 41363 45490 41397 45524
rect 41435 45490 41465 45524
rect 41465 45490 41469 45524
rect 41730 45504 41768 45901
rect 50192 45504 50230 45901
rect 50366 45846 50400 45852
rect 50366 45818 50400 45846
rect 50366 45778 50400 45780
rect 50366 45746 50400 45778
rect 50366 45676 50400 45708
rect 50366 45674 50400 45676
rect 50366 45608 50400 45636
rect 50366 45602 50400 45608
rect 50477 45846 50511 45852
rect 50477 45818 50511 45846
rect 50477 45778 50511 45780
rect 50477 45746 50511 45778
rect 50477 45676 50511 45708
rect 50477 45674 50511 45676
rect 50477 45608 50511 45636
rect 50477 45602 50511 45608
rect 50563 45846 50597 45852
rect 50563 45818 50597 45846
rect 50563 45778 50597 45780
rect 50563 45746 50597 45778
rect 50563 45676 50597 45708
rect 50563 45674 50597 45676
rect 50563 45608 50597 45636
rect 50563 45602 50597 45608
rect 50649 45846 50683 45852
rect 50649 45818 50683 45846
rect 50649 45778 50683 45780
rect 50649 45746 50683 45778
rect 50649 45676 50683 45708
rect 50649 45674 50683 45676
rect 50649 45608 50683 45636
rect 50649 45602 50683 45608
rect 50760 45846 50794 45852
rect 50760 45818 50794 45846
rect 50760 45778 50794 45780
rect 50760 45746 50794 45778
rect 50760 45676 50794 45708
rect 50760 45674 50794 45676
rect 50760 45608 50794 45636
rect 50760 45602 50794 45608
rect 50491 45490 50495 45524
rect 50495 45490 50525 45524
rect 50563 45490 50597 45524
rect 50635 45490 50665 45524
rect 50665 45490 50669 45524
rect 50930 45504 50968 45901
rect 59392 45504 59430 45901
rect 59566 45846 59600 45852
rect 59566 45818 59600 45846
rect 59566 45778 59600 45780
rect 59566 45746 59600 45778
rect 59566 45676 59600 45708
rect 59566 45674 59600 45676
rect 59566 45608 59600 45636
rect 59566 45602 59600 45608
rect 59677 45846 59711 45852
rect 59677 45818 59711 45846
rect 59677 45778 59711 45780
rect 59677 45746 59711 45778
rect 59677 45676 59711 45708
rect 59677 45674 59711 45676
rect 59677 45608 59711 45636
rect 59677 45602 59711 45608
rect 59763 45846 59797 45852
rect 59763 45818 59797 45846
rect 59763 45778 59797 45780
rect 59763 45746 59797 45778
rect 59763 45676 59797 45708
rect 59763 45674 59797 45676
rect 59763 45608 59797 45636
rect 59763 45602 59797 45608
rect 59849 45846 59883 45852
rect 59849 45818 59883 45846
rect 59849 45778 59883 45780
rect 59849 45746 59883 45778
rect 59849 45676 59883 45708
rect 59849 45674 59883 45676
rect 59849 45608 59883 45636
rect 59849 45602 59883 45608
rect 59960 45846 59994 45852
rect 59960 45818 59994 45846
rect 59960 45778 59994 45780
rect 59960 45746 59994 45778
rect 59960 45676 59994 45708
rect 59960 45674 59994 45676
rect 59960 45608 59994 45636
rect 59960 45602 59994 45608
rect 59691 45490 59695 45524
rect 59695 45490 59725 45524
rect 59763 45490 59797 45524
rect 59835 45490 59865 45524
rect 59865 45490 59869 45524
rect 60130 45504 60168 45901
rect 68592 45504 68630 45901
rect 68766 45846 68800 45852
rect 68766 45818 68800 45846
rect 68766 45778 68800 45780
rect 68766 45746 68800 45778
rect 68766 45676 68800 45708
rect 68766 45674 68800 45676
rect 68766 45608 68800 45636
rect 68766 45602 68800 45608
rect 68877 45846 68911 45852
rect 68877 45818 68911 45846
rect 68877 45778 68911 45780
rect 68877 45746 68911 45778
rect 68877 45676 68911 45708
rect 68877 45674 68911 45676
rect 68877 45608 68911 45636
rect 68877 45602 68911 45608
rect 68963 45846 68997 45852
rect 68963 45818 68997 45846
rect 68963 45778 68997 45780
rect 68963 45746 68997 45778
rect 68963 45676 68997 45708
rect 68963 45674 68997 45676
rect 68963 45608 68997 45636
rect 68963 45602 68997 45608
rect 69049 45846 69083 45852
rect 69049 45818 69083 45846
rect 69049 45778 69083 45780
rect 69049 45746 69083 45778
rect 69049 45676 69083 45708
rect 69049 45674 69083 45676
rect 69049 45608 69083 45636
rect 69049 45602 69083 45608
rect 69160 45846 69194 45852
rect 69160 45818 69194 45846
rect 69160 45778 69194 45780
rect 69160 45746 69194 45778
rect 69160 45676 69194 45708
rect 69160 45674 69194 45676
rect 69160 45608 69194 45636
rect 69160 45602 69194 45608
rect 68891 45490 68895 45524
rect 68895 45490 68925 45524
rect 68963 45490 68997 45524
rect 69035 45490 69065 45524
rect 69065 45490 69069 45524
rect 69330 45504 69368 45901
rect -220 45300 -180 45340
rect -424 44978 -390 45254
rect -336 44978 -302 45254
rect -440 44876 -390 44890
rect -330 44876 -280 44890
rect -440 44840 -434 44876
rect -434 44840 -398 44876
rect -398 44840 -390 44876
rect -330 44840 -300 44876
rect -300 44840 -280 44876
rect 4192 36255 4230 36652
rect 4930 36255 4968 36652
rect 13392 36255 13430 36652
rect 14130 36255 14168 36652
rect 22592 36255 22630 36652
rect 23330 36255 23368 36652
rect 31792 36255 31830 36652
rect 32530 36255 32568 36652
rect 40992 36255 41030 36652
rect 41730 36255 41768 36652
rect 50192 36255 50230 36652
rect 50930 36255 50968 36652
rect 59392 36255 59430 36652
rect 60130 36255 60168 36652
rect 68592 36255 68630 36652
rect 69330 36255 69368 36652
rect 4491 36050 4495 36084
rect 4495 36050 4525 36084
rect 4563 36050 4597 36084
rect 4635 36050 4665 36084
rect 4665 36050 4669 36084
rect 13691 36050 13695 36084
rect 13695 36050 13725 36084
rect 13763 36050 13797 36084
rect 13835 36050 13865 36084
rect 13865 36050 13869 36084
rect 22891 36050 22895 36084
rect 22895 36050 22925 36084
rect 22963 36050 22997 36084
rect 23035 36050 23065 36084
rect 23065 36050 23069 36084
rect 32091 36050 32095 36084
rect 32095 36050 32125 36084
rect 32163 36050 32197 36084
rect 32235 36050 32265 36084
rect 32265 36050 32269 36084
rect 41291 36050 41295 36084
rect 41295 36050 41325 36084
rect 41363 36050 41397 36084
rect 41435 36050 41465 36084
rect 41465 36050 41469 36084
rect 50491 36050 50495 36084
rect 50495 36050 50525 36084
rect 50563 36050 50597 36084
rect 50635 36050 50665 36084
rect 50665 36050 50669 36084
rect 59691 36050 59695 36084
rect 59695 36050 59725 36084
rect 59763 36050 59797 36084
rect 59835 36050 59865 36084
rect 59865 36050 59869 36084
rect 68891 36050 68895 36084
rect 68895 36050 68925 36084
rect 68963 36050 68997 36084
rect 69035 36050 69065 36084
rect 69065 36050 69069 36084
rect 4192 35624 4230 36021
rect 4366 35966 4400 35972
rect 4366 35938 4400 35966
rect 4366 35898 4400 35900
rect 4366 35866 4400 35898
rect 4366 35796 4400 35828
rect 4366 35794 4400 35796
rect 4366 35728 4400 35756
rect 4366 35722 4400 35728
rect 4477 35966 4511 35972
rect 4477 35938 4511 35966
rect 4477 35898 4511 35900
rect 4477 35866 4511 35898
rect 4477 35796 4511 35828
rect 4477 35794 4511 35796
rect 4477 35728 4511 35756
rect 4477 35722 4511 35728
rect 4563 35966 4597 35972
rect 4563 35938 4597 35966
rect 4563 35898 4597 35900
rect 4563 35866 4597 35898
rect 4563 35796 4597 35828
rect 4563 35794 4597 35796
rect 4563 35728 4597 35756
rect 4563 35722 4597 35728
rect 4649 35966 4683 35972
rect 4649 35938 4683 35966
rect 4649 35898 4683 35900
rect 4649 35866 4683 35898
rect 4649 35796 4683 35828
rect 4649 35794 4683 35796
rect 4649 35728 4683 35756
rect 4649 35722 4683 35728
rect 4760 35966 4794 35972
rect 4760 35938 4794 35966
rect 4760 35898 4794 35900
rect 4760 35866 4794 35898
rect 4760 35796 4794 35828
rect 4760 35794 4794 35796
rect 4760 35728 4794 35756
rect 4760 35722 4794 35728
rect 4491 35610 4495 35644
rect 4495 35610 4525 35644
rect 4563 35610 4597 35644
rect 4635 35610 4665 35644
rect 4665 35610 4669 35644
rect 4930 35624 4968 36021
rect 13392 35624 13430 36021
rect 13566 35966 13600 35972
rect 13566 35938 13600 35966
rect 13566 35898 13600 35900
rect 13566 35866 13600 35898
rect 13566 35796 13600 35828
rect 13566 35794 13600 35796
rect 13566 35728 13600 35756
rect 13566 35722 13600 35728
rect 13677 35966 13711 35972
rect 13677 35938 13711 35966
rect 13677 35898 13711 35900
rect 13677 35866 13711 35898
rect 13677 35796 13711 35828
rect 13677 35794 13711 35796
rect 13677 35728 13711 35756
rect 13677 35722 13711 35728
rect 13763 35966 13797 35972
rect 13763 35938 13797 35966
rect 13763 35898 13797 35900
rect 13763 35866 13797 35898
rect 13763 35796 13797 35828
rect 13763 35794 13797 35796
rect 13763 35728 13797 35756
rect 13763 35722 13797 35728
rect 13849 35966 13883 35972
rect 13849 35938 13883 35966
rect 13849 35898 13883 35900
rect 13849 35866 13883 35898
rect 13849 35796 13883 35828
rect 13849 35794 13883 35796
rect 13849 35728 13883 35756
rect 13849 35722 13883 35728
rect 13960 35966 13994 35972
rect 13960 35938 13994 35966
rect 13960 35898 13994 35900
rect 13960 35866 13994 35898
rect 13960 35796 13994 35828
rect 13960 35794 13994 35796
rect 13960 35728 13994 35756
rect 13960 35722 13994 35728
rect 13691 35610 13695 35644
rect 13695 35610 13725 35644
rect 13763 35610 13797 35644
rect 13835 35610 13865 35644
rect 13865 35610 13869 35644
rect 14130 35624 14168 36021
rect 22592 35624 22630 36021
rect 22766 35966 22800 35972
rect 22766 35938 22800 35966
rect 22766 35898 22800 35900
rect 22766 35866 22800 35898
rect 22766 35796 22800 35828
rect 22766 35794 22800 35796
rect 22766 35728 22800 35756
rect 22766 35722 22800 35728
rect 22877 35966 22911 35972
rect 22877 35938 22911 35966
rect 22877 35898 22911 35900
rect 22877 35866 22911 35898
rect 22877 35796 22911 35828
rect 22877 35794 22911 35796
rect 22877 35728 22911 35756
rect 22877 35722 22911 35728
rect 22963 35966 22997 35972
rect 22963 35938 22997 35966
rect 22963 35898 22997 35900
rect 22963 35866 22997 35898
rect 22963 35796 22997 35828
rect 22963 35794 22997 35796
rect 22963 35728 22997 35756
rect 22963 35722 22997 35728
rect 23049 35966 23083 35972
rect 23049 35938 23083 35966
rect 23049 35898 23083 35900
rect 23049 35866 23083 35898
rect 23049 35796 23083 35828
rect 23049 35794 23083 35796
rect 23049 35728 23083 35756
rect 23049 35722 23083 35728
rect 23160 35966 23194 35972
rect 23160 35938 23194 35966
rect 23160 35898 23194 35900
rect 23160 35866 23194 35898
rect 23160 35796 23194 35828
rect 23160 35794 23194 35796
rect 23160 35728 23194 35756
rect 23160 35722 23194 35728
rect 22891 35610 22895 35644
rect 22895 35610 22925 35644
rect 22963 35610 22997 35644
rect 23035 35610 23065 35644
rect 23065 35610 23069 35644
rect 23330 35624 23368 36021
rect 31792 35624 31830 36021
rect 31966 35966 32000 35972
rect 31966 35938 32000 35966
rect 31966 35898 32000 35900
rect 31966 35866 32000 35898
rect 31966 35796 32000 35828
rect 31966 35794 32000 35796
rect 31966 35728 32000 35756
rect 31966 35722 32000 35728
rect 32077 35966 32111 35972
rect 32077 35938 32111 35966
rect 32077 35898 32111 35900
rect 32077 35866 32111 35898
rect 32077 35796 32111 35828
rect 32077 35794 32111 35796
rect 32077 35728 32111 35756
rect 32077 35722 32111 35728
rect 32163 35966 32197 35972
rect 32163 35938 32197 35966
rect 32163 35898 32197 35900
rect 32163 35866 32197 35898
rect 32163 35796 32197 35828
rect 32163 35794 32197 35796
rect 32163 35728 32197 35756
rect 32163 35722 32197 35728
rect 32249 35966 32283 35972
rect 32249 35938 32283 35966
rect 32249 35898 32283 35900
rect 32249 35866 32283 35898
rect 32249 35796 32283 35828
rect 32249 35794 32283 35796
rect 32249 35728 32283 35756
rect 32249 35722 32283 35728
rect 32360 35966 32394 35972
rect 32360 35938 32394 35966
rect 32360 35898 32394 35900
rect 32360 35866 32394 35898
rect 32360 35796 32394 35828
rect 32360 35794 32394 35796
rect 32360 35728 32394 35756
rect 32360 35722 32394 35728
rect 32091 35610 32095 35644
rect 32095 35610 32125 35644
rect 32163 35610 32197 35644
rect 32235 35610 32265 35644
rect 32265 35610 32269 35644
rect 32530 35624 32568 36021
rect 40992 35624 41030 36021
rect 41166 35966 41200 35972
rect 41166 35938 41200 35966
rect 41166 35898 41200 35900
rect 41166 35866 41200 35898
rect 41166 35796 41200 35828
rect 41166 35794 41200 35796
rect 41166 35728 41200 35756
rect 41166 35722 41200 35728
rect 41277 35966 41311 35972
rect 41277 35938 41311 35966
rect 41277 35898 41311 35900
rect 41277 35866 41311 35898
rect 41277 35796 41311 35828
rect 41277 35794 41311 35796
rect 41277 35728 41311 35756
rect 41277 35722 41311 35728
rect 41363 35966 41397 35972
rect 41363 35938 41397 35966
rect 41363 35898 41397 35900
rect 41363 35866 41397 35898
rect 41363 35796 41397 35828
rect 41363 35794 41397 35796
rect 41363 35728 41397 35756
rect 41363 35722 41397 35728
rect 41449 35966 41483 35972
rect 41449 35938 41483 35966
rect 41449 35898 41483 35900
rect 41449 35866 41483 35898
rect 41449 35796 41483 35828
rect 41449 35794 41483 35796
rect 41449 35728 41483 35756
rect 41449 35722 41483 35728
rect 41560 35966 41594 35972
rect 41560 35938 41594 35966
rect 41560 35898 41594 35900
rect 41560 35866 41594 35898
rect 41560 35796 41594 35828
rect 41560 35794 41594 35796
rect 41560 35728 41594 35756
rect 41560 35722 41594 35728
rect 41291 35610 41295 35644
rect 41295 35610 41325 35644
rect 41363 35610 41397 35644
rect 41435 35610 41465 35644
rect 41465 35610 41469 35644
rect 41730 35624 41768 36021
rect 50192 35624 50230 36021
rect 50366 35966 50400 35972
rect 50366 35938 50400 35966
rect 50366 35898 50400 35900
rect 50366 35866 50400 35898
rect 50366 35796 50400 35828
rect 50366 35794 50400 35796
rect 50366 35728 50400 35756
rect 50366 35722 50400 35728
rect 50477 35966 50511 35972
rect 50477 35938 50511 35966
rect 50477 35898 50511 35900
rect 50477 35866 50511 35898
rect 50477 35796 50511 35828
rect 50477 35794 50511 35796
rect 50477 35728 50511 35756
rect 50477 35722 50511 35728
rect 50563 35966 50597 35972
rect 50563 35938 50597 35966
rect 50563 35898 50597 35900
rect 50563 35866 50597 35898
rect 50563 35796 50597 35828
rect 50563 35794 50597 35796
rect 50563 35728 50597 35756
rect 50563 35722 50597 35728
rect 50649 35966 50683 35972
rect 50649 35938 50683 35966
rect 50649 35898 50683 35900
rect 50649 35866 50683 35898
rect 50649 35796 50683 35828
rect 50649 35794 50683 35796
rect 50649 35728 50683 35756
rect 50649 35722 50683 35728
rect 50760 35966 50794 35972
rect 50760 35938 50794 35966
rect 50760 35898 50794 35900
rect 50760 35866 50794 35898
rect 50760 35796 50794 35828
rect 50760 35794 50794 35796
rect 50760 35728 50794 35756
rect 50760 35722 50794 35728
rect 50491 35610 50495 35644
rect 50495 35610 50525 35644
rect 50563 35610 50597 35644
rect 50635 35610 50665 35644
rect 50665 35610 50669 35644
rect 50930 35624 50968 36021
rect 59392 35624 59430 36021
rect 59566 35966 59600 35972
rect 59566 35938 59600 35966
rect 59566 35898 59600 35900
rect 59566 35866 59600 35898
rect 59566 35796 59600 35828
rect 59566 35794 59600 35796
rect 59566 35728 59600 35756
rect 59566 35722 59600 35728
rect 59677 35966 59711 35972
rect 59677 35938 59711 35966
rect 59677 35898 59711 35900
rect 59677 35866 59711 35898
rect 59677 35796 59711 35828
rect 59677 35794 59711 35796
rect 59677 35728 59711 35756
rect 59677 35722 59711 35728
rect 59763 35966 59797 35972
rect 59763 35938 59797 35966
rect 59763 35898 59797 35900
rect 59763 35866 59797 35898
rect 59763 35796 59797 35828
rect 59763 35794 59797 35796
rect 59763 35728 59797 35756
rect 59763 35722 59797 35728
rect 59849 35966 59883 35972
rect 59849 35938 59883 35966
rect 59849 35898 59883 35900
rect 59849 35866 59883 35898
rect 59849 35796 59883 35828
rect 59849 35794 59883 35796
rect 59849 35728 59883 35756
rect 59849 35722 59883 35728
rect 59960 35966 59994 35972
rect 59960 35938 59994 35966
rect 59960 35898 59994 35900
rect 59960 35866 59994 35898
rect 59960 35796 59994 35828
rect 59960 35794 59994 35796
rect 59960 35728 59994 35756
rect 59960 35722 59994 35728
rect 59691 35610 59695 35644
rect 59695 35610 59725 35644
rect 59763 35610 59797 35644
rect 59835 35610 59865 35644
rect 59865 35610 59869 35644
rect 60130 35624 60168 36021
rect 68592 35624 68630 36021
rect 68766 35966 68800 35972
rect 68766 35938 68800 35966
rect 68766 35898 68800 35900
rect 68766 35866 68800 35898
rect 68766 35796 68800 35828
rect 68766 35794 68800 35796
rect 68766 35728 68800 35756
rect 68766 35722 68800 35728
rect 68877 35966 68911 35972
rect 68877 35938 68911 35966
rect 68877 35898 68911 35900
rect 68877 35866 68911 35898
rect 68877 35796 68911 35828
rect 68877 35794 68911 35796
rect 68877 35728 68911 35756
rect 68877 35722 68911 35728
rect 68963 35966 68997 35972
rect 68963 35938 68997 35966
rect 68963 35898 68997 35900
rect 68963 35866 68997 35898
rect 68963 35796 68997 35828
rect 68963 35794 68997 35796
rect 68963 35728 68997 35756
rect 68963 35722 68997 35728
rect 69049 35966 69083 35972
rect 69049 35938 69083 35966
rect 69049 35898 69083 35900
rect 69049 35866 69083 35898
rect 69049 35796 69083 35828
rect 69049 35794 69083 35796
rect 69049 35728 69083 35756
rect 69049 35722 69083 35728
rect 69160 35966 69194 35972
rect 69160 35938 69194 35966
rect 69160 35898 69194 35900
rect 69160 35866 69194 35898
rect 69160 35796 69194 35828
rect 69160 35794 69194 35796
rect 69160 35728 69194 35756
rect 69160 35722 69194 35728
rect 68891 35610 68895 35644
rect 68895 35610 68925 35644
rect 68963 35610 68997 35644
rect 69035 35610 69065 35644
rect 69065 35610 69069 35644
rect 69330 35624 69368 36021
rect 4192 26375 4230 26772
rect 4930 26375 4968 26772
rect 13392 26375 13430 26772
rect 14130 26375 14168 26772
rect 22592 26375 22630 26772
rect 23330 26375 23368 26772
rect 31792 26375 31830 26772
rect 32530 26375 32568 26772
rect 40992 26375 41030 26772
rect 41730 26375 41768 26772
rect 50192 26375 50230 26772
rect 50930 26375 50968 26772
rect 59392 26375 59430 26772
rect 60130 26375 60168 26772
rect 68592 26375 68630 26772
rect 69330 26375 69368 26772
rect 4491 26170 4495 26204
rect 4495 26170 4525 26204
rect 4563 26170 4597 26204
rect 4635 26170 4665 26204
rect 4665 26170 4669 26204
rect 13691 26170 13695 26204
rect 13695 26170 13725 26204
rect 13763 26170 13797 26204
rect 13835 26170 13865 26204
rect 13865 26170 13869 26204
rect 22891 26170 22895 26204
rect 22895 26170 22925 26204
rect 22963 26170 22997 26204
rect 23035 26170 23065 26204
rect 23065 26170 23069 26204
rect 32091 26170 32095 26204
rect 32095 26170 32125 26204
rect 32163 26170 32197 26204
rect 32235 26170 32265 26204
rect 32265 26170 32269 26204
rect 41291 26170 41295 26204
rect 41295 26170 41325 26204
rect 41363 26170 41397 26204
rect 41435 26170 41465 26204
rect 41465 26170 41469 26204
rect 50491 26170 50495 26204
rect 50495 26170 50525 26204
rect 50563 26170 50597 26204
rect 50635 26170 50665 26204
rect 50665 26170 50669 26204
rect 59691 26170 59695 26204
rect 59695 26170 59725 26204
rect 59763 26170 59797 26204
rect 59835 26170 59865 26204
rect 59865 26170 59869 26204
rect 68891 26170 68895 26204
rect 68895 26170 68925 26204
rect 68963 26170 68997 26204
rect 69035 26170 69065 26204
rect 69065 26170 69069 26204
rect 4192 25744 4230 26141
rect 4366 26086 4400 26092
rect 4366 26058 4400 26086
rect 4366 26018 4400 26020
rect 4366 25986 4400 26018
rect 4366 25916 4400 25948
rect 4366 25914 4400 25916
rect 4366 25848 4400 25876
rect 4366 25842 4400 25848
rect 4477 26086 4511 26092
rect 4477 26058 4511 26086
rect 4477 26018 4511 26020
rect 4477 25986 4511 26018
rect 4477 25916 4511 25948
rect 4477 25914 4511 25916
rect 4477 25848 4511 25876
rect 4477 25842 4511 25848
rect 4563 26086 4597 26092
rect 4563 26058 4597 26086
rect 4563 26018 4597 26020
rect 4563 25986 4597 26018
rect 4563 25916 4597 25948
rect 4563 25914 4597 25916
rect 4563 25848 4597 25876
rect 4563 25842 4597 25848
rect 4649 26086 4683 26092
rect 4649 26058 4683 26086
rect 4649 26018 4683 26020
rect 4649 25986 4683 26018
rect 4649 25916 4683 25948
rect 4649 25914 4683 25916
rect 4649 25848 4683 25876
rect 4649 25842 4683 25848
rect 4760 26086 4794 26092
rect 4760 26058 4794 26086
rect 4760 26018 4794 26020
rect 4760 25986 4794 26018
rect 4760 25916 4794 25948
rect 4760 25914 4794 25916
rect 4760 25848 4794 25876
rect 4760 25842 4794 25848
rect 4491 25730 4495 25764
rect 4495 25730 4525 25764
rect 4563 25730 4597 25764
rect 4635 25730 4665 25764
rect 4665 25730 4669 25764
rect 4930 25744 4968 26141
rect 13392 25744 13430 26141
rect 13566 26086 13600 26092
rect 13566 26058 13600 26086
rect 13566 26018 13600 26020
rect 13566 25986 13600 26018
rect 13566 25916 13600 25948
rect 13566 25914 13600 25916
rect 13566 25848 13600 25876
rect 13566 25842 13600 25848
rect 13677 26086 13711 26092
rect 13677 26058 13711 26086
rect 13677 26018 13711 26020
rect 13677 25986 13711 26018
rect 13677 25916 13711 25948
rect 13677 25914 13711 25916
rect 13677 25848 13711 25876
rect 13677 25842 13711 25848
rect 13763 26086 13797 26092
rect 13763 26058 13797 26086
rect 13763 26018 13797 26020
rect 13763 25986 13797 26018
rect 13763 25916 13797 25948
rect 13763 25914 13797 25916
rect 13763 25848 13797 25876
rect 13763 25842 13797 25848
rect 13849 26086 13883 26092
rect 13849 26058 13883 26086
rect 13849 26018 13883 26020
rect 13849 25986 13883 26018
rect 13849 25916 13883 25948
rect 13849 25914 13883 25916
rect 13849 25848 13883 25876
rect 13849 25842 13883 25848
rect 13960 26086 13994 26092
rect 13960 26058 13994 26086
rect 13960 26018 13994 26020
rect 13960 25986 13994 26018
rect 13960 25916 13994 25948
rect 13960 25914 13994 25916
rect 13960 25848 13994 25876
rect 13960 25842 13994 25848
rect 13691 25730 13695 25764
rect 13695 25730 13725 25764
rect 13763 25730 13797 25764
rect 13835 25730 13865 25764
rect 13865 25730 13869 25764
rect 14130 25744 14168 26141
rect 22592 25744 22630 26141
rect 22766 26086 22800 26092
rect 22766 26058 22800 26086
rect 22766 26018 22800 26020
rect 22766 25986 22800 26018
rect 22766 25916 22800 25948
rect 22766 25914 22800 25916
rect 22766 25848 22800 25876
rect 22766 25842 22800 25848
rect 22877 26086 22911 26092
rect 22877 26058 22911 26086
rect 22877 26018 22911 26020
rect 22877 25986 22911 26018
rect 22877 25916 22911 25948
rect 22877 25914 22911 25916
rect 22877 25848 22911 25876
rect 22877 25842 22911 25848
rect 22963 26086 22997 26092
rect 22963 26058 22997 26086
rect 22963 26018 22997 26020
rect 22963 25986 22997 26018
rect 22963 25916 22997 25948
rect 22963 25914 22997 25916
rect 22963 25848 22997 25876
rect 22963 25842 22997 25848
rect 23049 26086 23083 26092
rect 23049 26058 23083 26086
rect 23049 26018 23083 26020
rect 23049 25986 23083 26018
rect 23049 25916 23083 25948
rect 23049 25914 23083 25916
rect 23049 25848 23083 25876
rect 23049 25842 23083 25848
rect 23160 26086 23194 26092
rect 23160 26058 23194 26086
rect 23160 26018 23194 26020
rect 23160 25986 23194 26018
rect 23160 25916 23194 25948
rect 23160 25914 23194 25916
rect 23160 25848 23194 25876
rect 23160 25842 23194 25848
rect 22891 25730 22895 25764
rect 22895 25730 22925 25764
rect 22963 25730 22997 25764
rect 23035 25730 23065 25764
rect 23065 25730 23069 25764
rect 23330 25744 23368 26141
rect 31792 25744 31830 26141
rect 31966 26086 32000 26092
rect 31966 26058 32000 26086
rect 31966 26018 32000 26020
rect 31966 25986 32000 26018
rect 31966 25916 32000 25948
rect 31966 25914 32000 25916
rect 31966 25848 32000 25876
rect 31966 25842 32000 25848
rect 32077 26086 32111 26092
rect 32077 26058 32111 26086
rect 32077 26018 32111 26020
rect 32077 25986 32111 26018
rect 32077 25916 32111 25948
rect 32077 25914 32111 25916
rect 32077 25848 32111 25876
rect 32077 25842 32111 25848
rect 32163 26086 32197 26092
rect 32163 26058 32197 26086
rect 32163 26018 32197 26020
rect 32163 25986 32197 26018
rect 32163 25916 32197 25948
rect 32163 25914 32197 25916
rect 32163 25848 32197 25876
rect 32163 25842 32197 25848
rect 32249 26086 32283 26092
rect 32249 26058 32283 26086
rect 32249 26018 32283 26020
rect 32249 25986 32283 26018
rect 32249 25916 32283 25948
rect 32249 25914 32283 25916
rect 32249 25848 32283 25876
rect 32249 25842 32283 25848
rect 32360 26086 32394 26092
rect 32360 26058 32394 26086
rect 32360 26018 32394 26020
rect 32360 25986 32394 26018
rect 32360 25916 32394 25948
rect 32360 25914 32394 25916
rect 32360 25848 32394 25876
rect 32360 25842 32394 25848
rect 32091 25730 32095 25764
rect 32095 25730 32125 25764
rect 32163 25730 32197 25764
rect 32235 25730 32265 25764
rect 32265 25730 32269 25764
rect 32530 25744 32568 26141
rect 40992 25744 41030 26141
rect 41166 26086 41200 26092
rect 41166 26058 41200 26086
rect 41166 26018 41200 26020
rect 41166 25986 41200 26018
rect 41166 25916 41200 25948
rect 41166 25914 41200 25916
rect 41166 25848 41200 25876
rect 41166 25842 41200 25848
rect 41277 26086 41311 26092
rect 41277 26058 41311 26086
rect 41277 26018 41311 26020
rect 41277 25986 41311 26018
rect 41277 25916 41311 25948
rect 41277 25914 41311 25916
rect 41277 25848 41311 25876
rect 41277 25842 41311 25848
rect 41363 26086 41397 26092
rect 41363 26058 41397 26086
rect 41363 26018 41397 26020
rect 41363 25986 41397 26018
rect 41363 25916 41397 25948
rect 41363 25914 41397 25916
rect 41363 25848 41397 25876
rect 41363 25842 41397 25848
rect 41449 26086 41483 26092
rect 41449 26058 41483 26086
rect 41449 26018 41483 26020
rect 41449 25986 41483 26018
rect 41449 25916 41483 25948
rect 41449 25914 41483 25916
rect 41449 25848 41483 25876
rect 41449 25842 41483 25848
rect 41560 26086 41594 26092
rect 41560 26058 41594 26086
rect 41560 26018 41594 26020
rect 41560 25986 41594 26018
rect 41560 25916 41594 25948
rect 41560 25914 41594 25916
rect 41560 25848 41594 25876
rect 41560 25842 41594 25848
rect 41291 25730 41295 25764
rect 41295 25730 41325 25764
rect 41363 25730 41397 25764
rect 41435 25730 41465 25764
rect 41465 25730 41469 25764
rect 41730 25744 41768 26141
rect 50192 25744 50230 26141
rect 50366 26086 50400 26092
rect 50366 26058 50400 26086
rect 50366 26018 50400 26020
rect 50366 25986 50400 26018
rect 50366 25916 50400 25948
rect 50366 25914 50400 25916
rect 50366 25848 50400 25876
rect 50366 25842 50400 25848
rect 50477 26086 50511 26092
rect 50477 26058 50511 26086
rect 50477 26018 50511 26020
rect 50477 25986 50511 26018
rect 50477 25916 50511 25948
rect 50477 25914 50511 25916
rect 50477 25848 50511 25876
rect 50477 25842 50511 25848
rect 50563 26086 50597 26092
rect 50563 26058 50597 26086
rect 50563 26018 50597 26020
rect 50563 25986 50597 26018
rect 50563 25916 50597 25948
rect 50563 25914 50597 25916
rect 50563 25848 50597 25876
rect 50563 25842 50597 25848
rect 50649 26086 50683 26092
rect 50649 26058 50683 26086
rect 50649 26018 50683 26020
rect 50649 25986 50683 26018
rect 50649 25916 50683 25948
rect 50649 25914 50683 25916
rect 50649 25848 50683 25876
rect 50649 25842 50683 25848
rect 50760 26086 50794 26092
rect 50760 26058 50794 26086
rect 50760 26018 50794 26020
rect 50760 25986 50794 26018
rect 50760 25916 50794 25948
rect 50760 25914 50794 25916
rect 50760 25848 50794 25876
rect 50760 25842 50794 25848
rect 50491 25730 50495 25764
rect 50495 25730 50525 25764
rect 50563 25730 50597 25764
rect 50635 25730 50665 25764
rect 50665 25730 50669 25764
rect 50930 25744 50968 26141
rect 59392 25744 59430 26141
rect 59566 26086 59600 26092
rect 59566 26058 59600 26086
rect 59566 26018 59600 26020
rect 59566 25986 59600 26018
rect 59566 25916 59600 25948
rect 59566 25914 59600 25916
rect 59566 25848 59600 25876
rect 59566 25842 59600 25848
rect 59677 26086 59711 26092
rect 59677 26058 59711 26086
rect 59677 26018 59711 26020
rect 59677 25986 59711 26018
rect 59677 25916 59711 25948
rect 59677 25914 59711 25916
rect 59677 25848 59711 25876
rect 59677 25842 59711 25848
rect 59763 26086 59797 26092
rect 59763 26058 59797 26086
rect 59763 26018 59797 26020
rect 59763 25986 59797 26018
rect 59763 25916 59797 25948
rect 59763 25914 59797 25916
rect 59763 25848 59797 25876
rect 59763 25842 59797 25848
rect 59849 26086 59883 26092
rect 59849 26058 59883 26086
rect 59849 26018 59883 26020
rect 59849 25986 59883 26018
rect 59849 25916 59883 25948
rect 59849 25914 59883 25916
rect 59849 25848 59883 25876
rect 59849 25842 59883 25848
rect 59960 26086 59994 26092
rect 59960 26058 59994 26086
rect 59960 26018 59994 26020
rect 59960 25986 59994 26018
rect 59960 25916 59994 25948
rect 59960 25914 59994 25916
rect 59960 25848 59994 25876
rect 59960 25842 59994 25848
rect 59691 25730 59695 25764
rect 59695 25730 59725 25764
rect 59763 25730 59797 25764
rect 59835 25730 59865 25764
rect 59865 25730 59869 25764
rect 60130 25744 60168 26141
rect 68592 25744 68630 26141
rect 68766 26086 68800 26092
rect 68766 26058 68800 26086
rect 68766 26018 68800 26020
rect 68766 25986 68800 26018
rect 68766 25916 68800 25948
rect 68766 25914 68800 25916
rect 68766 25848 68800 25876
rect 68766 25842 68800 25848
rect 68877 26086 68911 26092
rect 68877 26058 68911 26086
rect 68877 26018 68911 26020
rect 68877 25986 68911 26018
rect 68877 25916 68911 25948
rect 68877 25914 68911 25916
rect 68877 25848 68911 25876
rect 68877 25842 68911 25848
rect 68963 26086 68997 26092
rect 68963 26058 68997 26086
rect 68963 26018 68997 26020
rect 68963 25986 68997 26018
rect 68963 25916 68997 25948
rect 68963 25914 68997 25916
rect 68963 25848 68997 25876
rect 68963 25842 68997 25848
rect 69049 26086 69083 26092
rect 69049 26058 69083 26086
rect 69049 26018 69083 26020
rect 69049 25986 69083 26018
rect 69049 25916 69083 25948
rect 69049 25914 69083 25916
rect 69049 25848 69083 25876
rect 69049 25842 69083 25848
rect 69160 26086 69194 26092
rect 69160 26058 69194 26086
rect 69160 26018 69194 26020
rect 69160 25986 69194 26018
rect 69160 25916 69194 25948
rect 69160 25914 69194 25916
rect 69160 25848 69194 25876
rect 69160 25842 69194 25848
rect 68891 25730 68895 25764
rect 68895 25730 68925 25764
rect 68963 25730 68997 25764
rect 69035 25730 69065 25764
rect 69065 25730 69069 25764
rect 69330 25744 69368 26141
rect 4192 16495 4230 16892
rect 4930 16495 4968 16892
rect 13392 16495 13430 16892
rect 14130 16495 14168 16892
rect 22592 16495 22630 16892
rect 23330 16495 23368 16892
rect 31792 16495 31830 16892
rect 32530 16495 32568 16892
rect 40992 16495 41030 16892
rect 41730 16495 41768 16892
rect 50192 16495 50230 16892
rect 50930 16495 50968 16892
rect 59392 16495 59430 16892
rect 60130 16495 60168 16892
rect 68592 16495 68630 16892
rect 69330 16495 69368 16892
rect 4491 16290 4495 16324
rect 4495 16290 4525 16324
rect 4563 16290 4597 16324
rect 4635 16290 4665 16324
rect 4665 16290 4669 16324
rect 13691 16290 13695 16324
rect 13695 16290 13725 16324
rect 13763 16290 13797 16324
rect 13835 16290 13865 16324
rect 13865 16290 13869 16324
rect 22891 16290 22895 16324
rect 22895 16290 22925 16324
rect 22963 16290 22997 16324
rect 23035 16290 23065 16324
rect 23065 16290 23069 16324
rect 32091 16290 32095 16324
rect 32095 16290 32125 16324
rect 32163 16290 32197 16324
rect 32235 16290 32265 16324
rect 32265 16290 32269 16324
rect 41291 16290 41295 16324
rect 41295 16290 41325 16324
rect 41363 16290 41397 16324
rect 41435 16290 41465 16324
rect 41465 16290 41469 16324
rect 50491 16290 50495 16324
rect 50495 16290 50525 16324
rect 50563 16290 50597 16324
rect 50635 16290 50665 16324
rect 50665 16290 50669 16324
rect 59691 16290 59695 16324
rect 59695 16290 59725 16324
rect 59763 16290 59797 16324
rect 59835 16290 59865 16324
rect 59865 16290 59869 16324
rect 68891 16290 68895 16324
rect 68895 16290 68925 16324
rect 68963 16290 68997 16324
rect 69035 16290 69065 16324
rect 69065 16290 69069 16324
rect 4192 15864 4230 16261
rect 4366 16206 4400 16212
rect 4366 16178 4400 16206
rect 4366 16138 4400 16140
rect 4366 16106 4400 16138
rect 4366 16036 4400 16068
rect 4366 16034 4400 16036
rect 4366 15968 4400 15996
rect 4366 15962 4400 15968
rect 4477 16206 4511 16212
rect 4477 16178 4511 16206
rect 4477 16138 4511 16140
rect 4477 16106 4511 16138
rect 4477 16036 4511 16068
rect 4477 16034 4511 16036
rect 4477 15968 4511 15996
rect 4477 15962 4511 15968
rect 4563 16206 4597 16212
rect 4563 16178 4597 16206
rect 4563 16138 4597 16140
rect 4563 16106 4597 16138
rect 4563 16036 4597 16068
rect 4563 16034 4597 16036
rect 4563 15968 4597 15996
rect 4563 15962 4597 15968
rect 4649 16206 4683 16212
rect 4649 16178 4683 16206
rect 4649 16138 4683 16140
rect 4649 16106 4683 16138
rect 4649 16036 4683 16068
rect 4649 16034 4683 16036
rect 4649 15968 4683 15996
rect 4649 15962 4683 15968
rect 4760 16206 4794 16212
rect 4760 16178 4794 16206
rect 4760 16138 4794 16140
rect 4760 16106 4794 16138
rect 4760 16036 4794 16068
rect 4760 16034 4794 16036
rect 4760 15968 4794 15996
rect 4760 15962 4794 15968
rect 4491 15850 4495 15884
rect 4495 15850 4525 15884
rect 4563 15850 4597 15884
rect 4635 15850 4665 15884
rect 4665 15850 4669 15884
rect 4930 15864 4968 16261
rect 13392 15864 13430 16261
rect 13566 16206 13600 16212
rect 13566 16178 13600 16206
rect 13566 16138 13600 16140
rect 13566 16106 13600 16138
rect 13566 16036 13600 16068
rect 13566 16034 13600 16036
rect 13566 15968 13600 15996
rect 13566 15962 13600 15968
rect 13677 16206 13711 16212
rect 13677 16178 13711 16206
rect 13677 16138 13711 16140
rect 13677 16106 13711 16138
rect 13677 16036 13711 16068
rect 13677 16034 13711 16036
rect 13677 15968 13711 15996
rect 13677 15962 13711 15968
rect 13763 16206 13797 16212
rect 13763 16178 13797 16206
rect 13763 16138 13797 16140
rect 13763 16106 13797 16138
rect 13763 16036 13797 16068
rect 13763 16034 13797 16036
rect 13763 15968 13797 15996
rect 13763 15962 13797 15968
rect 13849 16206 13883 16212
rect 13849 16178 13883 16206
rect 13849 16138 13883 16140
rect 13849 16106 13883 16138
rect 13849 16036 13883 16068
rect 13849 16034 13883 16036
rect 13849 15968 13883 15996
rect 13849 15962 13883 15968
rect 13960 16206 13994 16212
rect 13960 16178 13994 16206
rect 13960 16138 13994 16140
rect 13960 16106 13994 16138
rect 13960 16036 13994 16068
rect 13960 16034 13994 16036
rect 13960 15968 13994 15996
rect 13960 15962 13994 15968
rect 13691 15850 13695 15884
rect 13695 15850 13725 15884
rect 13763 15850 13797 15884
rect 13835 15850 13865 15884
rect 13865 15850 13869 15884
rect 14130 15864 14168 16261
rect 22592 15864 22630 16261
rect 22766 16206 22800 16212
rect 22766 16178 22800 16206
rect 22766 16138 22800 16140
rect 22766 16106 22800 16138
rect 22766 16036 22800 16068
rect 22766 16034 22800 16036
rect 22766 15968 22800 15996
rect 22766 15962 22800 15968
rect 22877 16206 22911 16212
rect 22877 16178 22911 16206
rect 22877 16138 22911 16140
rect 22877 16106 22911 16138
rect 22877 16036 22911 16068
rect 22877 16034 22911 16036
rect 22877 15968 22911 15996
rect 22877 15962 22911 15968
rect 22963 16206 22997 16212
rect 22963 16178 22997 16206
rect 22963 16138 22997 16140
rect 22963 16106 22997 16138
rect 22963 16036 22997 16068
rect 22963 16034 22997 16036
rect 22963 15968 22997 15996
rect 22963 15962 22997 15968
rect 23049 16206 23083 16212
rect 23049 16178 23083 16206
rect 23049 16138 23083 16140
rect 23049 16106 23083 16138
rect 23049 16036 23083 16068
rect 23049 16034 23083 16036
rect 23049 15968 23083 15996
rect 23049 15962 23083 15968
rect 23160 16206 23194 16212
rect 23160 16178 23194 16206
rect 23160 16138 23194 16140
rect 23160 16106 23194 16138
rect 23160 16036 23194 16068
rect 23160 16034 23194 16036
rect 23160 15968 23194 15996
rect 23160 15962 23194 15968
rect 22891 15850 22895 15884
rect 22895 15850 22925 15884
rect 22963 15850 22997 15884
rect 23035 15850 23065 15884
rect 23065 15850 23069 15884
rect 23330 15864 23368 16261
rect 31792 15864 31830 16261
rect 31966 16206 32000 16212
rect 31966 16178 32000 16206
rect 31966 16138 32000 16140
rect 31966 16106 32000 16138
rect 31966 16036 32000 16068
rect 31966 16034 32000 16036
rect 31966 15968 32000 15996
rect 31966 15962 32000 15968
rect 32077 16206 32111 16212
rect 32077 16178 32111 16206
rect 32077 16138 32111 16140
rect 32077 16106 32111 16138
rect 32077 16036 32111 16068
rect 32077 16034 32111 16036
rect 32077 15968 32111 15996
rect 32077 15962 32111 15968
rect 32163 16206 32197 16212
rect 32163 16178 32197 16206
rect 32163 16138 32197 16140
rect 32163 16106 32197 16138
rect 32163 16036 32197 16068
rect 32163 16034 32197 16036
rect 32163 15968 32197 15996
rect 32163 15962 32197 15968
rect 32249 16206 32283 16212
rect 32249 16178 32283 16206
rect 32249 16138 32283 16140
rect 32249 16106 32283 16138
rect 32249 16036 32283 16068
rect 32249 16034 32283 16036
rect 32249 15968 32283 15996
rect 32249 15962 32283 15968
rect 32360 16206 32394 16212
rect 32360 16178 32394 16206
rect 32360 16138 32394 16140
rect 32360 16106 32394 16138
rect 32360 16036 32394 16068
rect 32360 16034 32394 16036
rect 32360 15968 32394 15996
rect 32360 15962 32394 15968
rect 32091 15850 32095 15884
rect 32095 15850 32125 15884
rect 32163 15850 32197 15884
rect 32235 15850 32265 15884
rect 32265 15850 32269 15884
rect 32530 15864 32568 16261
rect 40992 15864 41030 16261
rect 41166 16206 41200 16212
rect 41166 16178 41200 16206
rect 41166 16138 41200 16140
rect 41166 16106 41200 16138
rect 41166 16036 41200 16068
rect 41166 16034 41200 16036
rect 41166 15968 41200 15996
rect 41166 15962 41200 15968
rect 41277 16206 41311 16212
rect 41277 16178 41311 16206
rect 41277 16138 41311 16140
rect 41277 16106 41311 16138
rect 41277 16036 41311 16068
rect 41277 16034 41311 16036
rect 41277 15968 41311 15996
rect 41277 15962 41311 15968
rect 41363 16206 41397 16212
rect 41363 16178 41397 16206
rect 41363 16138 41397 16140
rect 41363 16106 41397 16138
rect 41363 16036 41397 16068
rect 41363 16034 41397 16036
rect 41363 15968 41397 15996
rect 41363 15962 41397 15968
rect 41449 16206 41483 16212
rect 41449 16178 41483 16206
rect 41449 16138 41483 16140
rect 41449 16106 41483 16138
rect 41449 16036 41483 16068
rect 41449 16034 41483 16036
rect 41449 15968 41483 15996
rect 41449 15962 41483 15968
rect 41560 16206 41594 16212
rect 41560 16178 41594 16206
rect 41560 16138 41594 16140
rect 41560 16106 41594 16138
rect 41560 16036 41594 16068
rect 41560 16034 41594 16036
rect 41560 15968 41594 15996
rect 41560 15962 41594 15968
rect 41291 15850 41295 15884
rect 41295 15850 41325 15884
rect 41363 15850 41397 15884
rect 41435 15850 41465 15884
rect 41465 15850 41469 15884
rect 41730 15864 41768 16261
rect 50192 15864 50230 16261
rect 50366 16206 50400 16212
rect 50366 16178 50400 16206
rect 50366 16138 50400 16140
rect 50366 16106 50400 16138
rect 50366 16036 50400 16068
rect 50366 16034 50400 16036
rect 50366 15968 50400 15996
rect 50366 15962 50400 15968
rect 50477 16206 50511 16212
rect 50477 16178 50511 16206
rect 50477 16138 50511 16140
rect 50477 16106 50511 16138
rect 50477 16036 50511 16068
rect 50477 16034 50511 16036
rect 50477 15968 50511 15996
rect 50477 15962 50511 15968
rect 50563 16206 50597 16212
rect 50563 16178 50597 16206
rect 50563 16138 50597 16140
rect 50563 16106 50597 16138
rect 50563 16036 50597 16068
rect 50563 16034 50597 16036
rect 50563 15968 50597 15996
rect 50563 15962 50597 15968
rect 50649 16206 50683 16212
rect 50649 16178 50683 16206
rect 50649 16138 50683 16140
rect 50649 16106 50683 16138
rect 50649 16036 50683 16068
rect 50649 16034 50683 16036
rect 50649 15968 50683 15996
rect 50649 15962 50683 15968
rect 50760 16206 50794 16212
rect 50760 16178 50794 16206
rect 50760 16138 50794 16140
rect 50760 16106 50794 16138
rect 50760 16036 50794 16068
rect 50760 16034 50794 16036
rect 50760 15968 50794 15996
rect 50760 15962 50794 15968
rect 50491 15850 50495 15884
rect 50495 15850 50525 15884
rect 50563 15850 50597 15884
rect 50635 15850 50665 15884
rect 50665 15850 50669 15884
rect 50930 15864 50968 16261
rect 59392 15864 59430 16261
rect 59566 16206 59600 16212
rect 59566 16178 59600 16206
rect 59566 16138 59600 16140
rect 59566 16106 59600 16138
rect 59566 16036 59600 16068
rect 59566 16034 59600 16036
rect 59566 15968 59600 15996
rect 59566 15962 59600 15968
rect 59677 16206 59711 16212
rect 59677 16178 59711 16206
rect 59677 16138 59711 16140
rect 59677 16106 59711 16138
rect 59677 16036 59711 16068
rect 59677 16034 59711 16036
rect 59677 15968 59711 15996
rect 59677 15962 59711 15968
rect 59763 16206 59797 16212
rect 59763 16178 59797 16206
rect 59763 16138 59797 16140
rect 59763 16106 59797 16138
rect 59763 16036 59797 16068
rect 59763 16034 59797 16036
rect 59763 15968 59797 15996
rect 59763 15962 59797 15968
rect 59849 16206 59883 16212
rect 59849 16178 59883 16206
rect 59849 16138 59883 16140
rect 59849 16106 59883 16138
rect 59849 16036 59883 16068
rect 59849 16034 59883 16036
rect 59849 15968 59883 15996
rect 59849 15962 59883 15968
rect 59960 16206 59994 16212
rect 59960 16178 59994 16206
rect 59960 16138 59994 16140
rect 59960 16106 59994 16138
rect 59960 16036 59994 16068
rect 59960 16034 59994 16036
rect 59960 15968 59994 15996
rect 59960 15962 59994 15968
rect 59691 15850 59695 15884
rect 59695 15850 59725 15884
rect 59763 15850 59797 15884
rect 59835 15850 59865 15884
rect 59865 15850 59869 15884
rect 60130 15864 60168 16261
rect 68592 15864 68630 16261
rect 68766 16206 68800 16212
rect 68766 16178 68800 16206
rect 68766 16138 68800 16140
rect 68766 16106 68800 16138
rect 68766 16036 68800 16068
rect 68766 16034 68800 16036
rect 68766 15968 68800 15996
rect 68766 15962 68800 15968
rect 68877 16206 68911 16212
rect 68877 16178 68911 16206
rect 68877 16138 68911 16140
rect 68877 16106 68911 16138
rect 68877 16036 68911 16068
rect 68877 16034 68911 16036
rect 68877 15968 68911 15996
rect 68877 15962 68911 15968
rect 68963 16206 68997 16212
rect 68963 16178 68997 16206
rect 68963 16138 68997 16140
rect 68963 16106 68997 16138
rect 68963 16036 68997 16068
rect 68963 16034 68997 16036
rect 68963 15968 68997 15996
rect 68963 15962 68997 15968
rect 69049 16206 69083 16212
rect 69049 16178 69083 16206
rect 69049 16138 69083 16140
rect 69049 16106 69083 16138
rect 69049 16036 69083 16068
rect 69049 16034 69083 16036
rect 69049 15968 69083 15996
rect 69049 15962 69083 15968
rect 69160 16206 69194 16212
rect 69160 16178 69194 16206
rect 69160 16138 69194 16140
rect 69160 16106 69194 16138
rect 69160 16036 69194 16068
rect 69160 16034 69194 16036
rect 69160 15968 69194 15996
rect 69160 15962 69194 15968
rect 68891 15850 68895 15884
rect 68895 15850 68925 15884
rect 68963 15850 68997 15884
rect 69035 15850 69065 15884
rect 69065 15850 69069 15884
rect 69330 15864 69368 16261
rect -480 6570 -440 6610
rect -400 6574 -392 6610
rect -392 6574 -360 6610
rect -310 6574 -278 6610
rect -278 6574 -270 6610
rect -400 6570 -360 6574
rect -310 6570 -270 6574
rect 4192 6615 4230 7012
rect 4930 6615 4968 7012
rect 13392 6615 13430 7012
rect 14130 6615 14168 7012
rect 22592 6615 22630 7012
rect 23330 6615 23368 7012
rect 31792 6615 31830 7012
rect 32530 6615 32568 7012
rect 40992 6615 41030 7012
rect 41730 6615 41768 7012
rect 50192 6615 50230 7012
rect 50930 6615 50968 7012
rect 59392 6615 59430 7012
rect 60130 6615 60168 7012
rect 68592 6615 68630 7012
rect 69330 6615 69368 7012
rect -424 5888 -390 6464
rect -600 5800 -560 5840
rect -336 5888 -302 6464
rect 4491 6410 4495 6444
rect 4495 6410 4525 6444
rect 4563 6410 4597 6444
rect 4635 6410 4665 6444
rect 4665 6410 4669 6444
rect 13691 6410 13695 6444
rect 13695 6410 13725 6444
rect 13763 6410 13797 6444
rect 13835 6410 13865 6444
rect 13865 6410 13869 6444
rect 22891 6410 22895 6444
rect 22895 6410 22925 6444
rect 22963 6410 22997 6444
rect 23035 6410 23065 6444
rect 23065 6410 23069 6444
rect 32091 6410 32095 6444
rect 32095 6410 32125 6444
rect 32163 6410 32197 6444
rect 32235 6410 32265 6444
rect 32265 6410 32269 6444
rect 41291 6410 41295 6444
rect 41295 6410 41325 6444
rect 41363 6410 41397 6444
rect 41435 6410 41465 6444
rect 41465 6410 41469 6444
rect 50491 6410 50495 6444
rect 50495 6410 50525 6444
rect 50563 6410 50597 6444
rect 50635 6410 50665 6444
rect 50665 6410 50669 6444
rect 59691 6410 59695 6444
rect 59695 6410 59725 6444
rect 59763 6410 59797 6444
rect 59835 6410 59865 6444
rect 59865 6410 59869 6444
rect 68891 6410 68895 6444
rect 68895 6410 68925 6444
rect 68963 6410 68997 6444
rect 69035 6410 69065 6444
rect 69065 6410 69069 6444
rect 4192 5984 4230 6381
rect 4366 6326 4400 6332
rect 4366 6298 4400 6326
rect 4366 6258 4400 6260
rect 4366 6226 4400 6258
rect 4366 6156 4400 6188
rect 4366 6154 4400 6156
rect 4366 6088 4400 6116
rect 4366 6082 4400 6088
rect 4477 6326 4511 6332
rect 4477 6298 4511 6326
rect 4477 6258 4511 6260
rect 4477 6226 4511 6258
rect 4477 6156 4511 6188
rect 4477 6154 4511 6156
rect 4477 6088 4511 6116
rect 4477 6082 4511 6088
rect 4563 6326 4597 6332
rect 4563 6298 4597 6326
rect 4563 6258 4597 6260
rect 4563 6226 4597 6258
rect 4563 6156 4597 6188
rect 4563 6154 4597 6156
rect 4563 6088 4597 6116
rect 4563 6082 4597 6088
rect 4649 6326 4683 6332
rect 4649 6298 4683 6326
rect 4649 6258 4683 6260
rect 4649 6226 4683 6258
rect 4649 6156 4683 6188
rect 4649 6154 4683 6156
rect 4649 6088 4683 6116
rect 4649 6082 4683 6088
rect 4760 6326 4794 6332
rect 4760 6298 4794 6326
rect 4760 6258 4794 6260
rect 4760 6226 4794 6258
rect 4760 6156 4794 6188
rect 4760 6154 4794 6156
rect 4760 6088 4794 6116
rect 4760 6082 4794 6088
rect 4491 5970 4495 6004
rect 4495 5970 4525 6004
rect 4563 5970 4597 6004
rect 4635 5970 4665 6004
rect 4665 5970 4669 6004
rect 4930 5984 4968 6381
rect 13392 5984 13430 6381
rect 13566 6326 13600 6332
rect 13566 6298 13600 6326
rect 13566 6258 13600 6260
rect 13566 6226 13600 6258
rect 13566 6156 13600 6188
rect 13566 6154 13600 6156
rect 13566 6088 13600 6116
rect 13566 6082 13600 6088
rect 13677 6326 13711 6332
rect 13677 6298 13711 6326
rect 13677 6258 13711 6260
rect 13677 6226 13711 6258
rect 13677 6156 13711 6188
rect 13677 6154 13711 6156
rect 13677 6088 13711 6116
rect 13677 6082 13711 6088
rect 13763 6326 13797 6332
rect 13763 6298 13797 6326
rect 13763 6258 13797 6260
rect 13763 6226 13797 6258
rect 13763 6156 13797 6188
rect 13763 6154 13797 6156
rect 13763 6088 13797 6116
rect 13763 6082 13797 6088
rect 13849 6326 13883 6332
rect 13849 6298 13883 6326
rect 13849 6258 13883 6260
rect 13849 6226 13883 6258
rect 13849 6156 13883 6188
rect 13849 6154 13883 6156
rect 13849 6088 13883 6116
rect 13849 6082 13883 6088
rect 13960 6326 13994 6332
rect 13960 6298 13994 6326
rect 13960 6258 13994 6260
rect 13960 6226 13994 6258
rect 13960 6156 13994 6188
rect 13960 6154 13994 6156
rect 13960 6088 13994 6116
rect 13960 6082 13994 6088
rect 13691 5970 13695 6004
rect 13695 5970 13725 6004
rect 13763 5970 13797 6004
rect 13835 5970 13865 6004
rect 13865 5970 13869 6004
rect 14130 5984 14168 6381
rect 22592 5984 22630 6381
rect 22766 6326 22800 6332
rect 22766 6298 22800 6326
rect 22766 6258 22800 6260
rect 22766 6226 22800 6258
rect 22766 6156 22800 6188
rect 22766 6154 22800 6156
rect 22766 6088 22800 6116
rect 22766 6082 22800 6088
rect 22877 6326 22911 6332
rect 22877 6298 22911 6326
rect 22877 6258 22911 6260
rect 22877 6226 22911 6258
rect 22877 6156 22911 6188
rect 22877 6154 22911 6156
rect 22877 6088 22911 6116
rect 22877 6082 22911 6088
rect 22963 6326 22997 6332
rect 22963 6298 22997 6326
rect 22963 6258 22997 6260
rect 22963 6226 22997 6258
rect 22963 6156 22997 6188
rect 22963 6154 22997 6156
rect 22963 6088 22997 6116
rect 22963 6082 22997 6088
rect 23049 6326 23083 6332
rect 23049 6298 23083 6326
rect 23049 6258 23083 6260
rect 23049 6226 23083 6258
rect 23049 6156 23083 6188
rect 23049 6154 23083 6156
rect 23049 6088 23083 6116
rect 23049 6082 23083 6088
rect 23160 6326 23194 6332
rect 23160 6298 23194 6326
rect 23160 6258 23194 6260
rect 23160 6226 23194 6258
rect 23160 6156 23194 6188
rect 23160 6154 23194 6156
rect 23160 6088 23194 6116
rect 23160 6082 23194 6088
rect 22891 5970 22895 6004
rect 22895 5970 22925 6004
rect 22963 5970 22997 6004
rect 23035 5970 23065 6004
rect 23065 5970 23069 6004
rect 23330 5984 23368 6381
rect 31792 5984 31830 6381
rect 31966 6326 32000 6332
rect 31966 6298 32000 6326
rect 31966 6258 32000 6260
rect 31966 6226 32000 6258
rect 31966 6156 32000 6188
rect 31966 6154 32000 6156
rect 31966 6088 32000 6116
rect 31966 6082 32000 6088
rect 32077 6326 32111 6332
rect 32077 6298 32111 6326
rect 32077 6258 32111 6260
rect 32077 6226 32111 6258
rect 32077 6156 32111 6188
rect 32077 6154 32111 6156
rect 32077 6088 32111 6116
rect 32077 6082 32111 6088
rect 32163 6326 32197 6332
rect 32163 6298 32197 6326
rect 32163 6258 32197 6260
rect 32163 6226 32197 6258
rect 32163 6156 32197 6188
rect 32163 6154 32197 6156
rect 32163 6088 32197 6116
rect 32163 6082 32197 6088
rect 32249 6326 32283 6332
rect 32249 6298 32283 6326
rect 32249 6258 32283 6260
rect 32249 6226 32283 6258
rect 32249 6156 32283 6188
rect 32249 6154 32283 6156
rect 32249 6088 32283 6116
rect 32249 6082 32283 6088
rect 32360 6326 32394 6332
rect 32360 6298 32394 6326
rect 32360 6258 32394 6260
rect 32360 6226 32394 6258
rect 32360 6156 32394 6188
rect 32360 6154 32394 6156
rect 32360 6088 32394 6116
rect 32360 6082 32394 6088
rect 32091 5970 32095 6004
rect 32095 5970 32125 6004
rect 32163 5970 32197 6004
rect 32235 5970 32265 6004
rect 32265 5970 32269 6004
rect 32530 5984 32568 6381
rect 40992 5984 41030 6381
rect 41166 6326 41200 6332
rect 41166 6298 41200 6326
rect 41166 6258 41200 6260
rect 41166 6226 41200 6258
rect 41166 6156 41200 6188
rect 41166 6154 41200 6156
rect 41166 6088 41200 6116
rect 41166 6082 41200 6088
rect 41277 6326 41311 6332
rect 41277 6298 41311 6326
rect 41277 6258 41311 6260
rect 41277 6226 41311 6258
rect 41277 6156 41311 6188
rect 41277 6154 41311 6156
rect 41277 6088 41311 6116
rect 41277 6082 41311 6088
rect 41363 6326 41397 6332
rect 41363 6298 41397 6326
rect 41363 6258 41397 6260
rect 41363 6226 41397 6258
rect 41363 6156 41397 6188
rect 41363 6154 41397 6156
rect 41363 6088 41397 6116
rect 41363 6082 41397 6088
rect 41449 6326 41483 6332
rect 41449 6298 41483 6326
rect 41449 6258 41483 6260
rect 41449 6226 41483 6258
rect 41449 6156 41483 6188
rect 41449 6154 41483 6156
rect 41449 6088 41483 6116
rect 41449 6082 41483 6088
rect 41560 6326 41594 6332
rect 41560 6298 41594 6326
rect 41560 6258 41594 6260
rect 41560 6226 41594 6258
rect 41560 6156 41594 6188
rect 41560 6154 41594 6156
rect 41560 6088 41594 6116
rect 41560 6082 41594 6088
rect 41291 5970 41295 6004
rect 41295 5970 41325 6004
rect 41363 5970 41397 6004
rect 41435 5970 41465 6004
rect 41465 5970 41469 6004
rect 41730 5984 41768 6381
rect 50192 5984 50230 6381
rect 50366 6326 50400 6332
rect 50366 6298 50400 6326
rect 50366 6258 50400 6260
rect 50366 6226 50400 6258
rect 50366 6156 50400 6188
rect 50366 6154 50400 6156
rect 50366 6088 50400 6116
rect 50366 6082 50400 6088
rect 50477 6326 50511 6332
rect 50477 6298 50511 6326
rect 50477 6258 50511 6260
rect 50477 6226 50511 6258
rect 50477 6156 50511 6188
rect 50477 6154 50511 6156
rect 50477 6088 50511 6116
rect 50477 6082 50511 6088
rect 50563 6326 50597 6332
rect 50563 6298 50597 6326
rect 50563 6258 50597 6260
rect 50563 6226 50597 6258
rect 50563 6156 50597 6188
rect 50563 6154 50597 6156
rect 50563 6088 50597 6116
rect 50563 6082 50597 6088
rect 50649 6326 50683 6332
rect 50649 6298 50683 6326
rect 50649 6258 50683 6260
rect 50649 6226 50683 6258
rect 50649 6156 50683 6188
rect 50649 6154 50683 6156
rect 50649 6088 50683 6116
rect 50649 6082 50683 6088
rect 50760 6326 50794 6332
rect 50760 6298 50794 6326
rect 50760 6258 50794 6260
rect 50760 6226 50794 6258
rect 50760 6156 50794 6188
rect 50760 6154 50794 6156
rect 50760 6088 50794 6116
rect 50760 6082 50794 6088
rect 50491 5970 50495 6004
rect 50495 5970 50525 6004
rect 50563 5970 50597 6004
rect 50635 5970 50665 6004
rect 50665 5970 50669 6004
rect 50930 5984 50968 6381
rect 59392 5984 59430 6381
rect 59566 6326 59600 6332
rect 59566 6298 59600 6326
rect 59566 6258 59600 6260
rect 59566 6226 59600 6258
rect 59566 6156 59600 6188
rect 59566 6154 59600 6156
rect 59566 6088 59600 6116
rect 59566 6082 59600 6088
rect 59677 6326 59711 6332
rect 59677 6298 59711 6326
rect 59677 6258 59711 6260
rect 59677 6226 59711 6258
rect 59677 6156 59711 6188
rect 59677 6154 59711 6156
rect 59677 6088 59711 6116
rect 59677 6082 59711 6088
rect 59763 6326 59797 6332
rect 59763 6298 59797 6326
rect 59763 6258 59797 6260
rect 59763 6226 59797 6258
rect 59763 6156 59797 6188
rect 59763 6154 59797 6156
rect 59763 6088 59797 6116
rect 59763 6082 59797 6088
rect 59849 6326 59883 6332
rect 59849 6298 59883 6326
rect 59849 6258 59883 6260
rect 59849 6226 59883 6258
rect 59849 6156 59883 6188
rect 59849 6154 59883 6156
rect 59849 6088 59883 6116
rect 59849 6082 59883 6088
rect 59960 6326 59994 6332
rect 59960 6298 59994 6326
rect 59960 6258 59994 6260
rect 59960 6226 59994 6258
rect 59960 6156 59994 6188
rect 59960 6154 59994 6156
rect 59960 6088 59994 6116
rect 59960 6082 59994 6088
rect 59691 5970 59695 6004
rect 59695 5970 59725 6004
rect 59763 5970 59797 6004
rect 59835 5970 59865 6004
rect 59865 5970 59869 6004
rect 60130 5984 60168 6381
rect 68592 5984 68630 6381
rect 68766 6326 68800 6332
rect 68766 6298 68800 6326
rect 68766 6258 68800 6260
rect 68766 6226 68800 6258
rect 68766 6156 68800 6188
rect 68766 6154 68800 6156
rect 68766 6088 68800 6116
rect 68766 6082 68800 6088
rect 68877 6326 68911 6332
rect 68877 6298 68911 6326
rect 68877 6258 68911 6260
rect 68877 6226 68911 6258
rect 68877 6156 68911 6188
rect 68877 6154 68911 6156
rect 68877 6088 68911 6116
rect 68877 6082 68911 6088
rect 68963 6326 68997 6332
rect 68963 6298 68997 6326
rect 68963 6258 68997 6260
rect 68963 6226 68997 6258
rect 68963 6156 68997 6188
rect 68963 6154 68997 6156
rect 68963 6088 68997 6116
rect 68963 6082 68997 6088
rect 69049 6326 69083 6332
rect 69049 6298 69083 6326
rect 69049 6258 69083 6260
rect 69049 6226 69083 6258
rect 69049 6156 69083 6188
rect 69049 6154 69083 6156
rect 69049 6088 69083 6116
rect 69049 6082 69083 6088
rect 69160 6326 69194 6332
rect 69160 6298 69194 6326
rect 69160 6258 69194 6260
rect 69160 6226 69194 6258
rect 69160 6156 69194 6188
rect 69160 6154 69194 6156
rect 69160 6088 69194 6116
rect 69160 6082 69194 6088
rect 68891 5970 68895 6004
rect 68895 5970 68925 6004
rect 68963 5970 68997 6004
rect 69035 5970 69065 6004
rect 69065 5970 69069 6004
rect 69330 5984 69368 6381
rect -220 5780 -180 5820
rect -424 5458 -390 5734
rect -336 5458 -302 5734
rect -440 5356 -390 5370
rect -330 5356 -280 5370
rect -440 5320 -434 5356
rect -434 5320 -398 5356
rect -398 5320 -390 5356
rect -330 5320 -300 5356
rect -300 5320 -280 5356
<< metal1 >>
rect -3880 98790 -1880 110790
rect -3880 94300 -1870 98790
rect -610 95932 9200 97790
rect -610 95790 4192 95932
rect -610 94760 -550 95790
rect -510 95540 -220 95560
rect -510 95480 -490 95540
rect -240 95480 -220 95540
rect 4186 95535 4192 95790
rect 4230 95790 4930 95932
rect 4230 95535 4236 95790
rect 4186 95523 4236 95535
rect 4924 95535 4930 95790
rect 4968 95790 9200 95932
rect 4968 95535 4974 95790
rect 4924 95523 4974 95535
rect -510 95460 -220 95480
rect -430 95384 -384 95396
rect -430 94808 -424 95384
rect -390 94808 -384 95384
rect -430 94796 -384 94808
rect -342 95384 -296 95396
rect -342 94808 -336 95384
rect -302 94808 -296 95384
rect 4479 95364 4681 95384
rect 4479 95330 4491 95364
rect 4525 95330 4563 95364
rect 4597 95330 4635 95364
rect 4669 95330 4681 95364
rect 4479 95318 4681 95330
rect 4166 94886 4176 95318
rect 4246 94886 4256 95318
rect 4354 95252 4412 95280
rect 4354 95218 4366 95252
rect 4400 95218 4412 95252
rect 4354 95180 4412 95218
rect 4354 95146 4366 95180
rect 4400 95146 4412 95180
rect 4354 95108 4412 95146
rect 4354 95074 4366 95108
rect 4400 95074 4412 95108
rect 4354 95036 4412 95074
rect 4354 95002 4366 95036
rect 4400 95002 4412 95036
rect 4354 94974 4412 95002
rect 4468 95252 4520 95280
rect 4468 95218 4477 95252
rect 4511 95218 4520 95252
rect 4468 95180 4520 95218
rect 4468 95146 4477 95180
rect 4511 95146 4520 95180
rect 4468 95108 4520 95146
rect 4468 95096 4477 95108
rect 4511 95096 4520 95108
rect 4468 95036 4520 95044
rect 4468 95032 4477 95036
rect 4511 95032 4520 95036
rect 4468 94974 4520 94980
rect 4554 95274 4606 95280
rect 4554 95218 4563 95222
rect 4597 95218 4606 95222
rect 4554 95210 4606 95218
rect 4554 95146 4563 95158
rect 4597 95146 4606 95158
rect 4554 95108 4606 95146
rect 4554 95074 4563 95108
rect 4597 95074 4606 95108
rect 4554 95036 4606 95074
rect 4554 95002 4563 95036
rect 4597 95002 4606 95036
rect 4554 94974 4606 95002
rect 4640 95252 4692 95280
rect 4640 95218 4649 95252
rect 4683 95218 4692 95252
rect 4640 95180 4692 95218
rect 4640 95146 4649 95180
rect 4683 95146 4692 95180
rect 4640 95108 4692 95146
rect 4640 95096 4649 95108
rect 4683 95096 4692 95108
rect 4640 95036 4692 95044
rect 4640 95032 4649 95036
rect 4683 95032 4692 95036
rect 4640 94974 4692 94980
rect 4748 95252 4806 95280
rect 4748 95218 4760 95252
rect 4794 95218 4806 95252
rect 4748 95180 4806 95218
rect 4748 95146 4760 95180
rect 4794 95146 4806 95180
rect 4748 95108 4806 95146
rect 4748 95074 4760 95108
rect 4794 95074 4806 95108
rect 4748 95036 4806 95074
rect 4748 95002 4760 95036
rect 4794 95002 4806 95036
rect 4748 94974 4806 95002
rect -342 94796 -296 94808
rect 4366 94800 4400 94974
rect 4479 94924 4681 94936
rect 4479 94890 4491 94924
rect 4525 94890 4563 94924
rect 4597 94890 4635 94924
rect 4669 94890 4681 94924
rect 4479 94870 4681 94890
rect 4479 94810 4493 94870
rect 4667 94810 4681 94870
rect -610 94720 -600 94760
rect -560 94750 -550 94760
rect -240 94750 -160 94760
rect -560 94720 -430 94750
rect -610 94710 -430 94720
rect -610 94700 -550 94710
rect -240 94690 -230 94750
rect -170 94690 -160 94750
rect -240 94680 -160 94690
rect 4360 94740 4400 94800
rect 4760 94800 4794 94974
rect 4904 94886 4914 95318
rect 4984 94886 4994 95318
rect 4760 94740 4800 94800
rect -430 94654 -384 94666
rect -430 94378 -424 94654
rect -390 94378 -384 94654
rect -430 94366 -384 94378
rect -342 94654 -296 94666
rect -342 94378 -336 94654
rect -302 94378 -296 94654
rect -342 94366 -296 94378
rect -3880 94290 0 94300
rect -3880 94240 -440 94290
rect -390 94240 -330 94290
rect -280 94240 0 94290
rect -3880 94220 0 94240
rect -3880 91910 -1870 94220
rect 4360 91910 4800 94740
rect -3880 89910 9200 91910
rect -3880 84420 -1870 89910
rect -610 86052 18400 87910
rect -610 85910 4192 86052
rect -610 84880 -550 85910
rect -510 85660 -220 85680
rect -510 85600 -490 85660
rect -240 85600 -220 85660
rect 4186 85655 4192 85910
rect 4230 85910 4930 86052
rect 4230 85655 4236 85910
rect 4186 85643 4236 85655
rect 4924 85655 4930 85910
rect 4968 85910 13392 86052
rect 4968 85655 4974 85910
rect 4924 85643 4974 85655
rect 13386 85655 13392 85910
rect 13430 85910 14130 86052
rect 13430 85655 13436 85910
rect 13386 85643 13436 85655
rect 14124 85655 14130 85910
rect 14168 85910 18400 86052
rect 14168 85655 14174 85910
rect 14124 85643 14174 85655
rect -510 85580 -220 85600
rect -430 85504 -384 85516
rect -430 84928 -424 85504
rect -390 84928 -384 85504
rect -430 84916 -384 84928
rect -342 85504 -296 85516
rect -342 84928 -336 85504
rect -302 84928 -296 85504
rect 4479 85484 4681 85504
rect 4479 85450 4491 85484
rect 4525 85450 4563 85484
rect 4597 85450 4635 85484
rect 4669 85450 4681 85484
rect 4479 85438 4681 85450
rect 13679 85484 13881 85504
rect 13679 85450 13691 85484
rect 13725 85450 13763 85484
rect 13797 85450 13835 85484
rect 13869 85450 13881 85484
rect 13679 85438 13881 85450
rect 4166 85006 4176 85438
rect 4246 85006 4256 85438
rect 4354 85372 4412 85400
rect 4354 85338 4366 85372
rect 4400 85338 4412 85372
rect 4354 85300 4412 85338
rect 4354 85266 4366 85300
rect 4400 85266 4412 85300
rect 4354 85228 4412 85266
rect 4354 85194 4366 85228
rect 4400 85194 4412 85228
rect 4354 85156 4412 85194
rect 4354 85122 4366 85156
rect 4400 85122 4412 85156
rect 4354 85094 4412 85122
rect 4468 85372 4520 85400
rect 4468 85338 4477 85372
rect 4511 85338 4520 85372
rect 4468 85300 4520 85338
rect 4468 85266 4477 85300
rect 4511 85266 4520 85300
rect 4468 85228 4520 85266
rect 4468 85216 4477 85228
rect 4511 85216 4520 85228
rect 4468 85156 4520 85164
rect 4468 85152 4477 85156
rect 4511 85152 4520 85156
rect 4468 85094 4520 85100
rect 4554 85394 4606 85400
rect 4554 85338 4563 85342
rect 4597 85338 4606 85342
rect 4554 85330 4606 85338
rect 4554 85266 4563 85278
rect 4597 85266 4606 85278
rect 4554 85228 4606 85266
rect 4554 85194 4563 85228
rect 4597 85194 4606 85228
rect 4554 85156 4606 85194
rect 4554 85122 4563 85156
rect 4597 85122 4606 85156
rect 4554 85094 4606 85122
rect 4640 85372 4692 85400
rect 4640 85338 4649 85372
rect 4683 85338 4692 85372
rect 4640 85300 4692 85338
rect 4640 85266 4649 85300
rect 4683 85266 4692 85300
rect 4640 85228 4692 85266
rect 4640 85216 4649 85228
rect 4683 85216 4692 85228
rect 4640 85156 4692 85164
rect 4640 85152 4649 85156
rect 4683 85152 4692 85156
rect 4640 85094 4692 85100
rect 4748 85372 4806 85400
rect 4748 85338 4760 85372
rect 4794 85338 4806 85372
rect 4748 85300 4806 85338
rect 4748 85266 4760 85300
rect 4794 85266 4806 85300
rect 4748 85228 4806 85266
rect 4748 85194 4760 85228
rect 4794 85194 4806 85228
rect 4748 85156 4806 85194
rect 4748 85122 4760 85156
rect 4794 85122 4806 85156
rect 4748 85094 4806 85122
rect -342 84916 -296 84928
rect 4366 84920 4400 85094
rect 4479 85044 4681 85056
rect 4479 85010 4491 85044
rect 4525 85010 4563 85044
rect 4597 85010 4635 85044
rect 4669 85010 4681 85044
rect 4479 84990 4681 85010
rect 4479 84930 4493 84990
rect 4667 84930 4681 84990
rect -610 84840 -600 84880
rect -560 84870 -550 84880
rect -240 84870 -160 84880
rect -560 84840 -430 84870
rect -610 84830 -430 84840
rect -610 84820 -550 84830
rect -240 84810 -230 84870
rect -170 84810 -160 84870
rect -240 84800 -160 84810
rect 4360 84860 4400 84920
rect 4760 84920 4794 85094
rect 4904 85006 4914 85438
rect 4984 85006 4994 85438
rect 13366 85006 13376 85438
rect 13446 85006 13456 85438
rect 13554 85372 13612 85400
rect 13554 85338 13566 85372
rect 13600 85338 13612 85372
rect 13554 85300 13612 85338
rect 13554 85266 13566 85300
rect 13600 85266 13612 85300
rect 13554 85228 13612 85266
rect 13554 85194 13566 85228
rect 13600 85194 13612 85228
rect 13554 85156 13612 85194
rect 13554 85122 13566 85156
rect 13600 85122 13612 85156
rect 13554 85094 13612 85122
rect 13668 85372 13720 85400
rect 13668 85338 13677 85372
rect 13711 85338 13720 85372
rect 13668 85300 13720 85338
rect 13668 85266 13677 85300
rect 13711 85266 13720 85300
rect 13668 85228 13720 85266
rect 13668 85216 13677 85228
rect 13711 85216 13720 85228
rect 13668 85156 13720 85164
rect 13668 85152 13677 85156
rect 13711 85152 13720 85156
rect 13668 85094 13720 85100
rect 13754 85394 13806 85400
rect 13754 85338 13763 85342
rect 13797 85338 13806 85342
rect 13754 85330 13806 85338
rect 13754 85266 13763 85278
rect 13797 85266 13806 85278
rect 13754 85228 13806 85266
rect 13754 85194 13763 85228
rect 13797 85194 13806 85228
rect 13754 85156 13806 85194
rect 13754 85122 13763 85156
rect 13797 85122 13806 85156
rect 13754 85094 13806 85122
rect 13840 85372 13892 85400
rect 13840 85338 13849 85372
rect 13883 85338 13892 85372
rect 13840 85300 13892 85338
rect 13840 85266 13849 85300
rect 13883 85266 13892 85300
rect 13840 85228 13892 85266
rect 13840 85216 13849 85228
rect 13883 85216 13892 85228
rect 13840 85156 13892 85164
rect 13840 85152 13849 85156
rect 13883 85152 13892 85156
rect 13840 85094 13892 85100
rect 13948 85372 14006 85400
rect 13948 85338 13960 85372
rect 13994 85338 14006 85372
rect 13948 85300 14006 85338
rect 13948 85266 13960 85300
rect 13994 85266 14006 85300
rect 13948 85228 14006 85266
rect 13948 85194 13960 85228
rect 13994 85194 14006 85228
rect 13948 85156 14006 85194
rect 13948 85122 13960 85156
rect 13994 85122 14006 85156
rect 13948 85094 14006 85122
rect 13566 84920 13600 85094
rect 13679 85044 13881 85056
rect 13679 85010 13691 85044
rect 13725 85010 13763 85044
rect 13797 85010 13835 85044
rect 13869 85010 13881 85044
rect 13679 84990 13881 85010
rect 13679 84930 13693 84990
rect 13867 84930 13881 84990
rect 4760 84860 4800 84920
rect -430 84774 -384 84786
rect -430 84498 -424 84774
rect -390 84498 -384 84774
rect -430 84486 -384 84498
rect -342 84774 -296 84786
rect -342 84498 -336 84774
rect -302 84498 -296 84774
rect -342 84486 -296 84498
rect -3880 84410 0 84420
rect -3880 84360 -440 84410
rect -390 84360 -330 84410
rect -280 84360 0 84410
rect -3880 84340 0 84360
rect -3880 82030 -1870 84340
rect 4360 82030 4800 84860
rect 13560 84860 13600 84920
rect 13960 84920 13994 85094
rect 14104 85006 14114 85438
rect 14184 85006 14194 85438
rect 13960 84860 14000 84920
rect 13560 82030 14000 84860
rect -3880 80030 18400 82030
rect -3880 74540 -1870 80030
rect -610 76172 36800 78030
rect -610 76030 4192 76172
rect -610 75000 -550 76030
rect -510 75780 -220 75800
rect -510 75720 -490 75780
rect -240 75720 -220 75780
rect 4186 75775 4192 76030
rect 4230 76030 4930 76172
rect 4230 75775 4236 76030
rect 4186 75763 4236 75775
rect 4924 75775 4930 76030
rect 4968 76030 13392 76172
rect 4968 75775 4974 76030
rect 4924 75763 4974 75775
rect 13386 75775 13392 76030
rect 13430 76030 14130 76172
rect 13430 75775 13436 76030
rect 13386 75763 13436 75775
rect 14124 75775 14130 76030
rect 14168 76030 22592 76172
rect 14168 75775 14174 76030
rect 14124 75763 14174 75775
rect 22586 75775 22592 76030
rect 22630 76030 23330 76172
rect 22630 75775 22636 76030
rect 22586 75763 22636 75775
rect 23324 75775 23330 76030
rect 23368 76030 31792 76172
rect 23368 75775 23374 76030
rect 23324 75763 23374 75775
rect 31786 75775 31792 76030
rect 31830 76030 32530 76172
rect 31830 75775 31836 76030
rect 31786 75763 31836 75775
rect 32524 75775 32530 76030
rect 32568 76030 36800 76172
rect 32568 75775 32574 76030
rect 32524 75763 32574 75775
rect -510 75700 -220 75720
rect -430 75624 -384 75636
rect -430 75048 -424 75624
rect -390 75048 -384 75624
rect -430 75036 -384 75048
rect -342 75624 -296 75636
rect -342 75048 -336 75624
rect -302 75048 -296 75624
rect 4479 75604 4681 75624
rect 4479 75570 4491 75604
rect 4525 75570 4563 75604
rect 4597 75570 4635 75604
rect 4669 75570 4681 75604
rect 4479 75558 4681 75570
rect 13679 75604 13881 75624
rect 13679 75570 13691 75604
rect 13725 75570 13763 75604
rect 13797 75570 13835 75604
rect 13869 75570 13881 75604
rect 13679 75558 13881 75570
rect 22879 75604 23081 75624
rect 22879 75570 22891 75604
rect 22925 75570 22963 75604
rect 22997 75570 23035 75604
rect 23069 75570 23081 75604
rect 22879 75558 23081 75570
rect 32079 75604 32281 75624
rect 32079 75570 32091 75604
rect 32125 75570 32163 75604
rect 32197 75570 32235 75604
rect 32269 75570 32281 75604
rect 32079 75558 32281 75570
rect 4166 75126 4176 75558
rect 4246 75126 4256 75558
rect 4354 75492 4412 75520
rect 4354 75458 4366 75492
rect 4400 75458 4412 75492
rect 4354 75420 4412 75458
rect 4354 75386 4366 75420
rect 4400 75386 4412 75420
rect 4354 75348 4412 75386
rect 4354 75314 4366 75348
rect 4400 75314 4412 75348
rect 4354 75276 4412 75314
rect 4354 75242 4366 75276
rect 4400 75242 4412 75276
rect 4354 75214 4412 75242
rect 4468 75492 4520 75520
rect 4468 75458 4477 75492
rect 4511 75458 4520 75492
rect 4468 75420 4520 75458
rect 4468 75386 4477 75420
rect 4511 75386 4520 75420
rect 4468 75348 4520 75386
rect 4468 75336 4477 75348
rect 4511 75336 4520 75348
rect 4468 75276 4520 75284
rect 4468 75272 4477 75276
rect 4511 75272 4520 75276
rect 4468 75214 4520 75220
rect 4554 75514 4606 75520
rect 4554 75458 4563 75462
rect 4597 75458 4606 75462
rect 4554 75450 4606 75458
rect 4554 75386 4563 75398
rect 4597 75386 4606 75398
rect 4554 75348 4606 75386
rect 4554 75314 4563 75348
rect 4597 75314 4606 75348
rect 4554 75276 4606 75314
rect 4554 75242 4563 75276
rect 4597 75242 4606 75276
rect 4554 75214 4606 75242
rect 4640 75492 4692 75520
rect 4640 75458 4649 75492
rect 4683 75458 4692 75492
rect 4640 75420 4692 75458
rect 4640 75386 4649 75420
rect 4683 75386 4692 75420
rect 4640 75348 4692 75386
rect 4640 75336 4649 75348
rect 4683 75336 4692 75348
rect 4640 75276 4692 75284
rect 4640 75272 4649 75276
rect 4683 75272 4692 75276
rect 4640 75214 4692 75220
rect 4748 75492 4806 75520
rect 4748 75458 4760 75492
rect 4794 75458 4806 75492
rect 4748 75420 4806 75458
rect 4748 75386 4760 75420
rect 4794 75386 4806 75420
rect 4748 75348 4806 75386
rect 4748 75314 4760 75348
rect 4794 75314 4806 75348
rect 4748 75276 4806 75314
rect 4748 75242 4760 75276
rect 4794 75242 4806 75276
rect 4748 75214 4806 75242
rect -342 75036 -296 75048
rect 4366 75040 4400 75214
rect 4479 75164 4681 75176
rect 4479 75130 4491 75164
rect 4525 75130 4563 75164
rect 4597 75130 4635 75164
rect 4669 75130 4681 75164
rect 4479 75110 4681 75130
rect 4479 75050 4493 75110
rect 4667 75050 4681 75110
rect -610 74960 -600 75000
rect -560 74990 -550 75000
rect -240 74990 -160 75000
rect -560 74960 -430 74990
rect -610 74950 -430 74960
rect -610 74940 -550 74950
rect -240 74930 -230 74990
rect -170 74930 -160 74990
rect -240 74920 -160 74930
rect 4360 74980 4400 75040
rect 4760 75040 4794 75214
rect 4904 75126 4914 75558
rect 4984 75126 4994 75558
rect 13366 75126 13376 75558
rect 13446 75126 13456 75558
rect 13554 75492 13612 75520
rect 13554 75458 13566 75492
rect 13600 75458 13612 75492
rect 13554 75420 13612 75458
rect 13554 75386 13566 75420
rect 13600 75386 13612 75420
rect 13554 75348 13612 75386
rect 13554 75314 13566 75348
rect 13600 75314 13612 75348
rect 13554 75276 13612 75314
rect 13554 75242 13566 75276
rect 13600 75242 13612 75276
rect 13554 75214 13612 75242
rect 13668 75492 13720 75520
rect 13668 75458 13677 75492
rect 13711 75458 13720 75492
rect 13668 75420 13720 75458
rect 13668 75386 13677 75420
rect 13711 75386 13720 75420
rect 13668 75348 13720 75386
rect 13668 75336 13677 75348
rect 13711 75336 13720 75348
rect 13668 75276 13720 75284
rect 13668 75272 13677 75276
rect 13711 75272 13720 75276
rect 13668 75214 13720 75220
rect 13754 75514 13806 75520
rect 13754 75458 13763 75462
rect 13797 75458 13806 75462
rect 13754 75450 13806 75458
rect 13754 75386 13763 75398
rect 13797 75386 13806 75398
rect 13754 75348 13806 75386
rect 13754 75314 13763 75348
rect 13797 75314 13806 75348
rect 13754 75276 13806 75314
rect 13754 75242 13763 75276
rect 13797 75242 13806 75276
rect 13754 75214 13806 75242
rect 13840 75492 13892 75520
rect 13840 75458 13849 75492
rect 13883 75458 13892 75492
rect 13840 75420 13892 75458
rect 13840 75386 13849 75420
rect 13883 75386 13892 75420
rect 13840 75348 13892 75386
rect 13840 75336 13849 75348
rect 13883 75336 13892 75348
rect 13840 75276 13892 75284
rect 13840 75272 13849 75276
rect 13883 75272 13892 75276
rect 13840 75214 13892 75220
rect 13948 75492 14006 75520
rect 13948 75458 13960 75492
rect 13994 75458 14006 75492
rect 13948 75420 14006 75458
rect 13948 75386 13960 75420
rect 13994 75386 14006 75420
rect 13948 75348 14006 75386
rect 13948 75314 13960 75348
rect 13994 75314 14006 75348
rect 13948 75276 14006 75314
rect 13948 75242 13960 75276
rect 13994 75242 14006 75276
rect 13948 75214 14006 75242
rect 13566 75040 13600 75214
rect 13679 75164 13881 75176
rect 13679 75130 13691 75164
rect 13725 75130 13763 75164
rect 13797 75130 13835 75164
rect 13869 75130 13881 75164
rect 13679 75110 13881 75130
rect 13679 75050 13693 75110
rect 13867 75050 13881 75110
rect 4760 74980 4800 75040
rect -430 74894 -384 74906
rect -430 74618 -424 74894
rect -390 74618 -384 74894
rect -430 74606 -384 74618
rect -342 74894 -296 74906
rect -342 74618 -336 74894
rect -302 74618 -296 74894
rect -342 74606 -296 74618
rect -3880 74530 0 74540
rect -3880 74480 -440 74530
rect -390 74480 -330 74530
rect -280 74480 0 74530
rect -3880 74460 0 74480
rect -3880 72150 -1870 74460
rect 4360 72150 4800 74980
rect 13560 74980 13600 75040
rect 13960 75040 13994 75214
rect 14104 75126 14114 75558
rect 14184 75126 14194 75558
rect 22566 75126 22576 75558
rect 22646 75126 22656 75558
rect 22754 75492 22812 75520
rect 22754 75458 22766 75492
rect 22800 75458 22812 75492
rect 22754 75420 22812 75458
rect 22754 75386 22766 75420
rect 22800 75386 22812 75420
rect 22754 75348 22812 75386
rect 22754 75314 22766 75348
rect 22800 75314 22812 75348
rect 22754 75276 22812 75314
rect 22754 75242 22766 75276
rect 22800 75242 22812 75276
rect 22754 75214 22812 75242
rect 22868 75492 22920 75520
rect 22868 75458 22877 75492
rect 22911 75458 22920 75492
rect 22868 75420 22920 75458
rect 22868 75386 22877 75420
rect 22911 75386 22920 75420
rect 22868 75348 22920 75386
rect 22868 75336 22877 75348
rect 22911 75336 22920 75348
rect 22868 75276 22920 75284
rect 22868 75272 22877 75276
rect 22911 75272 22920 75276
rect 22868 75214 22920 75220
rect 22954 75514 23006 75520
rect 22954 75458 22963 75462
rect 22997 75458 23006 75462
rect 22954 75450 23006 75458
rect 22954 75386 22963 75398
rect 22997 75386 23006 75398
rect 22954 75348 23006 75386
rect 22954 75314 22963 75348
rect 22997 75314 23006 75348
rect 22954 75276 23006 75314
rect 22954 75242 22963 75276
rect 22997 75242 23006 75276
rect 22954 75214 23006 75242
rect 23040 75492 23092 75520
rect 23040 75458 23049 75492
rect 23083 75458 23092 75492
rect 23040 75420 23092 75458
rect 23040 75386 23049 75420
rect 23083 75386 23092 75420
rect 23040 75348 23092 75386
rect 23040 75336 23049 75348
rect 23083 75336 23092 75348
rect 23040 75276 23092 75284
rect 23040 75272 23049 75276
rect 23083 75272 23092 75276
rect 23040 75214 23092 75220
rect 23148 75492 23206 75520
rect 23148 75458 23160 75492
rect 23194 75458 23206 75492
rect 23148 75420 23206 75458
rect 23148 75386 23160 75420
rect 23194 75386 23206 75420
rect 23148 75348 23206 75386
rect 23148 75314 23160 75348
rect 23194 75314 23206 75348
rect 23148 75276 23206 75314
rect 23148 75242 23160 75276
rect 23194 75242 23206 75276
rect 23148 75214 23206 75242
rect 22766 75040 22800 75214
rect 22879 75164 23081 75176
rect 22879 75130 22891 75164
rect 22925 75130 22963 75164
rect 22997 75130 23035 75164
rect 23069 75130 23081 75164
rect 22879 75110 23081 75130
rect 22879 75050 22893 75110
rect 23067 75050 23081 75110
rect 13960 74980 14000 75040
rect 13560 72150 14000 74980
rect 22760 74980 22800 75040
rect 23160 75040 23194 75214
rect 23304 75126 23314 75558
rect 23384 75126 23394 75558
rect 31766 75126 31776 75558
rect 31846 75126 31856 75558
rect 31954 75492 32012 75520
rect 31954 75458 31966 75492
rect 32000 75458 32012 75492
rect 31954 75420 32012 75458
rect 31954 75386 31966 75420
rect 32000 75386 32012 75420
rect 31954 75348 32012 75386
rect 31954 75314 31966 75348
rect 32000 75314 32012 75348
rect 31954 75276 32012 75314
rect 31954 75242 31966 75276
rect 32000 75242 32012 75276
rect 31954 75214 32012 75242
rect 32068 75492 32120 75520
rect 32068 75458 32077 75492
rect 32111 75458 32120 75492
rect 32068 75420 32120 75458
rect 32068 75386 32077 75420
rect 32111 75386 32120 75420
rect 32068 75348 32120 75386
rect 32068 75336 32077 75348
rect 32111 75336 32120 75348
rect 32068 75276 32120 75284
rect 32068 75272 32077 75276
rect 32111 75272 32120 75276
rect 32068 75214 32120 75220
rect 32154 75514 32206 75520
rect 32154 75458 32163 75462
rect 32197 75458 32206 75462
rect 32154 75450 32206 75458
rect 32154 75386 32163 75398
rect 32197 75386 32206 75398
rect 32154 75348 32206 75386
rect 32154 75314 32163 75348
rect 32197 75314 32206 75348
rect 32154 75276 32206 75314
rect 32154 75242 32163 75276
rect 32197 75242 32206 75276
rect 32154 75214 32206 75242
rect 32240 75492 32292 75520
rect 32240 75458 32249 75492
rect 32283 75458 32292 75492
rect 32240 75420 32292 75458
rect 32240 75386 32249 75420
rect 32283 75386 32292 75420
rect 32240 75348 32292 75386
rect 32240 75336 32249 75348
rect 32283 75336 32292 75348
rect 32240 75276 32292 75284
rect 32240 75272 32249 75276
rect 32283 75272 32292 75276
rect 32240 75214 32292 75220
rect 32348 75492 32406 75520
rect 32348 75458 32360 75492
rect 32394 75458 32406 75492
rect 32348 75420 32406 75458
rect 32348 75386 32360 75420
rect 32394 75386 32406 75420
rect 32348 75348 32406 75386
rect 32348 75314 32360 75348
rect 32394 75314 32406 75348
rect 32348 75276 32406 75314
rect 32348 75242 32360 75276
rect 32394 75242 32406 75276
rect 32348 75214 32406 75242
rect 31966 75040 32000 75214
rect 32079 75164 32281 75176
rect 32079 75130 32091 75164
rect 32125 75130 32163 75164
rect 32197 75130 32235 75164
rect 32269 75130 32281 75164
rect 32079 75110 32281 75130
rect 32079 75050 32093 75110
rect 32267 75050 32281 75110
rect 23160 74980 23200 75040
rect 22760 72150 23200 74980
rect 31960 74980 32000 75040
rect 32360 75040 32394 75214
rect 32504 75126 32514 75558
rect 32584 75126 32594 75558
rect 32360 74980 32400 75040
rect 31960 72150 32400 74980
rect -3880 70150 36800 72150
rect -3880 64660 -1870 70150
rect -610 66292 73600 68150
rect -610 66150 4192 66292
rect -610 65120 -550 66150
rect -510 65900 -220 65920
rect -510 65840 -490 65900
rect -240 65840 -220 65900
rect 4186 65895 4192 66150
rect 4230 66150 4930 66292
rect 4230 65895 4236 66150
rect 4186 65883 4236 65895
rect 4924 65895 4930 66150
rect 4968 66150 13392 66292
rect 4968 65895 4974 66150
rect 4924 65883 4974 65895
rect 13386 65895 13392 66150
rect 13430 66150 14130 66292
rect 13430 65895 13436 66150
rect 13386 65883 13436 65895
rect 14124 65895 14130 66150
rect 14168 66150 22592 66292
rect 14168 65895 14174 66150
rect 14124 65883 14174 65895
rect 22586 65895 22592 66150
rect 22630 66150 23330 66292
rect 22630 65895 22636 66150
rect 22586 65883 22636 65895
rect 23324 65895 23330 66150
rect 23368 66150 31792 66292
rect 23368 65895 23374 66150
rect 23324 65883 23374 65895
rect 31786 65895 31792 66150
rect 31830 66150 32530 66292
rect 31830 65895 31836 66150
rect 31786 65883 31836 65895
rect 32524 65895 32530 66150
rect 32568 66150 40992 66292
rect 32568 65895 32574 66150
rect 32524 65883 32574 65895
rect 40986 65895 40992 66150
rect 41030 66150 41730 66292
rect 41030 65895 41036 66150
rect 40986 65883 41036 65895
rect 41724 65895 41730 66150
rect 41768 66150 50192 66292
rect 41768 65895 41774 66150
rect 41724 65883 41774 65895
rect 50186 65895 50192 66150
rect 50230 66150 50930 66292
rect 50230 65895 50236 66150
rect 50186 65883 50236 65895
rect 50924 65895 50930 66150
rect 50968 66150 59392 66292
rect 50968 65895 50974 66150
rect 50924 65883 50974 65895
rect 59386 65895 59392 66150
rect 59430 66150 60130 66292
rect 59430 65895 59436 66150
rect 59386 65883 59436 65895
rect 60124 65895 60130 66150
rect 60168 66150 68592 66292
rect 60168 65895 60174 66150
rect 60124 65883 60174 65895
rect 68586 65895 68592 66150
rect 68630 66150 69330 66292
rect 68630 65895 68636 66150
rect 68586 65883 68636 65895
rect 69324 65895 69330 66150
rect 69368 66150 73600 66292
rect 69368 65895 69374 66150
rect 69324 65883 69374 65895
rect -510 65820 -220 65840
rect -430 65744 -384 65756
rect -430 65168 -424 65744
rect -390 65168 -384 65744
rect -430 65156 -384 65168
rect -342 65744 -296 65756
rect -342 65168 -336 65744
rect -302 65168 -296 65744
rect 4479 65724 4681 65744
rect 4479 65690 4491 65724
rect 4525 65690 4563 65724
rect 4597 65690 4635 65724
rect 4669 65690 4681 65724
rect 4479 65678 4681 65690
rect 13679 65724 13881 65744
rect 13679 65690 13691 65724
rect 13725 65690 13763 65724
rect 13797 65690 13835 65724
rect 13869 65690 13881 65724
rect 13679 65678 13881 65690
rect 22879 65724 23081 65744
rect 22879 65690 22891 65724
rect 22925 65690 22963 65724
rect 22997 65690 23035 65724
rect 23069 65690 23081 65724
rect 22879 65678 23081 65690
rect 32079 65724 32281 65744
rect 32079 65690 32091 65724
rect 32125 65690 32163 65724
rect 32197 65690 32235 65724
rect 32269 65690 32281 65724
rect 32079 65678 32281 65690
rect 41279 65724 41481 65744
rect 41279 65690 41291 65724
rect 41325 65690 41363 65724
rect 41397 65690 41435 65724
rect 41469 65690 41481 65724
rect 41279 65678 41481 65690
rect 50479 65724 50681 65744
rect 50479 65690 50491 65724
rect 50525 65690 50563 65724
rect 50597 65690 50635 65724
rect 50669 65690 50681 65724
rect 50479 65678 50681 65690
rect 59679 65724 59881 65744
rect 59679 65690 59691 65724
rect 59725 65690 59763 65724
rect 59797 65690 59835 65724
rect 59869 65690 59881 65724
rect 59679 65678 59881 65690
rect 68879 65724 69081 65744
rect 68879 65690 68891 65724
rect 68925 65690 68963 65724
rect 68997 65690 69035 65724
rect 69069 65690 69081 65724
rect 68879 65678 69081 65690
rect 4166 65246 4176 65678
rect 4246 65246 4256 65678
rect 4354 65612 4412 65640
rect 4354 65578 4366 65612
rect 4400 65578 4412 65612
rect 4354 65540 4412 65578
rect 4354 65506 4366 65540
rect 4400 65506 4412 65540
rect 4354 65468 4412 65506
rect 4354 65434 4366 65468
rect 4400 65434 4412 65468
rect 4354 65396 4412 65434
rect 4354 65362 4366 65396
rect 4400 65362 4412 65396
rect 4354 65334 4412 65362
rect 4468 65612 4520 65640
rect 4468 65578 4477 65612
rect 4511 65578 4520 65612
rect 4468 65540 4520 65578
rect 4468 65506 4477 65540
rect 4511 65506 4520 65540
rect 4468 65468 4520 65506
rect 4468 65456 4477 65468
rect 4511 65456 4520 65468
rect 4468 65396 4520 65404
rect 4468 65392 4477 65396
rect 4511 65392 4520 65396
rect 4468 65334 4520 65340
rect 4554 65634 4606 65640
rect 4554 65578 4563 65582
rect 4597 65578 4606 65582
rect 4554 65570 4606 65578
rect 4554 65506 4563 65518
rect 4597 65506 4606 65518
rect 4554 65468 4606 65506
rect 4554 65434 4563 65468
rect 4597 65434 4606 65468
rect 4554 65396 4606 65434
rect 4554 65362 4563 65396
rect 4597 65362 4606 65396
rect 4554 65334 4606 65362
rect 4640 65612 4692 65640
rect 4640 65578 4649 65612
rect 4683 65578 4692 65612
rect 4640 65540 4692 65578
rect 4640 65506 4649 65540
rect 4683 65506 4692 65540
rect 4640 65468 4692 65506
rect 4640 65456 4649 65468
rect 4683 65456 4692 65468
rect 4640 65396 4692 65404
rect 4640 65392 4649 65396
rect 4683 65392 4692 65396
rect 4640 65334 4692 65340
rect 4748 65612 4806 65640
rect 4748 65578 4760 65612
rect 4794 65578 4806 65612
rect 4748 65540 4806 65578
rect 4748 65506 4760 65540
rect 4794 65506 4806 65540
rect 4748 65468 4806 65506
rect 4748 65434 4760 65468
rect 4794 65434 4806 65468
rect 4748 65396 4806 65434
rect 4748 65362 4760 65396
rect 4794 65362 4806 65396
rect 4748 65334 4806 65362
rect -342 65156 -296 65168
rect 4366 65160 4400 65334
rect 4479 65284 4681 65296
rect 4479 65250 4491 65284
rect 4525 65250 4563 65284
rect 4597 65250 4635 65284
rect 4669 65250 4681 65284
rect 4479 65230 4681 65250
rect 4479 65170 4493 65230
rect 4667 65170 4681 65230
rect -610 65080 -600 65120
rect -560 65110 -550 65120
rect -240 65110 -160 65120
rect -560 65080 -430 65110
rect -610 65070 -430 65080
rect -610 65060 -550 65070
rect -240 65050 -230 65110
rect -170 65050 -160 65110
rect -240 65040 -160 65050
rect 4360 65100 4400 65160
rect 4760 65160 4794 65334
rect 4904 65246 4914 65678
rect 4984 65246 4994 65678
rect 13366 65246 13376 65678
rect 13446 65246 13456 65678
rect 13554 65612 13612 65640
rect 13554 65578 13566 65612
rect 13600 65578 13612 65612
rect 13554 65540 13612 65578
rect 13554 65506 13566 65540
rect 13600 65506 13612 65540
rect 13554 65468 13612 65506
rect 13554 65434 13566 65468
rect 13600 65434 13612 65468
rect 13554 65396 13612 65434
rect 13554 65362 13566 65396
rect 13600 65362 13612 65396
rect 13554 65334 13612 65362
rect 13668 65612 13720 65640
rect 13668 65578 13677 65612
rect 13711 65578 13720 65612
rect 13668 65540 13720 65578
rect 13668 65506 13677 65540
rect 13711 65506 13720 65540
rect 13668 65468 13720 65506
rect 13668 65456 13677 65468
rect 13711 65456 13720 65468
rect 13668 65396 13720 65404
rect 13668 65392 13677 65396
rect 13711 65392 13720 65396
rect 13668 65334 13720 65340
rect 13754 65634 13806 65640
rect 13754 65578 13763 65582
rect 13797 65578 13806 65582
rect 13754 65570 13806 65578
rect 13754 65506 13763 65518
rect 13797 65506 13806 65518
rect 13754 65468 13806 65506
rect 13754 65434 13763 65468
rect 13797 65434 13806 65468
rect 13754 65396 13806 65434
rect 13754 65362 13763 65396
rect 13797 65362 13806 65396
rect 13754 65334 13806 65362
rect 13840 65612 13892 65640
rect 13840 65578 13849 65612
rect 13883 65578 13892 65612
rect 13840 65540 13892 65578
rect 13840 65506 13849 65540
rect 13883 65506 13892 65540
rect 13840 65468 13892 65506
rect 13840 65456 13849 65468
rect 13883 65456 13892 65468
rect 13840 65396 13892 65404
rect 13840 65392 13849 65396
rect 13883 65392 13892 65396
rect 13840 65334 13892 65340
rect 13948 65612 14006 65640
rect 13948 65578 13960 65612
rect 13994 65578 14006 65612
rect 13948 65540 14006 65578
rect 13948 65506 13960 65540
rect 13994 65506 14006 65540
rect 13948 65468 14006 65506
rect 13948 65434 13960 65468
rect 13994 65434 14006 65468
rect 13948 65396 14006 65434
rect 13948 65362 13960 65396
rect 13994 65362 14006 65396
rect 13948 65334 14006 65362
rect 13566 65160 13600 65334
rect 13679 65284 13881 65296
rect 13679 65250 13691 65284
rect 13725 65250 13763 65284
rect 13797 65250 13835 65284
rect 13869 65250 13881 65284
rect 13679 65230 13881 65250
rect 13679 65170 13693 65230
rect 13867 65170 13881 65230
rect 4760 65100 4800 65160
rect -430 65014 -384 65026
rect -430 64738 -424 65014
rect -390 64738 -384 65014
rect -430 64726 -384 64738
rect -342 65014 -296 65026
rect -342 64738 -336 65014
rect -302 64738 -296 65014
rect -342 64726 -296 64738
rect -3880 64650 0 64660
rect -3880 64600 -440 64650
rect -390 64600 -330 64650
rect -280 64600 0 64650
rect -3880 64580 0 64600
rect -3880 62270 -1870 64580
rect 4360 62270 4800 65100
rect 13560 65100 13600 65160
rect 13960 65160 13994 65334
rect 14104 65246 14114 65678
rect 14184 65246 14194 65678
rect 22566 65246 22576 65678
rect 22646 65246 22656 65678
rect 22754 65612 22812 65640
rect 22754 65578 22766 65612
rect 22800 65578 22812 65612
rect 22754 65540 22812 65578
rect 22754 65506 22766 65540
rect 22800 65506 22812 65540
rect 22754 65468 22812 65506
rect 22754 65434 22766 65468
rect 22800 65434 22812 65468
rect 22754 65396 22812 65434
rect 22754 65362 22766 65396
rect 22800 65362 22812 65396
rect 22754 65334 22812 65362
rect 22868 65612 22920 65640
rect 22868 65578 22877 65612
rect 22911 65578 22920 65612
rect 22868 65540 22920 65578
rect 22868 65506 22877 65540
rect 22911 65506 22920 65540
rect 22868 65468 22920 65506
rect 22868 65456 22877 65468
rect 22911 65456 22920 65468
rect 22868 65396 22920 65404
rect 22868 65392 22877 65396
rect 22911 65392 22920 65396
rect 22868 65334 22920 65340
rect 22954 65634 23006 65640
rect 22954 65578 22963 65582
rect 22997 65578 23006 65582
rect 22954 65570 23006 65578
rect 22954 65506 22963 65518
rect 22997 65506 23006 65518
rect 22954 65468 23006 65506
rect 22954 65434 22963 65468
rect 22997 65434 23006 65468
rect 22954 65396 23006 65434
rect 22954 65362 22963 65396
rect 22997 65362 23006 65396
rect 22954 65334 23006 65362
rect 23040 65612 23092 65640
rect 23040 65578 23049 65612
rect 23083 65578 23092 65612
rect 23040 65540 23092 65578
rect 23040 65506 23049 65540
rect 23083 65506 23092 65540
rect 23040 65468 23092 65506
rect 23040 65456 23049 65468
rect 23083 65456 23092 65468
rect 23040 65396 23092 65404
rect 23040 65392 23049 65396
rect 23083 65392 23092 65396
rect 23040 65334 23092 65340
rect 23148 65612 23206 65640
rect 23148 65578 23160 65612
rect 23194 65578 23206 65612
rect 23148 65540 23206 65578
rect 23148 65506 23160 65540
rect 23194 65506 23206 65540
rect 23148 65468 23206 65506
rect 23148 65434 23160 65468
rect 23194 65434 23206 65468
rect 23148 65396 23206 65434
rect 23148 65362 23160 65396
rect 23194 65362 23206 65396
rect 23148 65334 23206 65362
rect 22766 65160 22800 65334
rect 22879 65284 23081 65296
rect 22879 65250 22891 65284
rect 22925 65250 22963 65284
rect 22997 65250 23035 65284
rect 23069 65250 23081 65284
rect 22879 65230 23081 65250
rect 22879 65170 22893 65230
rect 23067 65170 23081 65230
rect 13960 65100 14000 65160
rect 13560 62270 14000 65100
rect 22760 65100 22800 65160
rect 23160 65160 23194 65334
rect 23304 65246 23314 65678
rect 23384 65246 23394 65678
rect 31766 65246 31776 65678
rect 31846 65246 31856 65678
rect 31954 65612 32012 65640
rect 31954 65578 31966 65612
rect 32000 65578 32012 65612
rect 31954 65540 32012 65578
rect 31954 65506 31966 65540
rect 32000 65506 32012 65540
rect 31954 65468 32012 65506
rect 31954 65434 31966 65468
rect 32000 65434 32012 65468
rect 31954 65396 32012 65434
rect 31954 65362 31966 65396
rect 32000 65362 32012 65396
rect 31954 65334 32012 65362
rect 32068 65612 32120 65640
rect 32068 65578 32077 65612
rect 32111 65578 32120 65612
rect 32068 65540 32120 65578
rect 32068 65506 32077 65540
rect 32111 65506 32120 65540
rect 32068 65468 32120 65506
rect 32068 65456 32077 65468
rect 32111 65456 32120 65468
rect 32068 65396 32120 65404
rect 32068 65392 32077 65396
rect 32111 65392 32120 65396
rect 32068 65334 32120 65340
rect 32154 65634 32206 65640
rect 32154 65578 32163 65582
rect 32197 65578 32206 65582
rect 32154 65570 32206 65578
rect 32154 65506 32163 65518
rect 32197 65506 32206 65518
rect 32154 65468 32206 65506
rect 32154 65434 32163 65468
rect 32197 65434 32206 65468
rect 32154 65396 32206 65434
rect 32154 65362 32163 65396
rect 32197 65362 32206 65396
rect 32154 65334 32206 65362
rect 32240 65612 32292 65640
rect 32240 65578 32249 65612
rect 32283 65578 32292 65612
rect 32240 65540 32292 65578
rect 32240 65506 32249 65540
rect 32283 65506 32292 65540
rect 32240 65468 32292 65506
rect 32240 65456 32249 65468
rect 32283 65456 32292 65468
rect 32240 65396 32292 65404
rect 32240 65392 32249 65396
rect 32283 65392 32292 65396
rect 32240 65334 32292 65340
rect 32348 65612 32406 65640
rect 32348 65578 32360 65612
rect 32394 65578 32406 65612
rect 32348 65540 32406 65578
rect 32348 65506 32360 65540
rect 32394 65506 32406 65540
rect 32348 65468 32406 65506
rect 32348 65434 32360 65468
rect 32394 65434 32406 65468
rect 32348 65396 32406 65434
rect 32348 65362 32360 65396
rect 32394 65362 32406 65396
rect 32348 65334 32406 65362
rect 31966 65160 32000 65334
rect 32079 65284 32281 65296
rect 32079 65250 32091 65284
rect 32125 65250 32163 65284
rect 32197 65250 32235 65284
rect 32269 65250 32281 65284
rect 32079 65230 32281 65250
rect 32079 65170 32093 65230
rect 32267 65170 32281 65230
rect 23160 65100 23200 65160
rect 22760 62270 23200 65100
rect 31960 65100 32000 65160
rect 32360 65160 32394 65334
rect 32504 65246 32514 65678
rect 32584 65246 32594 65678
rect 40966 65246 40976 65678
rect 41046 65246 41056 65678
rect 41154 65612 41212 65640
rect 41154 65578 41166 65612
rect 41200 65578 41212 65612
rect 41154 65540 41212 65578
rect 41154 65506 41166 65540
rect 41200 65506 41212 65540
rect 41154 65468 41212 65506
rect 41154 65434 41166 65468
rect 41200 65434 41212 65468
rect 41154 65396 41212 65434
rect 41154 65362 41166 65396
rect 41200 65362 41212 65396
rect 41154 65334 41212 65362
rect 41268 65612 41320 65640
rect 41268 65578 41277 65612
rect 41311 65578 41320 65612
rect 41268 65540 41320 65578
rect 41268 65506 41277 65540
rect 41311 65506 41320 65540
rect 41268 65468 41320 65506
rect 41268 65456 41277 65468
rect 41311 65456 41320 65468
rect 41268 65396 41320 65404
rect 41268 65392 41277 65396
rect 41311 65392 41320 65396
rect 41268 65334 41320 65340
rect 41354 65634 41406 65640
rect 41354 65578 41363 65582
rect 41397 65578 41406 65582
rect 41354 65570 41406 65578
rect 41354 65506 41363 65518
rect 41397 65506 41406 65518
rect 41354 65468 41406 65506
rect 41354 65434 41363 65468
rect 41397 65434 41406 65468
rect 41354 65396 41406 65434
rect 41354 65362 41363 65396
rect 41397 65362 41406 65396
rect 41354 65334 41406 65362
rect 41440 65612 41492 65640
rect 41440 65578 41449 65612
rect 41483 65578 41492 65612
rect 41440 65540 41492 65578
rect 41440 65506 41449 65540
rect 41483 65506 41492 65540
rect 41440 65468 41492 65506
rect 41440 65456 41449 65468
rect 41483 65456 41492 65468
rect 41440 65396 41492 65404
rect 41440 65392 41449 65396
rect 41483 65392 41492 65396
rect 41440 65334 41492 65340
rect 41548 65612 41606 65640
rect 41548 65578 41560 65612
rect 41594 65578 41606 65612
rect 41548 65540 41606 65578
rect 41548 65506 41560 65540
rect 41594 65506 41606 65540
rect 41548 65468 41606 65506
rect 41548 65434 41560 65468
rect 41594 65434 41606 65468
rect 41548 65396 41606 65434
rect 41548 65362 41560 65396
rect 41594 65362 41606 65396
rect 41548 65334 41606 65362
rect 41166 65160 41200 65334
rect 41279 65284 41481 65296
rect 41279 65250 41291 65284
rect 41325 65250 41363 65284
rect 41397 65250 41435 65284
rect 41469 65250 41481 65284
rect 41279 65230 41481 65250
rect 41279 65170 41293 65230
rect 41467 65170 41481 65230
rect 32360 65100 32400 65160
rect 31960 62270 32400 65100
rect 41160 65100 41200 65160
rect 41560 65160 41594 65334
rect 41704 65246 41714 65678
rect 41784 65246 41794 65678
rect 50166 65246 50176 65678
rect 50246 65246 50256 65678
rect 50354 65612 50412 65640
rect 50354 65578 50366 65612
rect 50400 65578 50412 65612
rect 50354 65540 50412 65578
rect 50354 65506 50366 65540
rect 50400 65506 50412 65540
rect 50354 65468 50412 65506
rect 50354 65434 50366 65468
rect 50400 65434 50412 65468
rect 50354 65396 50412 65434
rect 50354 65362 50366 65396
rect 50400 65362 50412 65396
rect 50354 65334 50412 65362
rect 50468 65612 50520 65640
rect 50468 65578 50477 65612
rect 50511 65578 50520 65612
rect 50468 65540 50520 65578
rect 50468 65506 50477 65540
rect 50511 65506 50520 65540
rect 50468 65468 50520 65506
rect 50468 65456 50477 65468
rect 50511 65456 50520 65468
rect 50468 65396 50520 65404
rect 50468 65392 50477 65396
rect 50511 65392 50520 65396
rect 50468 65334 50520 65340
rect 50554 65634 50606 65640
rect 50554 65578 50563 65582
rect 50597 65578 50606 65582
rect 50554 65570 50606 65578
rect 50554 65506 50563 65518
rect 50597 65506 50606 65518
rect 50554 65468 50606 65506
rect 50554 65434 50563 65468
rect 50597 65434 50606 65468
rect 50554 65396 50606 65434
rect 50554 65362 50563 65396
rect 50597 65362 50606 65396
rect 50554 65334 50606 65362
rect 50640 65612 50692 65640
rect 50640 65578 50649 65612
rect 50683 65578 50692 65612
rect 50640 65540 50692 65578
rect 50640 65506 50649 65540
rect 50683 65506 50692 65540
rect 50640 65468 50692 65506
rect 50640 65456 50649 65468
rect 50683 65456 50692 65468
rect 50640 65396 50692 65404
rect 50640 65392 50649 65396
rect 50683 65392 50692 65396
rect 50640 65334 50692 65340
rect 50748 65612 50806 65640
rect 50748 65578 50760 65612
rect 50794 65578 50806 65612
rect 50748 65540 50806 65578
rect 50748 65506 50760 65540
rect 50794 65506 50806 65540
rect 50748 65468 50806 65506
rect 50748 65434 50760 65468
rect 50794 65434 50806 65468
rect 50748 65396 50806 65434
rect 50748 65362 50760 65396
rect 50794 65362 50806 65396
rect 50748 65334 50806 65362
rect 50366 65160 50400 65334
rect 50479 65284 50681 65296
rect 50479 65250 50491 65284
rect 50525 65250 50563 65284
rect 50597 65250 50635 65284
rect 50669 65250 50681 65284
rect 50479 65230 50681 65250
rect 50479 65170 50493 65230
rect 50667 65170 50681 65230
rect 41560 65100 41600 65160
rect 41160 62270 41600 65100
rect 50360 65100 50400 65160
rect 50760 65160 50794 65334
rect 50904 65246 50914 65678
rect 50984 65246 50994 65678
rect 59366 65246 59376 65678
rect 59446 65246 59456 65678
rect 59554 65612 59612 65640
rect 59554 65578 59566 65612
rect 59600 65578 59612 65612
rect 59554 65540 59612 65578
rect 59554 65506 59566 65540
rect 59600 65506 59612 65540
rect 59554 65468 59612 65506
rect 59554 65434 59566 65468
rect 59600 65434 59612 65468
rect 59554 65396 59612 65434
rect 59554 65362 59566 65396
rect 59600 65362 59612 65396
rect 59554 65334 59612 65362
rect 59668 65612 59720 65640
rect 59668 65578 59677 65612
rect 59711 65578 59720 65612
rect 59668 65540 59720 65578
rect 59668 65506 59677 65540
rect 59711 65506 59720 65540
rect 59668 65468 59720 65506
rect 59668 65456 59677 65468
rect 59711 65456 59720 65468
rect 59668 65396 59720 65404
rect 59668 65392 59677 65396
rect 59711 65392 59720 65396
rect 59668 65334 59720 65340
rect 59754 65634 59806 65640
rect 59754 65578 59763 65582
rect 59797 65578 59806 65582
rect 59754 65570 59806 65578
rect 59754 65506 59763 65518
rect 59797 65506 59806 65518
rect 59754 65468 59806 65506
rect 59754 65434 59763 65468
rect 59797 65434 59806 65468
rect 59754 65396 59806 65434
rect 59754 65362 59763 65396
rect 59797 65362 59806 65396
rect 59754 65334 59806 65362
rect 59840 65612 59892 65640
rect 59840 65578 59849 65612
rect 59883 65578 59892 65612
rect 59840 65540 59892 65578
rect 59840 65506 59849 65540
rect 59883 65506 59892 65540
rect 59840 65468 59892 65506
rect 59840 65456 59849 65468
rect 59883 65456 59892 65468
rect 59840 65396 59892 65404
rect 59840 65392 59849 65396
rect 59883 65392 59892 65396
rect 59840 65334 59892 65340
rect 59948 65612 60006 65640
rect 59948 65578 59960 65612
rect 59994 65578 60006 65612
rect 59948 65540 60006 65578
rect 59948 65506 59960 65540
rect 59994 65506 60006 65540
rect 59948 65468 60006 65506
rect 59948 65434 59960 65468
rect 59994 65434 60006 65468
rect 59948 65396 60006 65434
rect 59948 65362 59960 65396
rect 59994 65362 60006 65396
rect 59948 65334 60006 65362
rect 59566 65160 59600 65334
rect 59679 65284 59881 65296
rect 59679 65250 59691 65284
rect 59725 65250 59763 65284
rect 59797 65250 59835 65284
rect 59869 65250 59881 65284
rect 59679 65230 59881 65250
rect 59679 65170 59693 65230
rect 59867 65170 59881 65230
rect 50760 65100 50800 65160
rect 50360 62270 50800 65100
rect 59560 65100 59600 65160
rect 59960 65160 59994 65334
rect 60104 65246 60114 65678
rect 60184 65246 60194 65678
rect 68566 65246 68576 65678
rect 68646 65246 68656 65678
rect 68754 65612 68812 65640
rect 68754 65578 68766 65612
rect 68800 65578 68812 65612
rect 68754 65540 68812 65578
rect 68754 65506 68766 65540
rect 68800 65506 68812 65540
rect 68754 65468 68812 65506
rect 68754 65434 68766 65468
rect 68800 65434 68812 65468
rect 68754 65396 68812 65434
rect 68754 65362 68766 65396
rect 68800 65362 68812 65396
rect 68754 65334 68812 65362
rect 68868 65612 68920 65640
rect 68868 65578 68877 65612
rect 68911 65578 68920 65612
rect 68868 65540 68920 65578
rect 68868 65506 68877 65540
rect 68911 65506 68920 65540
rect 68868 65468 68920 65506
rect 68868 65456 68877 65468
rect 68911 65456 68920 65468
rect 68868 65396 68920 65404
rect 68868 65392 68877 65396
rect 68911 65392 68920 65396
rect 68868 65334 68920 65340
rect 68954 65634 69006 65640
rect 68954 65578 68963 65582
rect 68997 65578 69006 65582
rect 68954 65570 69006 65578
rect 68954 65506 68963 65518
rect 68997 65506 69006 65518
rect 68954 65468 69006 65506
rect 68954 65434 68963 65468
rect 68997 65434 69006 65468
rect 68954 65396 69006 65434
rect 68954 65362 68963 65396
rect 68997 65362 69006 65396
rect 68954 65334 69006 65362
rect 69040 65612 69092 65640
rect 69040 65578 69049 65612
rect 69083 65578 69092 65612
rect 69040 65540 69092 65578
rect 69040 65506 69049 65540
rect 69083 65506 69092 65540
rect 69040 65468 69092 65506
rect 69040 65456 69049 65468
rect 69083 65456 69092 65468
rect 69040 65396 69092 65404
rect 69040 65392 69049 65396
rect 69083 65392 69092 65396
rect 69040 65334 69092 65340
rect 69148 65612 69206 65640
rect 69148 65578 69160 65612
rect 69194 65578 69206 65612
rect 69148 65540 69206 65578
rect 69148 65506 69160 65540
rect 69194 65506 69206 65540
rect 69148 65468 69206 65506
rect 69148 65434 69160 65468
rect 69194 65434 69206 65468
rect 69148 65396 69206 65434
rect 69148 65362 69160 65396
rect 69194 65362 69206 65396
rect 69148 65334 69206 65362
rect 68766 65160 68800 65334
rect 68879 65284 69081 65296
rect 68879 65250 68891 65284
rect 68925 65250 68963 65284
rect 68997 65250 69035 65284
rect 69069 65250 69081 65284
rect 68879 65230 69081 65250
rect 68879 65170 68893 65230
rect 69067 65170 69081 65230
rect 59960 65100 60000 65160
rect 59560 62270 60000 65100
rect 68760 65100 68800 65160
rect 69160 65160 69194 65334
rect 69304 65246 69314 65678
rect 69384 65246 69394 65678
rect 69160 65100 69200 65160
rect 68760 62270 69200 65100
rect -3880 60270 73600 62270
rect -3880 52390 -1870 60270
rect 0 56412 77600 58270
rect 0 56270 4192 56412
rect 4186 56015 4192 56270
rect 4230 56270 4930 56412
rect 4230 56015 4236 56270
rect 4186 56003 4236 56015
rect 4924 56015 4930 56270
rect 4968 56270 13392 56412
rect 4968 56015 4974 56270
rect 4924 56003 4974 56015
rect 13386 56015 13392 56270
rect 13430 56270 14130 56412
rect 13430 56015 13436 56270
rect 13386 56003 13436 56015
rect 14124 56015 14130 56270
rect 14168 56270 22592 56412
rect 14168 56015 14174 56270
rect 14124 56003 14174 56015
rect 22586 56015 22592 56270
rect 22630 56270 23330 56412
rect 22630 56015 22636 56270
rect 22586 56003 22636 56015
rect 23324 56015 23330 56270
rect 23368 56270 31792 56412
rect 23368 56015 23374 56270
rect 23324 56003 23374 56015
rect 31786 56015 31792 56270
rect 31830 56270 32530 56412
rect 31830 56015 31836 56270
rect 31786 56003 31836 56015
rect 32524 56015 32530 56270
rect 32568 56270 40992 56412
rect 32568 56015 32574 56270
rect 32524 56003 32574 56015
rect 40986 56015 40992 56270
rect 41030 56270 41730 56412
rect 41030 56015 41036 56270
rect 40986 56003 41036 56015
rect 41724 56015 41730 56270
rect 41768 56270 50192 56412
rect 41768 56015 41774 56270
rect 41724 56003 41774 56015
rect 50186 56015 50192 56270
rect 50230 56270 50930 56412
rect 50230 56015 50236 56270
rect 50186 56003 50236 56015
rect 50924 56015 50930 56270
rect 50968 56270 59392 56412
rect 50968 56015 50974 56270
rect 50924 56003 50974 56015
rect 59386 56015 59392 56270
rect 59430 56270 60130 56412
rect 59430 56015 59436 56270
rect 59386 56003 59436 56015
rect 60124 56015 60130 56270
rect 60168 56270 68592 56412
rect 60168 56015 60174 56270
rect 60124 56003 60174 56015
rect 68586 56015 68592 56270
rect 68630 56270 69330 56412
rect 68630 56015 68636 56270
rect 68586 56003 68636 56015
rect 69324 56015 69330 56270
rect 69368 56270 77600 56412
rect 69368 56015 69374 56270
rect 69324 56003 69374 56015
rect 4479 55844 4681 55864
rect 4479 55810 4491 55844
rect 4525 55810 4563 55844
rect 4597 55810 4635 55844
rect 4669 55810 4681 55844
rect 4479 55798 4681 55810
rect 13679 55844 13881 55864
rect 13679 55810 13691 55844
rect 13725 55810 13763 55844
rect 13797 55810 13835 55844
rect 13869 55810 13881 55844
rect 13679 55798 13881 55810
rect 22879 55844 23081 55864
rect 22879 55810 22891 55844
rect 22925 55810 22963 55844
rect 22997 55810 23035 55844
rect 23069 55810 23081 55844
rect 22879 55798 23081 55810
rect 32079 55844 32281 55864
rect 32079 55810 32091 55844
rect 32125 55810 32163 55844
rect 32197 55810 32235 55844
rect 32269 55810 32281 55844
rect 32079 55798 32281 55810
rect 41279 55844 41481 55864
rect 41279 55810 41291 55844
rect 41325 55810 41363 55844
rect 41397 55810 41435 55844
rect 41469 55810 41481 55844
rect 41279 55798 41481 55810
rect 50479 55844 50681 55864
rect 50479 55810 50491 55844
rect 50525 55810 50563 55844
rect 50597 55810 50635 55844
rect 50669 55810 50681 55844
rect 50479 55798 50681 55810
rect 59679 55844 59881 55864
rect 59679 55810 59691 55844
rect 59725 55810 59763 55844
rect 59797 55810 59835 55844
rect 59869 55810 59881 55844
rect 59679 55798 59881 55810
rect 68879 55844 69081 55864
rect 68879 55810 68891 55844
rect 68925 55810 68963 55844
rect 68997 55810 69035 55844
rect 69069 55810 69081 55844
rect 68879 55798 69081 55810
rect 4166 55366 4176 55798
rect 4246 55366 4256 55798
rect 4354 55732 4412 55760
rect 4354 55698 4366 55732
rect 4400 55698 4412 55732
rect 4354 55660 4412 55698
rect 4354 55626 4366 55660
rect 4400 55626 4412 55660
rect 4354 55588 4412 55626
rect 4354 55554 4366 55588
rect 4400 55554 4412 55588
rect 4354 55516 4412 55554
rect 4354 55482 4366 55516
rect 4400 55482 4412 55516
rect 4354 55454 4412 55482
rect 4468 55732 4520 55760
rect 4468 55698 4477 55732
rect 4511 55698 4520 55732
rect 4468 55660 4520 55698
rect 4468 55626 4477 55660
rect 4511 55626 4520 55660
rect 4468 55588 4520 55626
rect 4468 55576 4477 55588
rect 4511 55576 4520 55588
rect 4468 55516 4520 55524
rect 4468 55512 4477 55516
rect 4511 55512 4520 55516
rect 4468 55454 4520 55460
rect 4554 55754 4606 55760
rect 4554 55698 4563 55702
rect 4597 55698 4606 55702
rect 4554 55690 4606 55698
rect 4554 55626 4563 55638
rect 4597 55626 4606 55638
rect 4554 55588 4606 55626
rect 4554 55554 4563 55588
rect 4597 55554 4606 55588
rect 4554 55516 4606 55554
rect 4554 55482 4563 55516
rect 4597 55482 4606 55516
rect 4554 55454 4606 55482
rect 4640 55732 4692 55760
rect 4640 55698 4649 55732
rect 4683 55698 4692 55732
rect 4640 55660 4692 55698
rect 4640 55626 4649 55660
rect 4683 55626 4692 55660
rect 4640 55588 4692 55626
rect 4640 55576 4649 55588
rect 4683 55576 4692 55588
rect 4640 55516 4692 55524
rect 4640 55512 4649 55516
rect 4683 55512 4692 55516
rect 4640 55454 4692 55460
rect 4748 55732 4806 55760
rect 4748 55698 4760 55732
rect 4794 55698 4806 55732
rect 4748 55660 4806 55698
rect 4748 55626 4760 55660
rect 4794 55626 4806 55660
rect 4748 55588 4806 55626
rect 4748 55554 4760 55588
rect 4794 55554 4806 55588
rect 4748 55516 4806 55554
rect 4748 55482 4760 55516
rect 4794 55482 4806 55516
rect 4748 55454 4806 55482
rect 4366 55280 4400 55454
rect 4479 55404 4681 55416
rect 4479 55370 4491 55404
rect 4525 55370 4563 55404
rect 4597 55370 4635 55404
rect 4669 55370 4681 55404
rect 4479 55350 4681 55370
rect 4479 55290 4493 55350
rect 4667 55290 4681 55350
rect 4360 55220 4400 55280
rect 4760 55280 4794 55454
rect 4904 55366 4914 55798
rect 4984 55366 4994 55798
rect 13366 55366 13376 55798
rect 13446 55366 13456 55798
rect 13554 55732 13612 55760
rect 13554 55698 13566 55732
rect 13600 55698 13612 55732
rect 13554 55660 13612 55698
rect 13554 55626 13566 55660
rect 13600 55626 13612 55660
rect 13554 55588 13612 55626
rect 13554 55554 13566 55588
rect 13600 55554 13612 55588
rect 13554 55516 13612 55554
rect 13554 55482 13566 55516
rect 13600 55482 13612 55516
rect 13554 55454 13612 55482
rect 13668 55732 13720 55760
rect 13668 55698 13677 55732
rect 13711 55698 13720 55732
rect 13668 55660 13720 55698
rect 13668 55626 13677 55660
rect 13711 55626 13720 55660
rect 13668 55588 13720 55626
rect 13668 55576 13677 55588
rect 13711 55576 13720 55588
rect 13668 55516 13720 55524
rect 13668 55512 13677 55516
rect 13711 55512 13720 55516
rect 13668 55454 13720 55460
rect 13754 55754 13806 55760
rect 13754 55698 13763 55702
rect 13797 55698 13806 55702
rect 13754 55690 13806 55698
rect 13754 55626 13763 55638
rect 13797 55626 13806 55638
rect 13754 55588 13806 55626
rect 13754 55554 13763 55588
rect 13797 55554 13806 55588
rect 13754 55516 13806 55554
rect 13754 55482 13763 55516
rect 13797 55482 13806 55516
rect 13754 55454 13806 55482
rect 13840 55732 13892 55760
rect 13840 55698 13849 55732
rect 13883 55698 13892 55732
rect 13840 55660 13892 55698
rect 13840 55626 13849 55660
rect 13883 55626 13892 55660
rect 13840 55588 13892 55626
rect 13840 55576 13849 55588
rect 13883 55576 13892 55588
rect 13840 55516 13892 55524
rect 13840 55512 13849 55516
rect 13883 55512 13892 55516
rect 13840 55454 13892 55460
rect 13948 55732 14006 55760
rect 13948 55698 13960 55732
rect 13994 55698 14006 55732
rect 13948 55660 14006 55698
rect 13948 55626 13960 55660
rect 13994 55626 14006 55660
rect 13948 55588 14006 55626
rect 13948 55554 13960 55588
rect 13994 55554 14006 55588
rect 13948 55516 14006 55554
rect 13948 55482 13960 55516
rect 13994 55482 14006 55516
rect 13948 55454 14006 55482
rect 13566 55280 13600 55454
rect 13679 55404 13881 55416
rect 13679 55370 13691 55404
rect 13725 55370 13763 55404
rect 13797 55370 13835 55404
rect 13869 55370 13881 55404
rect 13679 55350 13881 55370
rect 13679 55290 13693 55350
rect 13867 55290 13881 55350
rect 4760 55220 4800 55280
rect 4360 52390 4800 55220
rect 13560 55220 13600 55280
rect 13960 55280 13994 55454
rect 14104 55366 14114 55798
rect 14184 55366 14194 55798
rect 22566 55366 22576 55798
rect 22646 55366 22656 55798
rect 22754 55732 22812 55760
rect 22754 55698 22766 55732
rect 22800 55698 22812 55732
rect 22754 55660 22812 55698
rect 22754 55626 22766 55660
rect 22800 55626 22812 55660
rect 22754 55588 22812 55626
rect 22754 55554 22766 55588
rect 22800 55554 22812 55588
rect 22754 55516 22812 55554
rect 22754 55482 22766 55516
rect 22800 55482 22812 55516
rect 22754 55454 22812 55482
rect 22868 55732 22920 55760
rect 22868 55698 22877 55732
rect 22911 55698 22920 55732
rect 22868 55660 22920 55698
rect 22868 55626 22877 55660
rect 22911 55626 22920 55660
rect 22868 55588 22920 55626
rect 22868 55576 22877 55588
rect 22911 55576 22920 55588
rect 22868 55516 22920 55524
rect 22868 55512 22877 55516
rect 22911 55512 22920 55516
rect 22868 55454 22920 55460
rect 22954 55754 23006 55760
rect 22954 55698 22963 55702
rect 22997 55698 23006 55702
rect 22954 55690 23006 55698
rect 22954 55626 22963 55638
rect 22997 55626 23006 55638
rect 22954 55588 23006 55626
rect 22954 55554 22963 55588
rect 22997 55554 23006 55588
rect 22954 55516 23006 55554
rect 22954 55482 22963 55516
rect 22997 55482 23006 55516
rect 22954 55454 23006 55482
rect 23040 55732 23092 55760
rect 23040 55698 23049 55732
rect 23083 55698 23092 55732
rect 23040 55660 23092 55698
rect 23040 55626 23049 55660
rect 23083 55626 23092 55660
rect 23040 55588 23092 55626
rect 23040 55576 23049 55588
rect 23083 55576 23092 55588
rect 23040 55516 23092 55524
rect 23040 55512 23049 55516
rect 23083 55512 23092 55516
rect 23040 55454 23092 55460
rect 23148 55732 23206 55760
rect 23148 55698 23160 55732
rect 23194 55698 23206 55732
rect 23148 55660 23206 55698
rect 23148 55626 23160 55660
rect 23194 55626 23206 55660
rect 23148 55588 23206 55626
rect 23148 55554 23160 55588
rect 23194 55554 23206 55588
rect 23148 55516 23206 55554
rect 23148 55482 23160 55516
rect 23194 55482 23206 55516
rect 23148 55454 23206 55482
rect 22766 55280 22800 55454
rect 22879 55404 23081 55416
rect 22879 55370 22891 55404
rect 22925 55370 22963 55404
rect 22997 55370 23035 55404
rect 23069 55370 23081 55404
rect 22879 55350 23081 55370
rect 22879 55290 22893 55350
rect 23067 55290 23081 55350
rect 13960 55220 14000 55280
rect 13560 52390 14000 55220
rect 22760 55220 22800 55280
rect 23160 55280 23194 55454
rect 23304 55366 23314 55798
rect 23384 55366 23394 55798
rect 31766 55366 31776 55798
rect 31846 55366 31856 55798
rect 31954 55732 32012 55760
rect 31954 55698 31966 55732
rect 32000 55698 32012 55732
rect 31954 55660 32012 55698
rect 31954 55626 31966 55660
rect 32000 55626 32012 55660
rect 31954 55588 32012 55626
rect 31954 55554 31966 55588
rect 32000 55554 32012 55588
rect 31954 55516 32012 55554
rect 31954 55482 31966 55516
rect 32000 55482 32012 55516
rect 31954 55454 32012 55482
rect 32068 55732 32120 55760
rect 32068 55698 32077 55732
rect 32111 55698 32120 55732
rect 32068 55660 32120 55698
rect 32068 55626 32077 55660
rect 32111 55626 32120 55660
rect 32068 55588 32120 55626
rect 32068 55576 32077 55588
rect 32111 55576 32120 55588
rect 32068 55516 32120 55524
rect 32068 55512 32077 55516
rect 32111 55512 32120 55516
rect 32068 55454 32120 55460
rect 32154 55754 32206 55760
rect 32154 55698 32163 55702
rect 32197 55698 32206 55702
rect 32154 55690 32206 55698
rect 32154 55626 32163 55638
rect 32197 55626 32206 55638
rect 32154 55588 32206 55626
rect 32154 55554 32163 55588
rect 32197 55554 32206 55588
rect 32154 55516 32206 55554
rect 32154 55482 32163 55516
rect 32197 55482 32206 55516
rect 32154 55454 32206 55482
rect 32240 55732 32292 55760
rect 32240 55698 32249 55732
rect 32283 55698 32292 55732
rect 32240 55660 32292 55698
rect 32240 55626 32249 55660
rect 32283 55626 32292 55660
rect 32240 55588 32292 55626
rect 32240 55576 32249 55588
rect 32283 55576 32292 55588
rect 32240 55516 32292 55524
rect 32240 55512 32249 55516
rect 32283 55512 32292 55516
rect 32240 55454 32292 55460
rect 32348 55732 32406 55760
rect 32348 55698 32360 55732
rect 32394 55698 32406 55732
rect 32348 55660 32406 55698
rect 32348 55626 32360 55660
rect 32394 55626 32406 55660
rect 32348 55588 32406 55626
rect 32348 55554 32360 55588
rect 32394 55554 32406 55588
rect 32348 55516 32406 55554
rect 32348 55482 32360 55516
rect 32394 55482 32406 55516
rect 32348 55454 32406 55482
rect 31966 55280 32000 55454
rect 32079 55404 32281 55416
rect 32079 55370 32091 55404
rect 32125 55370 32163 55404
rect 32197 55370 32235 55404
rect 32269 55370 32281 55404
rect 32079 55350 32281 55370
rect 32079 55290 32093 55350
rect 32267 55290 32281 55350
rect 23160 55220 23200 55280
rect 22760 52390 23200 55220
rect 31960 55220 32000 55280
rect 32360 55280 32394 55454
rect 32504 55366 32514 55798
rect 32584 55366 32594 55798
rect 40966 55366 40976 55798
rect 41046 55366 41056 55798
rect 41154 55732 41212 55760
rect 41154 55698 41166 55732
rect 41200 55698 41212 55732
rect 41154 55660 41212 55698
rect 41154 55626 41166 55660
rect 41200 55626 41212 55660
rect 41154 55588 41212 55626
rect 41154 55554 41166 55588
rect 41200 55554 41212 55588
rect 41154 55516 41212 55554
rect 41154 55482 41166 55516
rect 41200 55482 41212 55516
rect 41154 55454 41212 55482
rect 41268 55732 41320 55760
rect 41268 55698 41277 55732
rect 41311 55698 41320 55732
rect 41268 55660 41320 55698
rect 41268 55626 41277 55660
rect 41311 55626 41320 55660
rect 41268 55588 41320 55626
rect 41268 55576 41277 55588
rect 41311 55576 41320 55588
rect 41268 55516 41320 55524
rect 41268 55512 41277 55516
rect 41311 55512 41320 55516
rect 41268 55454 41320 55460
rect 41354 55754 41406 55760
rect 41354 55698 41363 55702
rect 41397 55698 41406 55702
rect 41354 55690 41406 55698
rect 41354 55626 41363 55638
rect 41397 55626 41406 55638
rect 41354 55588 41406 55626
rect 41354 55554 41363 55588
rect 41397 55554 41406 55588
rect 41354 55516 41406 55554
rect 41354 55482 41363 55516
rect 41397 55482 41406 55516
rect 41354 55454 41406 55482
rect 41440 55732 41492 55760
rect 41440 55698 41449 55732
rect 41483 55698 41492 55732
rect 41440 55660 41492 55698
rect 41440 55626 41449 55660
rect 41483 55626 41492 55660
rect 41440 55588 41492 55626
rect 41440 55576 41449 55588
rect 41483 55576 41492 55588
rect 41440 55516 41492 55524
rect 41440 55512 41449 55516
rect 41483 55512 41492 55516
rect 41440 55454 41492 55460
rect 41548 55732 41606 55760
rect 41548 55698 41560 55732
rect 41594 55698 41606 55732
rect 41548 55660 41606 55698
rect 41548 55626 41560 55660
rect 41594 55626 41606 55660
rect 41548 55588 41606 55626
rect 41548 55554 41560 55588
rect 41594 55554 41606 55588
rect 41548 55516 41606 55554
rect 41548 55482 41560 55516
rect 41594 55482 41606 55516
rect 41548 55454 41606 55482
rect 41166 55280 41200 55454
rect 41279 55404 41481 55416
rect 41279 55370 41291 55404
rect 41325 55370 41363 55404
rect 41397 55370 41435 55404
rect 41469 55370 41481 55404
rect 41279 55350 41481 55370
rect 41279 55290 41293 55350
rect 41467 55290 41481 55350
rect 32360 55220 32400 55280
rect 31960 52390 32400 55220
rect 41160 55220 41200 55280
rect 41560 55280 41594 55454
rect 41704 55366 41714 55798
rect 41784 55366 41794 55798
rect 50166 55366 50176 55798
rect 50246 55366 50256 55798
rect 50354 55732 50412 55760
rect 50354 55698 50366 55732
rect 50400 55698 50412 55732
rect 50354 55660 50412 55698
rect 50354 55626 50366 55660
rect 50400 55626 50412 55660
rect 50354 55588 50412 55626
rect 50354 55554 50366 55588
rect 50400 55554 50412 55588
rect 50354 55516 50412 55554
rect 50354 55482 50366 55516
rect 50400 55482 50412 55516
rect 50354 55454 50412 55482
rect 50468 55732 50520 55760
rect 50468 55698 50477 55732
rect 50511 55698 50520 55732
rect 50468 55660 50520 55698
rect 50468 55626 50477 55660
rect 50511 55626 50520 55660
rect 50468 55588 50520 55626
rect 50468 55576 50477 55588
rect 50511 55576 50520 55588
rect 50468 55516 50520 55524
rect 50468 55512 50477 55516
rect 50511 55512 50520 55516
rect 50468 55454 50520 55460
rect 50554 55754 50606 55760
rect 50554 55698 50563 55702
rect 50597 55698 50606 55702
rect 50554 55690 50606 55698
rect 50554 55626 50563 55638
rect 50597 55626 50606 55638
rect 50554 55588 50606 55626
rect 50554 55554 50563 55588
rect 50597 55554 50606 55588
rect 50554 55516 50606 55554
rect 50554 55482 50563 55516
rect 50597 55482 50606 55516
rect 50554 55454 50606 55482
rect 50640 55732 50692 55760
rect 50640 55698 50649 55732
rect 50683 55698 50692 55732
rect 50640 55660 50692 55698
rect 50640 55626 50649 55660
rect 50683 55626 50692 55660
rect 50640 55588 50692 55626
rect 50640 55576 50649 55588
rect 50683 55576 50692 55588
rect 50640 55516 50692 55524
rect 50640 55512 50649 55516
rect 50683 55512 50692 55516
rect 50640 55454 50692 55460
rect 50748 55732 50806 55760
rect 50748 55698 50760 55732
rect 50794 55698 50806 55732
rect 50748 55660 50806 55698
rect 50748 55626 50760 55660
rect 50794 55626 50806 55660
rect 50748 55588 50806 55626
rect 50748 55554 50760 55588
rect 50794 55554 50806 55588
rect 50748 55516 50806 55554
rect 50748 55482 50760 55516
rect 50794 55482 50806 55516
rect 50748 55454 50806 55482
rect 50366 55280 50400 55454
rect 50479 55404 50681 55416
rect 50479 55370 50491 55404
rect 50525 55370 50563 55404
rect 50597 55370 50635 55404
rect 50669 55370 50681 55404
rect 50479 55350 50681 55370
rect 50479 55290 50493 55350
rect 50667 55290 50681 55350
rect 41560 55220 41600 55280
rect 41160 52390 41600 55220
rect 50360 55220 50400 55280
rect 50760 55280 50794 55454
rect 50904 55366 50914 55798
rect 50984 55366 50994 55798
rect 59366 55366 59376 55798
rect 59446 55366 59456 55798
rect 59554 55732 59612 55760
rect 59554 55698 59566 55732
rect 59600 55698 59612 55732
rect 59554 55660 59612 55698
rect 59554 55626 59566 55660
rect 59600 55626 59612 55660
rect 59554 55588 59612 55626
rect 59554 55554 59566 55588
rect 59600 55554 59612 55588
rect 59554 55516 59612 55554
rect 59554 55482 59566 55516
rect 59600 55482 59612 55516
rect 59554 55454 59612 55482
rect 59668 55732 59720 55760
rect 59668 55698 59677 55732
rect 59711 55698 59720 55732
rect 59668 55660 59720 55698
rect 59668 55626 59677 55660
rect 59711 55626 59720 55660
rect 59668 55588 59720 55626
rect 59668 55576 59677 55588
rect 59711 55576 59720 55588
rect 59668 55516 59720 55524
rect 59668 55512 59677 55516
rect 59711 55512 59720 55516
rect 59668 55454 59720 55460
rect 59754 55754 59806 55760
rect 59754 55698 59763 55702
rect 59797 55698 59806 55702
rect 59754 55690 59806 55698
rect 59754 55626 59763 55638
rect 59797 55626 59806 55638
rect 59754 55588 59806 55626
rect 59754 55554 59763 55588
rect 59797 55554 59806 55588
rect 59754 55516 59806 55554
rect 59754 55482 59763 55516
rect 59797 55482 59806 55516
rect 59754 55454 59806 55482
rect 59840 55732 59892 55760
rect 59840 55698 59849 55732
rect 59883 55698 59892 55732
rect 59840 55660 59892 55698
rect 59840 55626 59849 55660
rect 59883 55626 59892 55660
rect 59840 55588 59892 55626
rect 59840 55576 59849 55588
rect 59883 55576 59892 55588
rect 59840 55516 59892 55524
rect 59840 55512 59849 55516
rect 59883 55512 59892 55516
rect 59840 55454 59892 55460
rect 59948 55732 60006 55760
rect 59948 55698 59960 55732
rect 59994 55698 60006 55732
rect 59948 55660 60006 55698
rect 59948 55626 59960 55660
rect 59994 55626 60006 55660
rect 59948 55588 60006 55626
rect 59948 55554 59960 55588
rect 59994 55554 60006 55588
rect 59948 55516 60006 55554
rect 59948 55482 59960 55516
rect 59994 55482 60006 55516
rect 59948 55454 60006 55482
rect 59566 55280 59600 55454
rect 59679 55404 59881 55416
rect 59679 55370 59691 55404
rect 59725 55370 59763 55404
rect 59797 55370 59835 55404
rect 59869 55370 59881 55404
rect 59679 55350 59881 55370
rect 59679 55290 59693 55350
rect 59867 55290 59881 55350
rect 50760 55220 50800 55280
rect 50360 52390 50800 55220
rect 59560 55220 59600 55280
rect 59960 55280 59994 55454
rect 60104 55366 60114 55798
rect 60184 55366 60194 55798
rect 68566 55366 68576 55798
rect 68646 55366 68656 55798
rect 68754 55732 68812 55760
rect 68754 55698 68766 55732
rect 68800 55698 68812 55732
rect 68754 55660 68812 55698
rect 68754 55626 68766 55660
rect 68800 55626 68812 55660
rect 68754 55588 68812 55626
rect 68754 55554 68766 55588
rect 68800 55554 68812 55588
rect 68754 55516 68812 55554
rect 68754 55482 68766 55516
rect 68800 55482 68812 55516
rect 68754 55454 68812 55482
rect 68868 55732 68920 55760
rect 68868 55698 68877 55732
rect 68911 55698 68920 55732
rect 68868 55660 68920 55698
rect 68868 55626 68877 55660
rect 68911 55626 68920 55660
rect 68868 55588 68920 55626
rect 68868 55576 68877 55588
rect 68911 55576 68920 55588
rect 68868 55516 68920 55524
rect 68868 55512 68877 55516
rect 68911 55512 68920 55516
rect 68868 55454 68920 55460
rect 68954 55754 69006 55760
rect 68954 55698 68963 55702
rect 68997 55698 69006 55702
rect 68954 55690 69006 55698
rect 68954 55626 68963 55638
rect 68997 55626 69006 55638
rect 68954 55588 69006 55626
rect 68954 55554 68963 55588
rect 68997 55554 69006 55588
rect 68954 55516 69006 55554
rect 68954 55482 68963 55516
rect 68997 55482 69006 55516
rect 68954 55454 69006 55482
rect 69040 55732 69092 55760
rect 69040 55698 69049 55732
rect 69083 55698 69092 55732
rect 69040 55660 69092 55698
rect 69040 55626 69049 55660
rect 69083 55626 69092 55660
rect 69040 55588 69092 55626
rect 69040 55576 69049 55588
rect 69083 55576 69092 55588
rect 69040 55516 69092 55524
rect 69040 55512 69049 55516
rect 69083 55512 69092 55516
rect 69040 55454 69092 55460
rect 69148 55732 69206 55760
rect 69148 55698 69160 55732
rect 69194 55698 69206 55732
rect 69148 55660 69206 55698
rect 69148 55626 69160 55660
rect 69194 55626 69206 55660
rect 69148 55588 69206 55626
rect 69148 55554 69160 55588
rect 69194 55554 69206 55588
rect 69148 55516 69206 55554
rect 69148 55482 69160 55516
rect 69194 55482 69206 55516
rect 69148 55454 69206 55482
rect 68766 55280 68800 55454
rect 68879 55404 69081 55416
rect 68879 55370 68891 55404
rect 68925 55370 68963 55404
rect 68997 55370 69035 55404
rect 69069 55370 69081 55404
rect 68879 55350 69081 55370
rect 68879 55290 68893 55350
rect 69067 55290 69081 55350
rect 59960 55220 60000 55280
rect 59560 52390 60000 55220
rect 68760 55220 68800 55280
rect 69160 55280 69194 55454
rect 69304 55366 69314 55798
rect 69384 55366 69394 55798
rect 69160 55220 69200 55280
rect 68760 52390 69200 55220
rect -3880 50390 73600 52390
rect -3880 44900 -1870 50390
rect 75600 48390 77600 56270
rect -610 46532 77600 48390
rect -610 46390 4192 46532
rect -610 45360 -550 46390
rect -510 46140 -220 46160
rect -510 46080 -490 46140
rect -240 46080 -220 46140
rect 4186 46135 4192 46390
rect 4230 46390 4930 46532
rect 4230 46135 4236 46390
rect 4186 46123 4236 46135
rect 4924 46135 4930 46390
rect 4968 46390 13392 46532
rect 4968 46135 4974 46390
rect 4924 46123 4974 46135
rect 13386 46135 13392 46390
rect 13430 46390 14130 46532
rect 13430 46135 13436 46390
rect 13386 46123 13436 46135
rect 14124 46135 14130 46390
rect 14168 46390 22592 46532
rect 14168 46135 14174 46390
rect 14124 46123 14174 46135
rect 22586 46135 22592 46390
rect 22630 46390 23330 46532
rect 22630 46135 22636 46390
rect 22586 46123 22636 46135
rect 23324 46135 23330 46390
rect 23368 46390 31792 46532
rect 23368 46135 23374 46390
rect 23324 46123 23374 46135
rect 31786 46135 31792 46390
rect 31830 46390 32530 46532
rect 31830 46135 31836 46390
rect 31786 46123 31836 46135
rect 32524 46135 32530 46390
rect 32568 46390 40992 46532
rect 32568 46135 32574 46390
rect 32524 46123 32574 46135
rect 40986 46135 40992 46390
rect 41030 46390 41730 46532
rect 41030 46135 41036 46390
rect 40986 46123 41036 46135
rect 41724 46135 41730 46390
rect 41768 46390 50192 46532
rect 41768 46135 41774 46390
rect 41724 46123 41774 46135
rect 50186 46135 50192 46390
rect 50230 46390 50930 46532
rect 50230 46135 50236 46390
rect 50186 46123 50236 46135
rect 50924 46135 50930 46390
rect 50968 46390 59392 46532
rect 50968 46135 50974 46390
rect 50924 46123 50974 46135
rect 59386 46135 59392 46390
rect 59430 46390 60130 46532
rect 59430 46135 59436 46390
rect 59386 46123 59436 46135
rect 60124 46135 60130 46390
rect 60168 46390 68592 46532
rect 60168 46135 60174 46390
rect 60124 46123 60174 46135
rect 68586 46135 68592 46390
rect 68630 46390 69330 46532
rect 68630 46135 68636 46390
rect 68586 46123 68636 46135
rect 69324 46135 69330 46390
rect 69368 46390 77600 46532
rect 69368 46135 69374 46390
rect 69324 46123 69374 46135
rect -510 46060 -220 46080
rect -430 45984 -384 45996
rect -430 45408 -424 45984
rect -390 45408 -384 45984
rect -430 45396 -384 45408
rect -342 45984 -296 45996
rect -342 45408 -336 45984
rect -302 45408 -296 45984
rect 4479 45964 4681 45984
rect 4479 45930 4491 45964
rect 4525 45930 4563 45964
rect 4597 45930 4635 45964
rect 4669 45930 4681 45964
rect 4479 45918 4681 45930
rect 13679 45964 13881 45984
rect 13679 45930 13691 45964
rect 13725 45930 13763 45964
rect 13797 45930 13835 45964
rect 13869 45930 13881 45964
rect 13679 45918 13881 45930
rect 22879 45964 23081 45984
rect 22879 45930 22891 45964
rect 22925 45930 22963 45964
rect 22997 45930 23035 45964
rect 23069 45930 23081 45964
rect 22879 45918 23081 45930
rect 32079 45964 32281 45984
rect 32079 45930 32091 45964
rect 32125 45930 32163 45964
rect 32197 45930 32235 45964
rect 32269 45930 32281 45964
rect 32079 45918 32281 45930
rect 41279 45964 41481 45984
rect 41279 45930 41291 45964
rect 41325 45930 41363 45964
rect 41397 45930 41435 45964
rect 41469 45930 41481 45964
rect 41279 45918 41481 45930
rect 50479 45964 50681 45984
rect 50479 45930 50491 45964
rect 50525 45930 50563 45964
rect 50597 45930 50635 45964
rect 50669 45930 50681 45964
rect 50479 45918 50681 45930
rect 59679 45964 59881 45984
rect 59679 45930 59691 45964
rect 59725 45930 59763 45964
rect 59797 45930 59835 45964
rect 59869 45930 59881 45964
rect 59679 45918 59881 45930
rect 68879 45964 69081 45984
rect 68879 45930 68891 45964
rect 68925 45930 68963 45964
rect 68997 45930 69035 45964
rect 69069 45930 69081 45964
rect 68879 45918 69081 45930
rect 4166 45486 4176 45918
rect 4246 45486 4256 45918
rect 4354 45852 4412 45880
rect 4354 45818 4366 45852
rect 4400 45818 4412 45852
rect 4354 45780 4412 45818
rect 4354 45746 4366 45780
rect 4400 45746 4412 45780
rect 4354 45708 4412 45746
rect 4354 45674 4366 45708
rect 4400 45674 4412 45708
rect 4354 45636 4412 45674
rect 4354 45602 4366 45636
rect 4400 45602 4412 45636
rect 4354 45574 4412 45602
rect 4468 45852 4520 45880
rect 4468 45818 4477 45852
rect 4511 45818 4520 45852
rect 4468 45780 4520 45818
rect 4468 45746 4477 45780
rect 4511 45746 4520 45780
rect 4468 45708 4520 45746
rect 4468 45696 4477 45708
rect 4511 45696 4520 45708
rect 4468 45636 4520 45644
rect 4468 45632 4477 45636
rect 4511 45632 4520 45636
rect 4468 45574 4520 45580
rect 4554 45874 4606 45880
rect 4554 45818 4563 45822
rect 4597 45818 4606 45822
rect 4554 45810 4606 45818
rect 4554 45746 4563 45758
rect 4597 45746 4606 45758
rect 4554 45708 4606 45746
rect 4554 45674 4563 45708
rect 4597 45674 4606 45708
rect 4554 45636 4606 45674
rect 4554 45602 4563 45636
rect 4597 45602 4606 45636
rect 4554 45574 4606 45602
rect 4640 45852 4692 45880
rect 4640 45818 4649 45852
rect 4683 45818 4692 45852
rect 4640 45780 4692 45818
rect 4640 45746 4649 45780
rect 4683 45746 4692 45780
rect 4640 45708 4692 45746
rect 4640 45696 4649 45708
rect 4683 45696 4692 45708
rect 4640 45636 4692 45644
rect 4640 45632 4649 45636
rect 4683 45632 4692 45636
rect 4640 45574 4692 45580
rect 4748 45852 4806 45880
rect 4748 45818 4760 45852
rect 4794 45818 4806 45852
rect 4748 45780 4806 45818
rect 4748 45746 4760 45780
rect 4794 45746 4806 45780
rect 4748 45708 4806 45746
rect 4748 45674 4760 45708
rect 4794 45674 4806 45708
rect 4748 45636 4806 45674
rect 4748 45602 4760 45636
rect 4794 45602 4806 45636
rect 4748 45574 4806 45602
rect -342 45396 -296 45408
rect 4366 45400 4400 45574
rect 4479 45524 4681 45536
rect 4479 45490 4491 45524
rect 4525 45490 4563 45524
rect 4597 45490 4635 45524
rect 4669 45490 4681 45524
rect 4479 45470 4681 45490
rect 4479 45410 4493 45470
rect 4667 45410 4681 45470
rect -610 45320 -600 45360
rect -560 45350 -550 45360
rect -240 45350 -160 45360
rect -560 45320 -430 45350
rect -610 45310 -430 45320
rect -610 45300 -550 45310
rect -240 45290 -230 45350
rect -170 45290 -160 45350
rect -240 45280 -160 45290
rect 4360 45340 4400 45400
rect 4760 45400 4794 45574
rect 4904 45486 4914 45918
rect 4984 45486 4994 45918
rect 13366 45486 13376 45918
rect 13446 45486 13456 45918
rect 13554 45852 13612 45880
rect 13554 45818 13566 45852
rect 13600 45818 13612 45852
rect 13554 45780 13612 45818
rect 13554 45746 13566 45780
rect 13600 45746 13612 45780
rect 13554 45708 13612 45746
rect 13554 45674 13566 45708
rect 13600 45674 13612 45708
rect 13554 45636 13612 45674
rect 13554 45602 13566 45636
rect 13600 45602 13612 45636
rect 13554 45574 13612 45602
rect 13668 45852 13720 45880
rect 13668 45818 13677 45852
rect 13711 45818 13720 45852
rect 13668 45780 13720 45818
rect 13668 45746 13677 45780
rect 13711 45746 13720 45780
rect 13668 45708 13720 45746
rect 13668 45696 13677 45708
rect 13711 45696 13720 45708
rect 13668 45636 13720 45644
rect 13668 45632 13677 45636
rect 13711 45632 13720 45636
rect 13668 45574 13720 45580
rect 13754 45874 13806 45880
rect 13754 45818 13763 45822
rect 13797 45818 13806 45822
rect 13754 45810 13806 45818
rect 13754 45746 13763 45758
rect 13797 45746 13806 45758
rect 13754 45708 13806 45746
rect 13754 45674 13763 45708
rect 13797 45674 13806 45708
rect 13754 45636 13806 45674
rect 13754 45602 13763 45636
rect 13797 45602 13806 45636
rect 13754 45574 13806 45602
rect 13840 45852 13892 45880
rect 13840 45818 13849 45852
rect 13883 45818 13892 45852
rect 13840 45780 13892 45818
rect 13840 45746 13849 45780
rect 13883 45746 13892 45780
rect 13840 45708 13892 45746
rect 13840 45696 13849 45708
rect 13883 45696 13892 45708
rect 13840 45636 13892 45644
rect 13840 45632 13849 45636
rect 13883 45632 13892 45636
rect 13840 45574 13892 45580
rect 13948 45852 14006 45880
rect 13948 45818 13960 45852
rect 13994 45818 14006 45852
rect 13948 45780 14006 45818
rect 13948 45746 13960 45780
rect 13994 45746 14006 45780
rect 13948 45708 14006 45746
rect 13948 45674 13960 45708
rect 13994 45674 14006 45708
rect 13948 45636 14006 45674
rect 13948 45602 13960 45636
rect 13994 45602 14006 45636
rect 13948 45574 14006 45602
rect 13566 45400 13600 45574
rect 13679 45524 13881 45536
rect 13679 45490 13691 45524
rect 13725 45490 13763 45524
rect 13797 45490 13835 45524
rect 13869 45490 13881 45524
rect 13679 45470 13881 45490
rect 13679 45410 13693 45470
rect 13867 45410 13881 45470
rect 4760 45340 4800 45400
rect -430 45254 -384 45266
rect -430 44978 -424 45254
rect -390 44978 -384 45254
rect -430 44966 -384 44978
rect -342 45254 -296 45266
rect -342 44978 -336 45254
rect -302 44978 -296 45254
rect -342 44966 -296 44978
rect -3880 44890 0 44900
rect -3880 44840 -440 44890
rect -390 44840 -330 44890
rect -280 44840 0 44890
rect -3880 44820 0 44840
rect -3880 42510 -1870 44820
rect 4360 42510 4800 45340
rect 13560 45340 13600 45400
rect 13960 45400 13994 45574
rect 14104 45486 14114 45918
rect 14184 45486 14194 45918
rect 22566 45486 22576 45918
rect 22646 45486 22656 45918
rect 22754 45852 22812 45880
rect 22754 45818 22766 45852
rect 22800 45818 22812 45852
rect 22754 45780 22812 45818
rect 22754 45746 22766 45780
rect 22800 45746 22812 45780
rect 22754 45708 22812 45746
rect 22754 45674 22766 45708
rect 22800 45674 22812 45708
rect 22754 45636 22812 45674
rect 22754 45602 22766 45636
rect 22800 45602 22812 45636
rect 22754 45574 22812 45602
rect 22868 45852 22920 45880
rect 22868 45818 22877 45852
rect 22911 45818 22920 45852
rect 22868 45780 22920 45818
rect 22868 45746 22877 45780
rect 22911 45746 22920 45780
rect 22868 45708 22920 45746
rect 22868 45696 22877 45708
rect 22911 45696 22920 45708
rect 22868 45636 22920 45644
rect 22868 45632 22877 45636
rect 22911 45632 22920 45636
rect 22868 45574 22920 45580
rect 22954 45874 23006 45880
rect 22954 45818 22963 45822
rect 22997 45818 23006 45822
rect 22954 45810 23006 45818
rect 22954 45746 22963 45758
rect 22997 45746 23006 45758
rect 22954 45708 23006 45746
rect 22954 45674 22963 45708
rect 22997 45674 23006 45708
rect 22954 45636 23006 45674
rect 22954 45602 22963 45636
rect 22997 45602 23006 45636
rect 22954 45574 23006 45602
rect 23040 45852 23092 45880
rect 23040 45818 23049 45852
rect 23083 45818 23092 45852
rect 23040 45780 23092 45818
rect 23040 45746 23049 45780
rect 23083 45746 23092 45780
rect 23040 45708 23092 45746
rect 23040 45696 23049 45708
rect 23083 45696 23092 45708
rect 23040 45636 23092 45644
rect 23040 45632 23049 45636
rect 23083 45632 23092 45636
rect 23040 45574 23092 45580
rect 23148 45852 23206 45880
rect 23148 45818 23160 45852
rect 23194 45818 23206 45852
rect 23148 45780 23206 45818
rect 23148 45746 23160 45780
rect 23194 45746 23206 45780
rect 23148 45708 23206 45746
rect 23148 45674 23160 45708
rect 23194 45674 23206 45708
rect 23148 45636 23206 45674
rect 23148 45602 23160 45636
rect 23194 45602 23206 45636
rect 23148 45574 23206 45602
rect 22766 45400 22800 45574
rect 22879 45524 23081 45536
rect 22879 45490 22891 45524
rect 22925 45490 22963 45524
rect 22997 45490 23035 45524
rect 23069 45490 23081 45524
rect 22879 45470 23081 45490
rect 22879 45410 22893 45470
rect 23067 45410 23081 45470
rect 13960 45340 14000 45400
rect 13560 42510 14000 45340
rect 22760 45340 22800 45400
rect 23160 45400 23194 45574
rect 23304 45486 23314 45918
rect 23384 45486 23394 45918
rect 31766 45486 31776 45918
rect 31846 45486 31856 45918
rect 31954 45852 32012 45880
rect 31954 45818 31966 45852
rect 32000 45818 32012 45852
rect 31954 45780 32012 45818
rect 31954 45746 31966 45780
rect 32000 45746 32012 45780
rect 31954 45708 32012 45746
rect 31954 45674 31966 45708
rect 32000 45674 32012 45708
rect 31954 45636 32012 45674
rect 31954 45602 31966 45636
rect 32000 45602 32012 45636
rect 31954 45574 32012 45602
rect 32068 45852 32120 45880
rect 32068 45818 32077 45852
rect 32111 45818 32120 45852
rect 32068 45780 32120 45818
rect 32068 45746 32077 45780
rect 32111 45746 32120 45780
rect 32068 45708 32120 45746
rect 32068 45696 32077 45708
rect 32111 45696 32120 45708
rect 32068 45636 32120 45644
rect 32068 45632 32077 45636
rect 32111 45632 32120 45636
rect 32068 45574 32120 45580
rect 32154 45874 32206 45880
rect 32154 45818 32163 45822
rect 32197 45818 32206 45822
rect 32154 45810 32206 45818
rect 32154 45746 32163 45758
rect 32197 45746 32206 45758
rect 32154 45708 32206 45746
rect 32154 45674 32163 45708
rect 32197 45674 32206 45708
rect 32154 45636 32206 45674
rect 32154 45602 32163 45636
rect 32197 45602 32206 45636
rect 32154 45574 32206 45602
rect 32240 45852 32292 45880
rect 32240 45818 32249 45852
rect 32283 45818 32292 45852
rect 32240 45780 32292 45818
rect 32240 45746 32249 45780
rect 32283 45746 32292 45780
rect 32240 45708 32292 45746
rect 32240 45696 32249 45708
rect 32283 45696 32292 45708
rect 32240 45636 32292 45644
rect 32240 45632 32249 45636
rect 32283 45632 32292 45636
rect 32240 45574 32292 45580
rect 32348 45852 32406 45880
rect 32348 45818 32360 45852
rect 32394 45818 32406 45852
rect 32348 45780 32406 45818
rect 32348 45746 32360 45780
rect 32394 45746 32406 45780
rect 32348 45708 32406 45746
rect 32348 45674 32360 45708
rect 32394 45674 32406 45708
rect 32348 45636 32406 45674
rect 32348 45602 32360 45636
rect 32394 45602 32406 45636
rect 32348 45574 32406 45602
rect 31966 45400 32000 45574
rect 32079 45524 32281 45536
rect 32079 45490 32091 45524
rect 32125 45490 32163 45524
rect 32197 45490 32235 45524
rect 32269 45490 32281 45524
rect 32079 45470 32281 45490
rect 32079 45410 32093 45470
rect 32267 45410 32281 45470
rect 23160 45340 23200 45400
rect 22760 42510 23200 45340
rect 31960 45340 32000 45400
rect 32360 45400 32394 45574
rect 32504 45486 32514 45918
rect 32584 45486 32594 45918
rect 40966 45486 40976 45918
rect 41046 45486 41056 45918
rect 41154 45852 41212 45880
rect 41154 45818 41166 45852
rect 41200 45818 41212 45852
rect 41154 45780 41212 45818
rect 41154 45746 41166 45780
rect 41200 45746 41212 45780
rect 41154 45708 41212 45746
rect 41154 45674 41166 45708
rect 41200 45674 41212 45708
rect 41154 45636 41212 45674
rect 41154 45602 41166 45636
rect 41200 45602 41212 45636
rect 41154 45574 41212 45602
rect 41268 45852 41320 45880
rect 41268 45818 41277 45852
rect 41311 45818 41320 45852
rect 41268 45780 41320 45818
rect 41268 45746 41277 45780
rect 41311 45746 41320 45780
rect 41268 45708 41320 45746
rect 41268 45696 41277 45708
rect 41311 45696 41320 45708
rect 41268 45636 41320 45644
rect 41268 45632 41277 45636
rect 41311 45632 41320 45636
rect 41268 45574 41320 45580
rect 41354 45874 41406 45880
rect 41354 45818 41363 45822
rect 41397 45818 41406 45822
rect 41354 45810 41406 45818
rect 41354 45746 41363 45758
rect 41397 45746 41406 45758
rect 41354 45708 41406 45746
rect 41354 45674 41363 45708
rect 41397 45674 41406 45708
rect 41354 45636 41406 45674
rect 41354 45602 41363 45636
rect 41397 45602 41406 45636
rect 41354 45574 41406 45602
rect 41440 45852 41492 45880
rect 41440 45818 41449 45852
rect 41483 45818 41492 45852
rect 41440 45780 41492 45818
rect 41440 45746 41449 45780
rect 41483 45746 41492 45780
rect 41440 45708 41492 45746
rect 41440 45696 41449 45708
rect 41483 45696 41492 45708
rect 41440 45636 41492 45644
rect 41440 45632 41449 45636
rect 41483 45632 41492 45636
rect 41440 45574 41492 45580
rect 41548 45852 41606 45880
rect 41548 45818 41560 45852
rect 41594 45818 41606 45852
rect 41548 45780 41606 45818
rect 41548 45746 41560 45780
rect 41594 45746 41606 45780
rect 41548 45708 41606 45746
rect 41548 45674 41560 45708
rect 41594 45674 41606 45708
rect 41548 45636 41606 45674
rect 41548 45602 41560 45636
rect 41594 45602 41606 45636
rect 41548 45574 41606 45602
rect 41166 45400 41200 45574
rect 41279 45524 41481 45536
rect 41279 45490 41291 45524
rect 41325 45490 41363 45524
rect 41397 45490 41435 45524
rect 41469 45490 41481 45524
rect 41279 45470 41481 45490
rect 41279 45410 41293 45470
rect 41467 45410 41481 45470
rect 32360 45340 32400 45400
rect 31960 42510 32400 45340
rect 41160 45340 41200 45400
rect 41560 45400 41594 45574
rect 41704 45486 41714 45918
rect 41784 45486 41794 45918
rect 50166 45486 50176 45918
rect 50246 45486 50256 45918
rect 50354 45852 50412 45880
rect 50354 45818 50366 45852
rect 50400 45818 50412 45852
rect 50354 45780 50412 45818
rect 50354 45746 50366 45780
rect 50400 45746 50412 45780
rect 50354 45708 50412 45746
rect 50354 45674 50366 45708
rect 50400 45674 50412 45708
rect 50354 45636 50412 45674
rect 50354 45602 50366 45636
rect 50400 45602 50412 45636
rect 50354 45574 50412 45602
rect 50468 45852 50520 45880
rect 50468 45818 50477 45852
rect 50511 45818 50520 45852
rect 50468 45780 50520 45818
rect 50468 45746 50477 45780
rect 50511 45746 50520 45780
rect 50468 45708 50520 45746
rect 50468 45696 50477 45708
rect 50511 45696 50520 45708
rect 50468 45636 50520 45644
rect 50468 45632 50477 45636
rect 50511 45632 50520 45636
rect 50468 45574 50520 45580
rect 50554 45874 50606 45880
rect 50554 45818 50563 45822
rect 50597 45818 50606 45822
rect 50554 45810 50606 45818
rect 50554 45746 50563 45758
rect 50597 45746 50606 45758
rect 50554 45708 50606 45746
rect 50554 45674 50563 45708
rect 50597 45674 50606 45708
rect 50554 45636 50606 45674
rect 50554 45602 50563 45636
rect 50597 45602 50606 45636
rect 50554 45574 50606 45602
rect 50640 45852 50692 45880
rect 50640 45818 50649 45852
rect 50683 45818 50692 45852
rect 50640 45780 50692 45818
rect 50640 45746 50649 45780
rect 50683 45746 50692 45780
rect 50640 45708 50692 45746
rect 50640 45696 50649 45708
rect 50683 45696 50692 45708
rect 50640 45636 50692 45644
rect 50640 45632 50649 45636
rect 50683 45632 50692 45636
rect 50640 45574 50692 45580
rect 50748 45852 50806 45880
rect 50748 45818 50760 45852
rect 50794 45818 50806 45852
rect 50748 45780 50806 45818
rect 50748 45746 50760 45780
rect 50794 45746 50806 45780
rect 50748 45708 50806 45746
rect 50748 45674 50760 45708
rect 50794 45674 50806 45708
rect 50748 45636 50806 45674
rect 50748 45602 50760 45636
rect 50794 45602 50806 45636
rect 50748 45574 50806 45602
rect 50366 45400 50400 45574
rect 50479 45524 50681 45536
rect 50479 45490 50491 45524
rect 50525 45490 50563 45524
rect 50597 45490 50635 45524
rect 50669 45490 50681 45524
rect 50479 45470 50681 45490
rect 50479 45410 50493 45470
rect 50667 45410 50681 45470
rect 41560 45340 41600 45400
rect 41160 42510 41600 45340
rect 50360 45340 50400 45400
rect 50760 45400 50794 45574
rect 50904 45486 50914 45918
rect 50984 45486 50994 45918
rect 59366 45486 59376 45918
rect 59446 45486 59456 45918
rect 59554 45852 59612 45880
rect 59554 45818 59566 45852
rect 59600 45818 59612 45852
rect 59554 45780 59612 45818
rect 59554 45746 59566 45780
rect 59600 45746 59612 45780
rect 59554 45708 59612 45746
rect 59554 45674 59566 45708
rect 59600 45674 59612 45708
rect 59554 45636 59612 45674
rect 59554 45602 59566 45636
rect 59600 45602 59612 45636
rect 59554 45574 59612 45602
rect 59668 45852 59720 45880
rect 59668 45818 59677 45852
rect 59711 45818 59720 45852
rect 59668 45780 59720 45818
rect 59668 45746 59677 45780
rect 59711 45746 59720 45780
rect 59668 45708 59720 45746
rect 59668 45696 59677 45708
rect 59711 45696 59720 45708
rect 59668 45636 59720 45644
rect 59668 45632 59677 45636
rect 59711 45632 59720 45636
rect 59668 45574 59720 45580
rect 59754 45874 59806 45880
rect 59754 45818 59763 45822
rect 59797 45818 59806 45822
rect 59754 45810 59806 45818
rect 59754 45746 59763 45758
rect 59797 45746 59806 45758
rect 59754 45708 59806 45746
rect 59754 45674 59763 45708
rect 59797 45674 59806 45708
rect 59754 45636 59806 45674
rect 59754 45602 59763 45636
rect 59797 45602 59806 45636
rect 59754 45574 59806 45602
rect 59840 45852 59892 45880
rect 59840 45818 59849 45852
rect 59883 45818 59892 45852
rect 59840 45780 59892 45818
rect 59840 45746 59849 45780
rect 59883 45746 59892 45780
rect 59840 45708 59892 45746
rect 59840 45696 59849 45708
rect 59883 45696 59892 45708
rect 59840 45636 59892 45644
rect 59840 45632 59849 45636
rect 59883 45632 59892 45636
rect 59840 45574 59892 45580
rect 59948 45852 60006 45880
rect 59948 45818 59960 45852
rect 59994 45818 60006 45852
rect 59948 45780 60006 45818
rect 59948 45746 59960 45780
rect 59994 45746 60006 45780
rect 59948 45708 60006 45746
rect 59948 45674 59960 45708
rect 59994 45674 60006 45708
rect 59948 45636 60006 45674
rect 59948 45602 59960 45636
rect 59994 45602 60006 45636
rect 59948 45574 60006 45602
rect 59566 45400 59600 45574
rect 59679 45524 59881 45536
rect 59679 45490 59691 45524
rect 59725 45490 59763 45524
rect 59797 45490 59835 45524
rect 59869 45490 59881 45524
rect 59679 45470 59881 45490
rect 59679 45410 59693 45470
rect 59867 45410 59881 45470
rect 50760 45340 50800 45400
rect 50360 42510 50800 45340
rect 59560 45340 59600 45400
rect 59960 45400 59994 45574
rect 60104 45486 60114 45918
rect 60184 45486 60194 45918
rect 68566 45486 68576 45918
rect 68646 45486 68656 45918
rect 68754 45852 68812 45880
rect 68754 45818 68766 45852
rect 68800 45818 68812 45852
rect 68754 45780 68812 45818
rect 68754 45746 68766 45780
rect 68800 45746 68812 45780
rect 68754 45708 68812 45746
rect 68754 45674 68766 45708
rect 68800 45674 68812 45708
rect 68754 45636 68812 45674
rect 68754 45602 68766 45636
rect 68800 45602 68812 45636
rect 68754 45574 68812 45602
rect 68868 45852 68920 45880
rect 68868 45818 68877 45852
rect 68911 45818 68920 45852
rect 68868 45780 68920 45818
rect 68868 45746 68877 45780
rect 68911 45746 68920 45780
rect 68868 45708 68920 45746
rect 68868 45696 68877 45708
rect 68911 45696 68920 45708
rect 68868 45636 68920 45644
rect 68868 45632 68877 45636
rect 68911 45632 68920 45636
rect 68868 45574 68920 45580
rect 68954 45874 69006 45880
rect 68954 45818 68963 45822
rect 68997 45818 69006 45822
rect 68954 45810 69006 45818
rect 68954 45746 68963 45758
rect 68997 45746 69006 45758
rect 68954 45708 69006 45746
rect 68954 45674 68963 45708
rect 68997 45674 69006 45708
rect 68954 45636 69006 45674
rect 68954 45602 68963 45636
rect 68997 45602 69006 45636
rect 68954 45574 69006 45602
rect 69040 45852 69092 45880
rect 69040 45818 69049 45852
rect 69083 45818 69092 45852
rect 69040 45780 69092 45818
rect 69040 45746 69049 45780
rect 69083 45746 69092 45780
rect 69040 45708 69092 45746
rect 69040 45696 69049 45708
rect 69083 45696 69092 45708
rect 69040 45636 69092 45644
rect 69040 45632 69049 45636
rect 69083 45632 69092 45636
rect 69040 45574 69092 45580
rect 69148 45852 69206 45880
rect 69148 45818 69160 45852
rect 69194 45818 69206 45852
rect 69148 45780 69206 45818
rect 69148 45746 69160 45780
rect 69194 45746 69206 45780
rect 69148 45708 69206 45746
rect 69148 45674 69160 45708
rect 69194 45674 69206 45708
rect 69148 45636 69206 45674
rect 69148 45602 69160 45636
rect 69194 45602 69206 45636
rect 69148 45574 69206 45602
rect 68766 45400 68800 45574
rect 68879 45524 69081 45536
rect 68879 45490 68891 45524
rect 68925 45490 68963 45524
rect 68997 45490 69035 45524
rect 69069 45490 69081 45524
rect 68879 45470 69081 45490
rect 68879 45410 68893 45470
rect 69067 45410 69081 45470
rect 59960 45340 60000 45400
rect 59560 42510 60000 45340
rect 68760 45340 68800 45400
rect 69160 45400 69194 45574
rect 69304 45486 69314 45918
rect 69384 45486 69394 45918
rect 69160 45340 69200 45400
rect 68760 42510 69200 45340
rect -3880 40510 73600 42510
rect -3880 32630 -1870 40510
rect 0 36652 77600 38510
rect 0 36510 4192 36652
rect 4186 36255 4192 36510
rect 4230 36510 4930 36652
rect 4230 36255 4236 36510
rect 4186 36243 4236 36255
rect 4924 36255 4930 36510
rect 4968 36510 13392 36652
rect 4968 36255 4974 36510
rect 4924 36243 4974 36255
rect 13386 36255 13392 36510
rect 13430 36510 14130 36652
rect 13430 36255 13436 36510
rect 13386 36243 13436 36255
rect 14124 36255 14130 36510
rect 14168 36510 22592 36652
rect 14168 36255 14174 36510
rect 14124 36243 14174 36255
rect 22586 36255 22592 36510
rect 22630 36510 23330 36652
rect 22630 36255 22636 36510
rect 22586 36243 22636 36255
rect 23324 36255 23330 36510
rect 23368 36510 31792 36652
rect 23368 36255 23374 36510
rect 23324 36243 23374 36255
rect 31786 36255 31792 36510
rect 31830 36510 32530 36652
rect 31830 36255 31836 36510
rect 31786 36243 31836 36255
rect 32524 36255 32530 36510
rect 32568 36510 40992 36652
rect 32568 36255 32574 36510
rect 32524 36243 32574 36255
rect 40986 36255 40992 36510
rect 41030 36510 41730 36652
rect 41030 36255 41036 36510
rect 40986 36243 41036 36255
rect 41724 36255 41730 36510
rect 41768 36510 50192 36652
rect 41768 36255 41774 36510
rect 41724 36243 41774 36255
rect 50186 36255 50192 36510
rect 50230 36510 50930 36652
rect 50230 36255 50236 36510
rect 50186 36243 50236 36255
rect 50924 36255 50930 36510
rect 50968 36510 59392 36652
rect 50968 36255 50974 36510
rect 50924 36243 50974 36255
rect 59386 36255 59392 36510
rect 59430 36510 60130 36652
rect 59430 36255 59436 36510
rect 59386 36243 59436 36255
rect 60124 36255 60130 36510
rect 60168 36510 68592 36652
rect 60168 36255 60174 36510
rect 60124 36243 60174 36255
rect 68586 36255 68592 36510
rect 68630 36510 69330 36652
rect 68630 36255 68636 36510
rect 68586 36243 68636 36255
rect 69324 36255 69330 36510
rect 69368 36510 77600 36652
rect 69368 36255 69374 36510
rect 69324 36243 69374 36255
rect 4479 36084 4681 36104
rect 4479 36050 4491 36084
rect 4525 36050 4563 36084
rect 4597 36050 4635 36084
rect 4669 36050 4681 36084
rect 4479 36038 4681 36050
rect 13679 36084 13881 36104
rect 13679 36050 13691 36084
rect 13725 36050 13763 36084
rect 13797 36050 13835 36084
rect 13869 36050 13881 36084
rect 13679 36038 13881 36050
rect 22879 36084 23081 36104
rect 22879 36050 22891 36084
rect 22925 36050 22963 36084
rect 22997 36050 23035 36084
rect 23069 36050 23081 36084
rect 22879 36038 23081 36050
rect 32079 36084 32281 36104
rect 32079 36050 32091 36084
rect 32125 36050 32163 36084
rect 32197 36050 32235 36084
rect 32269 36050 32281 36084
rect 32079 36038 32281 36050
rect 41279 36084 41481 36104
rect 41279 36050 41291 36084
rect 41325 36050 41363 36084
rect 41397 36050 41435 36084
rect 41469 36050 41481 36084
rect 41279 36038 41481 36050
rect 50479 36084 50681 36104
rect 50479 36050 50491 36084
rect 50525 36050 50563 36084
rect 50597 36050 50635 36084
rect 50669 36050 50681 36084
rect 50479 36038 50681 36050
rect 59679 36084 59881 36104
rect 59679 36050 59691 36084
rect 59725 36050 59763 36084
rect 59797 36050 59835 36084
rect 59869 36050 59881 36084
rect 59679 36038 59881 36050
rect 68879 36084 69081 36104
rect 68879 36050 68891 36084
rect 68925 36050 68963 36084
rect 68997 36050 69035 36084
rect 69069 36050 69081 36084
rect 68879 36038 69081 36050
rect 4166 35606 4176 36038
rect 4246 35606 4256 36038
rect 4354 35972 4412 36000
rect 4354 35938 4366 35972
rect 4400 35938 4412 35972
rect 4354 35900 4412 35938
rect 4354 35866 4366 35900
rect 4400 35866 4412 35900
rect 4354 35828 4412 35866
rect 4354 35794 4366 35828
rect 4400 35794 4412 35828
rect 4354 35756 4412 35794
rect 4354 35722 4366 35756
rect 4400 35722 4412 35756
rect 4354 35694 4412 35722
rect 4468 35972 4520 36000
rect 4468 35938 4477 35972
rect 4511 35938 4520 35972
rect 4468 35900 4520 35938
rect 4468 35866 4477 35900
rect 4511 35866 4520 35900
rect 4468 35828 4520 35866
rect 4468 35816 4477 35828
rect 4511 35816 4520 35828
rect 4468 35756 4520 35764
rect 4468 35752 4477 35756
rect 4511 35752 4520 35756
rect 4468 35694 4520 35700
rect 4554 35994 4606 36000
rect 4554 35938 4563 35942
rect 4597 35938 4606 35942
rect 4554 35930 4606 35938
rect 4554 35866 4563 35878
rect 4597 35866 4606 35878
rect 4554 35828 4606 35866
rect 4554 35794 4563 35828
rect 4597 35794 4606 35828
rect 4554 35756 4606 35794
rect 4554 35722 4563 35756
rect 4597 35722 4606 35756
rect 4554 35694 4606 35722
rect 4640 35972 4692 36000
rect 4640 35938 4649 35972
rect 4683 35938 4692 35972
rect 4640 35900 4692 35938
rect 4640 35866 4649 35900
rect 4683 35866 4692 35900
rect 4640 35828 4692 35866
rect 4640 35816 4649 35828
rect 4683 35816 4692 35828
rect 4640 35756 4692 35764
rect 4640 35752 4649 35756
rect 4683 35752 4692 35756
rect 4640 35694 4692 35700
rect 4748 35972 4806 36000
rect 4748 35938 4760 35972
rect 4794 35938 4806 35972
rect 4748 35900 4806 35938
rect 4748 35866 4760 35900
rect 4794 35866 4806 35900
rect 4748 35828 4806 35866
rect 4748 35794 4760 35828
rect 4794 35794 4806 35828
rect 4748 35756 4806 35794
rect 4748 35722 4760 35756
rect 4794 35722 4806 35756
rect 4748 35694 4806 35722
rect 4366 35520 4400 35694
rect 4479 35644 4681 35656
rect 4479 35610 4491 35644
rect 4525 35610 4563 35644
rect 4597 35610 4635 35644
rect 4669 35610 4681 35644
rect 4479 35590 4681 35610
rect 4479 35530 4493 35590
rect 4667 35530 4681 35590
rect 4360 35460 4400 35520
rect 4760 35520 4794 35694
rect 4904 35606 4914 36038
rect 4984 35606 4994 36038
rect 13366 35606 13376 36038
rect 13446 35606 13456 36038
rect 13554 35972 13612 36000
rect 13554 35938 13566 35972
rect 13600 35938 13612 35972
rect 13554 35900 13612 35938
rect 13554 35866 13566 35900
rect 13600 35866 13612 35900
rect 13554 35828 13612 35866
rect 13554 35794 13566 35828
rect 13600 35794 13612 35828
rect 13554 35756 13612 35794
rect 13554 35722 13566 35756
rect 13600 35722 13612 35756
rect 13554 35694 13612 35722
rect 13668 35972 13720 36000
rect 13668 35938 13677 35972
rect 13711 35938 13720 35972
rect 13668 35900 13720 35938
rect 13668 35866 13677 35900
rect 13711 35866 13720 35900
rect 13668 35828 13720 35866
rect 13668 35816 13677 35828
rect 13711 35816 13720 35828
rect 13668 35756 13720 35764
rect 13668 35752 13677 35756
rect 13711 35752 13720 35756
rect 13668 35694 13720 35700
rect 13754 35994 13806 36000
rect 13754 35938 13763 35942
rect 13797 35938 13806 35942
rect 13754 35930 13806 35938
rect 13754 35866 13763 35878
rect 13797 35866 13806 35878
rect 13754 35828 13806 35866
rect 13754 35794 13763 35828
rect 13797 35794 13806 35828
rect 13754 35756 13806 35794
rect 13754 35722 13763 35756
rect 13797 35722 13806 35756
rect 13754 35694 13806 35722
rect 13840 35972 13892 36000
rect 13840 35938 13849 35972
rect 13883 35938 13892 35972
rect 13840 35900 13892 35938
rect 13840 35866 13849 35900
rect 13883 35866 13892 35900
rect 13840 35828 13892 35866
rect 13840 35816 13849 35828
rect 13883 35816 13892 35828
rect 13840 35756 13892 35764
rect 13840 35752 13849 35756
rect 13883 35752 13892 35756
rect 13840 35694 13892 35700
rect 13948 35972 14006 36000
rect 13948 35938 13960 35972
rect 13994 35938 14006 35972
rect 13948 35900 14006 35938
rect 13948 35866 13960 35900
rect 13994 35866 14006 35900
rect 13948 35828 14006 35866
rect 13948 35794 13960 35828
rect 13994 35794 14006 35828
rect 13948 35756 14006 35794
rect 13948 35722 13960 35756
rect 13994 35722 14006 35756
rect 13948 35694 14006 35722
rect 13566 35520 13600 35694
rect 13679 35644 13881 35656
rect 13679 35610 13691 35644
rect 13725 35610 13763 35644
rect 13797 35610 13835 35644
rect 13869 35610 13881 35644
rect 13679 35590 13881 35610
rect 13679 35530 13693 35590
rect 13867 35530 13881 35590
rect 4760 35460 4800 35520
rect 4360 32630 4800 35460
rect 13560 35460 13600 35520
rect 13960 35520 13994 35694
rect 14104 35606 14114 36038
rect 14184 35606 14194 36038
rect 22566 35606 22576 36038
rect 22646 35606 22656 36038
rect 22754 35972 22812 36000
rect 22754 35938 22766 35972
rect 22800 35938 22812 35972
rect 22754 35900 22812 35938
rect 22754 35866 22766 35900
rect 22800 35866 22812 35900
rect 22754 35828 22812 35866
rect 22754 35794 22766 35828
rect 22800 35794 22812 35828
rect 22754 35756 22812 35794
rect 22754 35722 22766 35756
rect 22800 35722 22812 35756
rect 22754 35694 22812 35722
rect 22868 35972 22920 36000
rect 22868 35938 22877 35972
rect 22911 35938 22920 35972
rect 22868 35900 22920 35938
rect 22868 35866 22877 35900
rect 22911 35866 22920 35900
rect 22868 35828 22920 35866
rect 22868 35816 22877 35828
rect 22911 35816 22920 35828
rect 22868 35756 22920 35764
rect 22868 35752 22877 35756
rect 22911 35752 22920 35756
rect 22868 35694 22920 35700
rect 22954 35994 23006 36000
rect 22954 35938 22963 35942
rect 22997 35938 23006 35942
rect 22954 35930 23006 35938
rect 22954 35866 22963 35878
rect 22997 35866 23006 35878
rect 22954 35828 23006 35866
rect 22954 35794 22963 35828
rect 22997 35794 23006 35828
rect 22954 35756 23006 35794
rect 22954 35722 22963 35756
rect 22997 35722 23006 35756
rect 22954 35694 23006 35722
rect 23040 35972 23092 36000
rect 23040 35938 23049 35972
rect 23083 35938 23092 35972
rect 23040 35900 23092 35938
rect 23040 35866 23049 35900
rect 23083 35866 23092 35900
rect 23040 35828 23092 35866
rect 23040 35816 23049 35828
rect 23083 35816 23092 35828
rect 23040 35756 23092 35764
rect 23040 35752 23049 35756
rect 23083 35752 23092 35756
rect 23040 35694 23092 35700
rect 23148 35972 23206 36000
rect 23148 35938 23160 35972
rect 23194 35938 23206 35972
rect 23148 35900 23206 35938
rect 23148 35866 23160 35900
rect 23194 35866 23206 35900
rect 23148 35828 23206 35866
rect 23148 35794 23160 35828
rect 23194 35794 23206 35828
rect 23148 35756 23206 35794
rect 23148 35722 23160 35756
rect 23194 35722 23206 35756
rect 23148 35694 23206 35722
rect 22766 35520 22800 35694
rect 22879 35644 23081 35656
rect 22879 35610 22891 35644
rect 22925 35610 22963 35644
rect 22997 35610 23035 35644
rect 23069 35610 23081 35644
rect 22879 35590 23081 35610
rect 22879 35530 22893 35590
rect 23067 35530 23081 35590
rect 13960 35460 14000 35520
rect 13560 32630 14000 35460
rect 22760 35460 22800 35520
rect 23160 35520 23194 35694
rect 23304 35606 23314 36038
rect 23384 35606 23394 36038
rect 31766 35606 31776 36038
rect 31846 35606 31856 36038
rect 31954 35972 32012 36000
rect 31954 35938 31966 35972
rect 32000 35938 32012 35972
rect 31954 35900 32012 35938
rect 31954 35866 31966 35900
rect 32000 35866 32012 35900
rect 31954 35828 32012 35866
rect 31954 35794 31966 35828
rect 32000 35794 32012 35828
rect 31954 35756 32012 35794
rect 31954 35722 31966 35756
rect 32000 35722 32012 35756
rect 31954 35694 32012 35722
rect 32068 35972 32120 36000
rect 32068 35938 32077 35972
rect 32111 35938 32120 35972
rect 32068 35900 32120 35938
rect 32068 35866 32077 35900
rect 32111 35866 32120 35900
rect 32068 35828 32120 35866
rect 32068 35816 32077 35828
rect 32111 35816 32120 35828
rect 32068 35756 32120 35764
rect 32068 35752 32077 35756
rect 32111 35752 32120 35756
rect 32068 35694 32120 35700
rect 32154 35994 32206 36000
rect 32154 35938 32163 35942
rect 32197 35938 32206 35942
rect 32154 35930 32206 35938
rect 32154 35866 32163 35878
rect 32197 35866 32206 35878
rect 32154 35828 32206 35866
rect 32154 35794 32163 35828
rect 32197 35794 32206 35828
rect 32154 35756 32206 35794
rect 32154 35722 32163 35756
rect 32197 35722 32206 35756
rect 32154 35694 32206 35722
rect 32240 35972 32292 36000
rect 32240 35938 32249 35972
rect 32283 35938 32292 35972
rect 32240 35900 32292 35938
rect 32240 35866 32249 35900
rect 32283 35866 32292 35900
rect 32240 35828 32292 35866
rect 32240 35816 32249 35828
rect 32283 35816 32292 35828
rect 32240 35756 32292 35764
rect 32240 35752 32249 35756
rect 32283 35752 32292 35756
rect 32240 35694 32292 35700
rect 32348 35972 32406 36000
rect 32348 35938 32360 35972
rect 32394 35938 32406 35972
rect 32348 35900 32406 35938
rect 32348 35866 32360 35900
rect 32394 35866 32406 35900
rect 32348 35828 32406 35866
rect 32348 35794 32360 35828
rect 32394 35794 32406 35828
rect 32348 35756 32406 35794
rect 32348 35722 32360 35756
rect 32394 35722 32406 35756
rect 32348 35694 32406 35722
rect 31966 35520 32000 35694
rect 32079 35644 32281 35656
rect 32079 35610 32091 35644
rect 32125 35610 32163 35644
rect 32197 35610 32235 35644
rect 32269 35610 32281 35644
rect 32079 35590 32281 35610
rect 32079 35530 32093 35590
rect 32267 35530 32281 35590
rect 23160 35460 23200 35520
rect 22760 32630 23200 35460
rect 31960 35460 32000 35520
rect 32360 35520 32394 35694
rect 32504 35606 32514 36038
rect 32584 35606 32594 36038
rect 40966 35606 40976 36038
rect 41046 35606 41056 36038
rect 41154 35972 41212 36000
rect 41154 35938 41166 35972
rect 41200 35938 41212 35972
rect 41154 35900 41212 35938
rect 41154 35866 41166 35900
rect 41200 35866 41212 35900
rect 41154 35828 41212 35866
rect 41154 35794 41166 35828
rect 41200 35794 41212 35828
rect 41154 35756 41212 35794
rect 41154 35722 41166 35756
rect 41200 35722 41212 35756
rect 41154 35694 41212 35722
rect 41268 35972 41320 36000
rect 41268 35938 41277 35972
rect 41311 35938 41320 35972
rect 41268 35900 41320 35938
rect 41268 35866 41277 35900
rect 41311 35866 41320 35900
rect 41268 35828 41320 35866
rect 41268 35816 41277 35828
rect 41311 35816 41320 35828
rect 41268 35756 41320 35764
rect 41268 35752 41277 35756
rect 41311 35752 41320 35756
rect 41268 35694 41320 35700
rect 41354 35994 41406 36000
rect 41354 35938 41363 35942
rect 41397 35938 41406 35942
rect 41354 35930 41406 35938
rect 41354 35866 41363 35878
rect 41397 35866 41406 35878
rect 41354 35828 41406 35866
rect 41354 35794 41363 35828
rect 41397 35794 41406 35828
rect 41354 35756 41406 35794
rect 41354 35722 41363 35756
rect 41397 35722 41406 35756
rect 41354 35694 41406 35722
rect 41440 35972 41492 36000
rect 41440 35938 41449 35972
rect 41483 35938 41492 35972
rect 41440 35900 41492 35938
rect 41440 35866 41449 35900
rect 41483 35866 41492 35900
rect 41440 35828 41492 35866
rect 41440 35816 41449 35828
rect 41483 35816 41492 35828
rect 41440 35756 41492 35764
rect 41440 35752 41449 35756
rect 41483 35752 41492 35756
rect 41440 35694 41492 35700
rect 41548 35972 41606 36000
rect 41548 35938 41560 35972
rect 41594 35938 41606 35972
rect 41548 35900 41606 35938
rect 41548 35866 41560 35900
rect 41594 35866 41606 35900
rect 41548 35828 41606 35866
rect 41548 35794 41560 35828
rect 41594 35794 41606 35828
rect 41548 35756 41606 35794
rect 41548 35722 41560 35756
rect 41594 35722 41606 35756
rect 41548 35694 41606 35722
rect 41166 35520 41200 35694
rect 41279 35644 41481 35656
rect 41279 35610 41291 35644
rect 41325 35610 41363 35644
rect 41397 35610 41435 35644
rect 41469 35610 41481 35644
rect 41279 35590 41481 35610
rect 41279 35530 41293 35590
rect 41467 35530 41481 35590
rect 32360 35460 32400 35520
rect 31960 32630 32400 35460
rect 41160 35460 41200 35520
rect 41560 35520 41594 35694
rect 41704 35606 41714 36038
rect 41784 35606 41794 36038
rect 50166 35606 50176 36038
rect 50246 35606 50256 36038
rect 50354 35972 50412 36000
rect 50354 35938 50366 35972
rect 50400 35938 50412 35972
rect 50354 35900 50412 35938
rect 50354 35866 50366 35900
rect 50400 35866 50412 35900
rect 50354 35828 50412 35866
rect 50354 35794 50366 35828
rect 50400 35794 50412 35828
rect 50354 35756 50412 35794
rect 50354 35722 50366 35756
rect 50400 35722 50412 35756
rect 50354 35694 50412 35722
rect 50468 35972 50520 36000
rect 50468 35938 50477 35972
rect 50511 35938 50520 35972
rect 50468 35900 50520 35938
rect 50468 35866 50477 35900
rect 50511 35866 50520 35900
rect 50468 35828 50520 35866
rect 50468 35816 50477 35828
rect 50511 35816 50520 35828
rect 50468 35756 50520 35764
rect 50468 35752 50477 35756
rect 50511 35752 50520 35756
rect 50468 35694 50520 35700
rect 50554 35994 50606 36000
rect 50554 35938 50563 35942
rect 50597 35938 50606 35942
rect 50554 35930 50606 35938
rect 50554 35866 50563 35878
rect 50597 35866 50606 35878
rect 50554 35828 50606 35866
rect 50554 35794 50563 35828
rect 50597 35794 50606 35828
rect 50554 35756 50606 35794
rect 50554 35722 50563 35756
rect 50597 35722 50606 35756
rect 50554 35694 50606 35722
rect 50640 35972 50692 36000
rect 50640 35938 50649 35972
rect 50683 35938 50692 35972
rect 50640 35900 50692 35938
rect 50640 35866 50649 35900
rect 50683 35866 50692 35900
rect 50640 35828 50692 35866
rect 50640 35816 50649 35828
rect 50683 35816 50692 35828
rect 50640 35756 50692 35764
rect 50640 35752 50649 35756
rect 50683 35752 50692 35756
rect 50640 35694 50692 35700
rect 50748 35972 50806 36000
rect 50748 35938 50760 35972
rect 50794 35938 50806 35972
rect 50748 35900 50806 35938
rect 50748 35866 50760 35900
rect 50794 35866 50806 35900
rect 50748 35828 50806 35866
rect 50748 35794 50760 35828
rect 50794 35794 50806 35828
rect 50748 35756 50806 35794
rect 50748 35722 50760 35756
rect 50794 35722 50806 35756
rect 50748 35694 50806 35722
rect 50366 35520 50400 35694
rect 50479 35644 50681 35656
rect 50479 35610 50491 35644
rect 50525 35610 50563 35644
rect 50597 35610 50635 35644
rect 50669 35610 50681 35644
rect 50479 35590 50681 35610
rect 50479 35530 50493 35590
rect 50667 35530 50681 35590
rect 41560 35460 41600 35520
rect 41160 32630 41600 35460
rect 50360 35460 50400 35520
rect 50760 35520 50794 35694
rect 50904 35606 50914 36038
rect 50984 35606 50994 36038
rect 59366 35606 59376 36038
rect 59446 35606 59456 36038
rect 59554 35972 59612 36000
rect 59554 35938 59566 35972
rect 59600 35938 59612 35972
rect 59554 35900 59612 35938
rect 59554 35866 59566 35900
rect 59600 35866 59612 35900
rect 59554 35828 59612 35866
rect 59554 35794 59566 35828
rect 59600 35794 59612 35828
rect 59554 35756 59612 35794
rect 59554 35722 59566 35756
rect 59600 35722 59612 35756
rect 59554 35694 59612 35722
rect 59668 35972 59720 36000
rect 59668 35938 59677 35972
rect 59711 35938 59720 35972
rect 59668 35900 59720 35938
rect 59668 35866 59677 35900
rect 59711 35866 59720 35900
rect 59668 35828 59720 35866
rect 59668 35816 59677 35828
rect 59711 35816 59720 35828
rect 59668 35756 59720 35764
rect 59668 35752 59677 35756
rect 59711 35752 59720 35756
rect 59668 35694 59720 35700
rect 59754 35994 59806 36000
rect 59754 35938 59763 35942
rect 59797 35938 59806 35942
rect 59754 35930 59806 35938
rect 59754 35866 59763 35878
rect 59797 35866 59806 35878
rect 59754 35828 59806 35866
rect 59754 35794 59763 35828
rect 59797 35794 59806 35828
rect 59754 35756 59806 35794
rect 59754 35722 59763 35756
rect 59797 35722 59806 35756
rect 59754 35694 59806 35722
rect 59840 35972 59892 36000
rect 59840 35938 59849 35972
rect 59883 35938 59892 35972
rect 59840 35900 59892 35938
rect 59840 35866 59849 35900
rect 59883 35866 59892 35900
rect 59840 35828 59892 35866
rect 59840 35816 59849 35828
rect 59883 35816 59892 35828
rect 59840 35756 59892 35764
rect 59840 35752 59849 35756
rect 59883 35752 59892 35756
rect 59840 35694 59892 35700
rect 59948 35972 60006 36000
rect 59948 35938 59960 35972
rect 59994 35938 60006 35972
rect 59948 35900 60006 35938
rect 59948 35866 59960 35900
rect 59994 35866 60006 35900
rect 59948 35828 60006 35866
rect 59948 35794 59960 35828
rect 59994 35794 60006 35828
rect 59948 35756 60006 35794
rect 59948 35722 59960 35756
rect 59994 35722 60006 35756
rect 59948 35694 60006 35722
rect 59566 35520 59600 35694
rect 59679 35644 59881 35656
rect 59679 35610 59691 35644
rect 59725 35610 59763 35644
rect 59797 35610 59835 35644
rect 59869 35610 59881 35644
rect 59679 35590 59881 35610
rect 59679 35530 59693 35590
rect 59867 35530 59881 35590
rect 50760 35460 50800 35520
rect 50360 32630 50800 35460
rect 59560 35460 59600 35520
rect 59960 35520 59994 35694
rect 60104 35606 60114 36038
rect 60184 35606 60194 36038
rect 68566 35606 68576 36038
rect 68646 35606 68656 36038
rect 68754 35972 68812 36000
rect 68754 35938 68766 35972
rect 68800 35938 68812 35972
rect 68754 35900 68812 35938
rect 68754 35866 68766 35900
rect 68800 35866 68812 35900
rect 68754 35828 68812 35866
rect 68754 35794 68766 35828
rect 68800 35794 68812 35828
rect 68754 35756 68812 35794
rect 68754 35722 68766 35756
rect 68800 35722 68812 35756
rect 68754 35694 68812 35722
rect 68868 35972 68920 36000
rect 68868 35938 68877 35972
rect 68911 35938 68920 35972
rect 68868 35900 68920 35938
rect 68868 35866 68877 35900
rect 68911 35866 68920 35900
rect 68868 35828 68920 35866
rect 68868 35816 68877 35828
rect 68911 35816 68920 35828
rect 68868 35756 68920 35764
rect 68868 35752 68877 35756
rect 68911 35752 68920 35756
rect 68868 35694 68920 35700
rect 68954 35994 69006 36000
rect 68954 35938 68963 35942
rect 68997 35938 69006 35942
rect 68954 35930 69006 35938
rect 68954 35866 68963 35878
rect 68997 35866 69006 35878
rect 68954 35828 69006 35866
rect 68954 35794 68963 35828
rect 68997 35794 69006 35828
rect 68954 35756 69006 35794
rect 68954 35722 68963 35756
rect 68997 35722 69006 35756
rect 68954 35694 69006 35722
rect 69040 35972 69092 36000
rect 69040 35938 69049 35972
rect 69083 35938 69092 35972
rect 69040 35900 69092 35938
rect 69040 35866 69049 35900
rect 69083 35866 69092 35900
rect 69040 35828 69092 35866
rect 69040 35816 69049 35828
rect 69083 35816 69092 35828
rect 69040 35756 69092 35764
rect 69040 35752 69049 35756
rect 69083 35752 69092 35756
rect 69040 35694 69092 35700
rect 69148 35972 69206 36000
rect 69148 35938 69160 35972
rect 69194 35938 69206 35972
rect 69148 35900 69206 35938
rect 69148 35866 69160 35900
rect 69194 35866 69206 35900
rect 69148 35828 69206 35866
rect 69148 35794 69160 35828
rect 69194 35794 69206 35828
rect 69148 35756 69206 35794
rect 69148 35722 69160 35756
rect 69194 35722 69206 35756
rect 69148 35694 69206 35722
rect 68766 35520 68800 35694
rect 68879 35644 69081 35656
rect 68879 35610 68891 35644
rect 68925 35610 68963 35644
rect 68997 35610 69035 35644
rect 69069 35610 69081 35644
rect 68879 35590 69081 35610
rect 68879 35530 68893 35590
rect 69067 35530 69081 35590
rect 59960 35460 60000 35520
rect 59560 32630 60000 35460
rect 68760 35460 68800 35520
rect 69160 35520 69194 35694
rect 69304 35606 69314 36038
rect 69384 35606 69394 36038
rect 69160 35460 69200 35520
rect 68760 32630 69200 35460
rect -3880 30630 73600 32630
rect -3880 22750 -1870 30630
rect 75600 28630 77600 36510
rect 0 26772 77600 28630
rect 0 26630 4192 26772
rect 4186 26375 4192 26630
rect 4230 26630 4930 26772
rect 4230 26375 4236 26630
rect 4186 26363 4236 26375
rect 4924 26375 4930 26630
rect 4968 26630 13392 26772
rect 4968 26375 4974 26630
rect 4924 26363 4974 26375
rect 13386 26375 13392 26630
rect 13430 26630 14130 26772
rect 13430 26375 13436 26630
rect 13386 26363 13436 26375
rect 14124 26375 14130 26630
rect 14168 26630 22592 26772
rect 14168 26375 14174 26630
rect 14124 26363 14174 26375
rect 22586 26375 22592 26630
rect 22630 26630 23330 26772
rect 22630 26375 22636 26630
rect 22586 26363 22636 26375
rect 23324 26375 23330 26630
rect 23368 26630 31792 26772
rect 23368 26375 23374 26630
rect 23324 26363 23374 26375
rect 31786 26375 31792 26630
rect 31830 26630 32530 26772
rect 31830 26375 31836 26630
rect 31786 26363 31836 26375
rect 32524 26375 32530 26630
rect 32568 26630 40992 26772
rect 32568 26375 32574 26630
rect 32524 26363 32574 26375
rect 40986 26375 40992 26630
rect 41030 26630 41730 26772
rect 41030 26375 41036 26630
rect 40986 26363 41036 26375
rect 41724 26375 41730 26630
rect 41768 26630 50192 26772
rect 41768 26375 41774 26630
rect 41724 26363 41774 26375
rect 50186 26375 50192 26630
rect 50230 26630 50930 26772
rect 50230 26375 50236 26630
rect 50186 26363 50236 26375
rect 50924 26375 50930 26630
rect 50968 26630 59392 26772
rect 50968 26375 50974 26630
rect 50924 26363 50974 26375
rect 59386 26375 59392 26630
rect 59430 26630 60130 26772
rect 59430 26375 59436 26630
rect 59386 26363 59436 26375
rect 60124 26375 60130 26630
rect 60168 26630 68592 26772
rect 60168 26375 60174 26630
rect 60124 26363 60174 26375
rect 68586 26375 68592 26630
rect 68630 26630 69330 26772
rect 68630 26375 68636 26630
rect 68586 26363 68636 26375
rect 69324 26375 69330 26630
rect 69368 26630 77600 26772
rect 69368 26375 69374 26630
rect 69324 26363 69374 26375
rect 4479 26204 4681 26224
rect 4479 26170 4491 26204
rect 4525 26170 4563 26204
rect 4597 26170 4635 26204
rect 4669 26170 4681 26204
rect 4479 26158 4681 26170
rect 13679 26204 13881 26224
rect 13679 26170 13691 26204
rect 13725 26170 13763 26204
rect 13797 26170 13835 26204
rect 13869 26170 13881 26204
rect 13679 26158 13881 26170
rect 22879 26204 23081 26224
rect 22879 26170 22891 26204
rect 22925 26170 22963 26204
rect 22997 26170 23035 26204
rect 23069 26170 23081 26204
rect 22879 26158 23081 26170
rect 32079 26204 32281 26224
rect 32079 26170 32091 26204
rect 32125 26170 32163 26204
rect 32197 26170 32235 26204
rect 32269 26170 32281 26204
rect 32079 26158 32281 26170
rect 41279 26204 41481 26224
rect 41279 26170 41291 26204
rect 41325 26170 41363 26204
rect 41397 26170 41435 26204
rect 41469 26170 41481 26204
rect 41279 26158 41481 26170
rect 50479 26204 50681 26224
rect 50479 26170 50491 26204
rect 50525 26170 50563 26204
rect 50597 26170 50635 26204
rect 50669 26170 50681 26204
rect 50479 26158 50681 26170
rect 59679 26204 59881 26224
rect 59679 26170 59691 26204
rect 59725 26170 59763 26204
rect 59797 26170 59835 26204
rect 59869 26170 59881 26204
rect 59679 26158 59881 26170
rect 68879 26204 69081 26224
rect 68879 26170 68891 26204
rect 68925 26170 68963 26204
rect 68997 26170 69035 26204
rect 69069 26170 69081 26204
rect 68879 26158 69081 26170
rect 4166 25726 4176 26158
rect 4246 25726 4256 26158
rect 4354 26092 4412 26120
rect 4354 26058 4366 26092
rect 4400 26058 4412 26092
rect 4354 26020 4412 26058
rect 4354 25986 4366 26020
rect 4400 25986 4412 26020
rect 4354 25948 4412 25986
rect 4354 25914 4366 25948
rect 4400 25914 4412 25948
rect 4354 25876 4412 25914
rect 4354 25842 4366 25876
rect 4400 25842 4412 25876
rect 4354 25814 4412 25842
rect 4468 26092 4520 26120
rect 4468 26058 4477 26092
rect 4511 26058 4520 26092
rect 4468 26020 4520 26058
rect 4468 25986 4477 26020
rect 4511 25986 4520 26020
rect 4468 25948 4520 25986
rect 4468 25936 4477 25948
rect 4511 25936 4520 25948
rect 4468 25876 4520 25884
rect 4468 25872 4477 25876
rect 4511 25872 4520 25876
rect 4468 25814 4520 25820
rect 4554 26114 4606 26120
rect 4554 26058 4563 26062
rect 4597 26058 4606 26062
rect 4554 26050 4606 26058
rect 4554 25986 4563 25998
rect 4597 25986 4606 25998
rect 4554 25948 4606 25986
rect 4554 25914 4563 25948
rect 4597 25914 4606 25948
rect 4554 25876 4606 25914
rect 4554 25842 4563 25876
rect 4597 25842 4606 25876
rect 4554 25814 4606 25842
rect 4640 26092 4692 26120
rect 4640 26058 4649 26092
rect 4683 26058 4692 26092
rect 4640 26020 4692 26058
rect 4640 25986 4649 26020
rect 4683 25986 4692 26020
rect 4640 25948 4692 25986
rect 4640 25936 4649 25948
rect 4683 25936 4692 25948
rect 4640 25876 4692 25884
rect 4640 25872 4649 25876
rect 4683 25872 4692 25876
rect 4640 25814 4692 25820
rect 4748 26092 4806 26120
rect 4748 26058 4760 26092
rect 4794 26058 4806 26092
rect 4748 26020 4806 26058
rect 4748 25986 4760 26020
rect 4794 25986 4806 26020
rect 4748 25948 4806 25986
rect 4748 25914 4760 25948
rect 4794 25914 4806 25948
rect 4748 25876 4806 25914
rect 4748 25842 4760 25876
rect 4794 25842 4806 25876
rect 4748 25814 4806 25842
rect 4366 25640 4400 25814
rect 4479 25764 4681 25776
rect 4479 25730 4491 25764
rect 4525 25730 4563 25764
rect 4597 25730 4635 25764
rect 4669 25730 4681 25764
rect 4479 25710 4681 25730
rect 4479 25650 4493 25710
rect 4667 25650 4681 25710
rect 4360 25580 4400 25640
rect 4760 25640 4794 25814
rect 4904 25726 4914 26158
rect 4984 25726 4994 26158
rect 13366 25726 13376 26158
rect 13446 25726 13456 26158
rect 13554 26092 13612 26120
rect 13554 26058 13566 26092
rect 13600 26058 13612 26092
rect 13554 26020 13612 26058
rect 13554 25986 13566 26020
rect 13600 25986 13612 26020
rect 13554 25948 13612 25986
rect 13554 25914 13566 25948
rect 13600 25914 13612 25948
rect 13554 25876 13612 25914
rect 13554 25842 13566 25876
rect 13600 25842 13612 25876
rect 13554 25814 13612 25842
rect 13668 26092 13720 26120
rect 13668 26058 13677 26092
rect 13711 26058 13720 26092
rect 13668 26020 13720 26058
rect 13668 25986 13677 26020
rect 13711 25986 13720 26020
rect 13668 25948 13720 25986
rect 13668 25936 13677 25948
rect 13711 25936 13720 25948
rect 13668 25876 13720 25884
rect 13668 25872 13677 25876
rect 13711 25872 13720 25876
rect 13668 25814 13720 25820
rect 13754 26114 13806 26120
rect 13754 26058 13763 26062
rect 13797 26058 13806 26062
rect 13754 26050 13806 26058
rect 13754 25986 13763 25998
rect 13797 25986 13806 25998
rect 13754 25948 13806 25986
rect 13754 25914 13763 25948
rect 13797 25914 13806 25948
rect 13754 25876 13806 25914
rect 13754 25842 13763 25876
rect 13797 25842 13806 25876
rect 13754 25814 13806 25842
rect 13840 26092 13892 26120
rect 13840 26058 13849 26092
rect 13883 26058 13892 26092
rect 13840 26020 13892 26058
rect 13840 25986 13849 26020
rect 13883 25986 13892 26020
rect 13840 25948 13892 25986
rect 13840 25936 13849 25948
rect 13883 25936 13892 25948
rect 13840 25876 13892 25884
rect 13840 25872 13849 25876
rect 13883 25872 13892 25876
rect 13840 25814 13892 25820
rect 13948 26092 14006 26120
rect 13948 26058 13960 26092
rect 13994 26058 14006 26092
rect 13948 26020 14006 26058
rect 13948 25986 13960 26020
rect 13994 25986 14006 26020
rect 13948 25948 14006 25986
rect 13948 25914 13960 25948
rect 13994 25914 14006 25948
rect 13948 25876 14006 25914
rect 13948 25842 13960 25876
rect 13994 25842 14006 25876
rect 13948 25814 14006 25842
rect 13566 25640 13600 25814
rect 13679 25764 13881 25776
rect 13679 25730 13691 25764
rect 13725 25730 13763 25764
rect 13797 25730 13835 25764
rect 13869 25730 13881 25764
rect 13679 25710 13881 25730
rect 13679 25650 13693 25710
rect 13867 25650 13881 25710
rect 4760 25580 4800 25640
rect 4360 22750 4800 25580
rect 13560 25580 13600 25640
rect 13960 25640 13994 25814
rect 14104 25726 14114 26158
rect 14184 25726 14194 26158
rect 22566 25726 22576 26158
rect 22646 25726 22656 26158
rect 22754 26092 22812 26120
rect 22754 26058 22766 26092
rect 22800 26058 22812 26092
rect 22754 26020 22812 26058
rect 22754 25986 22766 26020
rect 22800 25986 22812 26020
rect 22754 25948 22812 25986
rect 22754 25914 22766 25948
rect 22800 25914 22812 25948
rect 22754 25876 22812 25914
rect 22754 25842 22766 25876
rect 22800 25842 22812 25876
rect 22754 25814 22812 25842
rect 22868 26092 22920 26120
rect 22868 26058 22877 26092
rect 22911 26058 22920 26092
rect 22868 26020 22920 26058
rect 22868 25986 22877 26020
rect 22911 25986 22920 26020
rect 22868 25948 22920 25986
rect 22868 25936 22877 25948
rect 22911 25936 22920 25948
rect 22868 25876 22920 25884
rect 22868 25872 22877 25876
rect 22911 25872 22920 25876
rect 22868 25814 22920 25820
rect 22954 26114 23006 26120
rect 22954 26058 22963 26062
rect 22997 26058 23006 26062
rect 22954 26050 23006 26058
rect 22954 25986 22963 25998
rect 22997 25986 23006 25998
rect 22954 25948 23006 25986
rect 22954 25914 22963 25948
rect 22997 25914 23006 25948
rect 22954 25876 23006 25914
rect 22954 25842 22963 25876
rect 22997 25842 23006 25876
rect 22954 25814 23006 25842
rect 23040 26092 23092 26120
rect 23040 26058 23049 26092
rect 23083 26058 23092 26092
rect 23040 26020 23092 26058
rect 23040 25986 23049 26020
rect 23083 25986 23092 26020
rect 23040 25948 23092 25986
rect 23040 25936 23049 25948
rect 23083 25936 23092 25948
rect 23040 25876 23092 25884
rect 23040 25872 23049 25876
rect 23083 25872 23092 25876
rect 23040 25814 23092 25820
rect 23148 26092 23206 26120
rect 23148 26058 23160 26092
rect 23194 26058 23206 26092
rect 23148 26020 23206 26058
rect 23148 25986 23160 26020
rect 23194 25986 23206 26020
rect 23148 25948 23206 25986
rect 23148 25914 23160 25948
rect 23194 25914 23206 25948
rect 23148 25876 23206 25914
rect 23148 25842 23160 25876
rect 23194 25842 23206 25876
rect 23148 25814 23206 25842
rect 22766 25640 22800 25814
rect 22879 25764 23081 25776
rect 22879 25730 22891 25764
rect 22925 25730 22963 25764
rect 22997 25730 23035 25764
rect 23069 25730 23081 25764
rect 22879 25710 23081 25730
rect 22879 25650 22893 25710
rect 23067 25650 23081 25710
rect 13960 25580 14000 25640
rect 13560 22750 14000 25580
rect 22760 25580 22800 25640
rect 23160 25640 23194 25814
rect 23304 25726 23314 26158
rect 23384 25726 23394 26158
rect 31766 25726 31776 26158
rect 31846 25726 31856 26158
rect 31954 26092 32012 26120
rect 31954 26058 31966 26092
rect 32000 26058 32012 26092
rect 31954 26020 32012 26058
rect 31954 25986 31966 26020
rect 32000 25986 32012 26020
rect 31954 25948 32012 25986
rect 31954 25914 31966 25948
rect 32000 25914 32012 25948
rect 31954 25876 32012 25914
rect 31954 25842 31966 25876
rect 32000 25842 32012 25876
rect 31954 25814 32012 25842
rect 32068 26092 32120 26120
rect 32068 26058 32077 26092
rect 32111 26058 32120 26092
rect 32068 26020 32120 26058
rect 32068 25986 32077 26020
rect 32111 25986 32120 26020
rect 32068 25948 32120 25986
rect 32068 25936 32077 25948
rect 32111 25936 32120 25948
rect 32068 25876 32120 25884
rect 32068 25872 32077 25876
rect 32111 25872 32120 25876
rect 32068 25814 32120 25820
rect 32154 26114 32206 26120
rect 32154 26058 32163 26062
rect 32197 26058 32206 26062
rect 32154 26050 32206 26058
rect 32154 25986 32163 25998
rect 32197 25986 32206 25998
rect 32154 25948 32206 25986
rect 32154 25914 32163 25948
rect 32197 25914 32206 25948
rect 32154 25876 32206 25914
rect 32154 25842 32163 25876
rect 32197 25842 32206 25876
rect 32154 25814 32206 25842
rect 32240 26092 32292 26120
rect 32240 26058 32249 26092
rect 32283 26058 32292 26092
rect 32240 26020 32292 26058
rect 32240 25986 32249 26020
rect 32283 25986 32292 26020
rect 32240 25948 32292 25986
rect 32240 25936 32249 25948
rect 32283 25936 32292 25948
rect 32240 25876 32292 25884
rect 32240 25872 32249 25876
rect 32283 25872 32292 25876
rect 32240 25814 32292 25820
rect 32348 26092 32406 26120
rect 32348 26058 32360 26092
rect 32394 26058 32406 26092
rect 32348 26020 32406 26058
rect 32348 25986 32360 26020
rect 32394 25986 32406 26020
rect 32348 25948 32406 25986
rect 32348 25914 32360 25948
rect 32394 25914 32406 25948
rect 32348 25876 32406 25914
rect 32348 25842 32360 25876
rect 32394 25842 32406 25876
rect 32348 25814 32406 25842
rect 31966 25640 32000 25814
rect 32079 25764 32281 25776
rect 32079 25730 32091 25764
rect 32125 25730 32163 25764
rect 32197 25730 32235 25764
rect 32269 25730 32281 25764
rect 32079 25710 32281 25730
rect 32079 25650 32093 25710
rect 32267 25650 32281 25710
rect 23160 25580 23200 25640
rect 22760 22750 23200 25580
rect 31960 25580 32000 25640
rect 32360 25640 32394 25814
rect 32504 25726 32514 26158
rect 32584 25726 32594 26158
rect 40966 25726 40976 26158
rect 41046 25726 41056 26158
rect 41154 26092 41212 26120
rect 41154 26058 41166 26092
rect 41200 26058 41212 26092
rect 41154 26020 41212 26058
rect 41154 25986 41166 26020
rect 41200 25986 41212 26020
rect 41154 25948 41212 25986
rect 41154 25914 41166 25948
rect 41200 25914 41212 25948
rect 41154 25876 41212 25914
rect 41154 25842 41166 25876
rect 41200 25842 41212 25876
rect 41154 25814 41212 25842
rect 41268 26092 41320 26120
rect 41268 26058 41277 26092
rect 41311 26058 41320 26092
rect 41268 26020 41320 26058
rect 41268 25986 41277 26020
rect 41311 25986 41320 26020
rect 41268 25948 41320 25986
rect 41268 25936 41277 25948
rect 41311 25936 41320 25948
rect 41268 25876 41320 25884
rect 41268 25872 41277 25876
rect 41311 25872 41320 25876
rect 41268 25814 41320 25820
rect 41354 26114 41406 26120
rect 41354 26058 41363 26062
rect 41397 26058 41406 26062
rect 41354 26050 41406 26058
rect 41354 25986 41363 25998
rect 41397 25986 41406 25998
rect 41354 25948 41406 25986
rect 41354 25914 41363 25948
rect 41397 25914 41406 25948
rect 41354 25876 41406 25914
rect 41354 25842 41363 25876
rect 41397 25842 41406 25876
rect 41354 25814 41406 25842
rect 41440 26092 41492 26120
rect 41440 26058 41449 26092
rect 41483 26058 41492 26092
rect 41440 26020 41492 26058
rect 41440 25986 41449 26020
rect 41483 25986 41492 26020
rect 41440 25948 41492 25986
rect 41440 25936 41449 25948
rect 41483 25936 41492 25948
rect 41440 25876 41492 25884
rect 41440 25872 41449 25876
rect 41483 25872 41492 25876
rect 41440 25814 41492 25820
rect 41548 26092 41606 26120
rect 41548 26058 41560 26092
rect 41594 26058 41606 26092
rect 41548 26020 41606 26058
rect 41548 25986 41560 26020
rect 41594 25986 41606 26020
rect 41548 25948 41606 25986
rect 41548 25914 41560 25948
rect 41594 25914 41606 25948
rect 41548 25876 41606 25914
rect 41548 25842 41560 25876
rect 41594 25842 41606 25876
rect 41548 25814 41606 25842
rect 41166 25640 41200 25814
rect 41279 25764 41481 25776
rect 41279 25730 41291 25764
rect 41325 25730 41363 25764
rect 41397 25730 41435 25764
rect 41469 25730 41481 25764
rect 41279 25710 41481 25730
rect 41279 25650 41293 25710
rect 41467 25650 41481 25710
rect 32360 25580 32400 25640
rect 31960 22750 32400 25580
rect 41160 25580 41200 25640
rect 41560 25640 41594 25814
rect 41704 25726 41714 26158
rect 41784 25726 41794 26158
rect 50166 25726 50176 26158
rect 50246 25726 50256 26158
rect 50354 26092 50412 26120
rect 50354 26058 50366 26092
rect 50400 26058 50412 26092
rect 50354 26020 50412 26058
rect 50354 25986 50366 26020
rect 50400 25986 50412 26020
rect 50354 25948 50412 25986
rect 50354 25914 50366 25948
rect 50400 25914 50412 25948
rect 50354 25876 50412 25914
rect 50354 25842 50366 25876
rect 50400 25842 50412 25876
rect 50354 25814 50412 25842
rect 50468 26092 50520 26120
rect 50468 26058 50477 26092
rect 50511 26058 50520 26092
rect 50468 26020 50520 26058
rect 50468 25986 50477 26020
rect 50511 25986 50520 26020
rect 50468 25948 50520 25986
rect 50468 25936 50477 25948
rect 50511 25936 50520 25948
rect 50468 25876 50520 25884
rect 50468 25872 50477 25876
rect 50511 25872 50520 25876
rect 50468 25814 50520 25820
rect 50554 26114 50606 26120
rect 50554 26058 50563 26062
rect 50597 26058 50606 26062
rect 50554 26050 50606 26058
rect 50554 25986 50563 25998
rect 50597 25986 50606 25998
rect 50554 25948 50606 25986
rect 50554 25914 50563 25948
rect 50597 25914 50606 25948
rect 50554 25876 50606 25914
rect 50554 25842 50563 25876
rect 50597 25842 50606 25876
rect 50554 25814 50606 25842
rect 50640 26092 50692 26120
rect 50640 26058 50649 26092
rect 50683 26058 50692 26092
rect 50640 26020 50692 26058
rect 50640 25986 50649 26020
rect 50683 25986 50692 26020
rect 50640 25948 50692 25986
rect 50640 25936 50649 25948
rect 50683 25936 50692 25948
rect 50640 25876 50692 25884
rect 50640 25872 50649 25876
rect 50683 25872 50692 25876
rect 50640 25814 50692 25820
rect 50748 26092 50806 26120
rect 50748 26058 50760 26092
rect 50794 26058 50806 26092
rect 50748 26020 50806 26058
rect 50748 25986 50760 26020
rect 50794 25986 50806 26020
rect 50748 25948 50806 25986
rect 50748 25914 50760 25948
rect 50794 25914 50806 25948
rect 50748 25876 50806 25914
rect 50748 25842 50760 25876
rect 50794 25842 50806 25876
rect 50748 25814 50806 25842
rect 50366 25640 50400 25814
rect 50479 25764 50681 25776
rect 50479 25730 50491 25764
rect 50525 25730 50563 25764
rect 50597 25730 50635 25764
rect 50669 25730 50681 25764
rect 50479 25710 50681 25730
rect 50479 25650 50493 25710
rect 50667 25650 50681 25710
rect 41560 25580 41600 25640
rect 41160 22750 41600 25580
rect 50360 25580 50400 25640
rect 50760 25640 50794 25814
rect 50904 25726 50914 26158
rect 50984 25726 50994 26158
rect 59366 25726 59376 26158
rect 59446 25726 59456 26158
rect 59554 26092 59612 26120
rect 59554 26058 59566 26092
rect 59600 26058 59612 26092
rect 59554 26020 59612 26058
rect 59554 25986 59566 26020
rect 59600 25986 59612 26020
rect 59554 25948 59612 25986
rect 59554 25914 59566 25948
rect 59600 25914 59612 25948
rect 59554 25876 59612 25914
rect 59554 25842 59566 25876
rect 59600 25842 59612 25876
rect 59554 25814 59612 25842
rect 59668 26092 59720 26120
rect 59668 26058 59677 26092
rect 59711 26058 59720 26092
rect 59668 26020 59720 26058
rect 59668 25986 59677 26020
rect 59711 25986 59720 26020
rect 59668 25948 59720 25986
rect 59668 25936 59677 25948
rect 59711 25936 59720 25948
rect 59668 25876 59720 25884
rect 59668 25872 59677 25876
rect 59711 25872 59720 25876
rect 59668 25814 59720 25820
rect 59754 26114 59806 26120
rect 59754 26058 59763 26062
rect 59797 26058 59806 26062
rect 59754 26050 59806 26058
rect 59754 25986 59763 25998
rect 59797 25986 59806 25998
rect 59754 25948 59806 25986
rect 59754 25914 59763 25948
rect 59797 25914 59806 25948
rect 59754 25876 59806 25914
rect 59754 25842 59763 25876
rect 59797 25842 59806 25876
rect 59754 25814 59806 25842
rect 59840 26092 59892 26120
rect 59840 26058 59849 26092
rect 59883 26058 59892 26092
rect 59840 26020 59892 26058
rect 59840 25986 59849 26020
rect 59883 25986 59892 26020
rect 59840 25948 59892 25986
rect 59840 25936 59849 25948
rect 59883 25936 59892 25948
rect 59840 25876 59892 25884
rect 59840 25872 59849 25876
rect 59883 25872 59892 25876
rect 59840 25814 59892 25820
rect 59948 26092 60006 26120
rect 59948 26058 59960 26092
rect 59994 26058 60006 26092
rect 59948 26020 60006 26058
rect 59948 25986 59960 26020
rect 59994 25986 60006 26020
rect 59948 25948 60006 25986
rect 59948 25914 59960 25948
rect 59994 25914 60006 25948
rect 59948 25876 60006 25914
rect 59948 25842 59960 25876
rect 59994 25842 60006 25876
rect 59948 25814 60006 25842
rect 59566 25640 59600 25814
rect 59679 25764 59881 25776
rect 59679 25730 59691 25764
rect 59725 25730 59763 25764
rect 59797 25730 59835 25764
rect 59869 25730 59881 25764
rect 59679 25710 59881 25730
rect 59679 25650 59693 25710
rect 59867 25650 59881 25710
rect 50760 25580 50800 25640
rect 50360 22750 50800 25580
rect 59560 25580 59600 25640
rect 59960 25640 59994 25814
rect 60104 25726 60114 26158
rect 60184 25726 60194 26158
rect 68566 25726 68576 26158
rect 68646 25726 68656 26158
rect 68754 26092 68812 26120
rect 68754 26058 68766 26092
rect 68800 26058 68812 26092
rect 68754 26020 68812 26058
rect 68754 25986 68766 26020
rect 68800 25986 68812 26020
rect 68754 25948 68812 25986
rect 68754 25914 68766 25948
rect 68800 25914 68812 25948
rect 68754 25876 68812 25914
rect 68754 25842 68766 25876
rect 68800 25842 68812 25876
rect 68754 25814 68812 25842
rect 68868 26092 68920 26120
rect 68868 26058 68877 26092
rect 68911 26058 68920 26092
rect 68868 26020 68920 26058
rect 68868 25986 68877 26020
rect 68911 25986 68920 26020
rect 68868 25948 68920 25986
rect 68868 25936 68877 25948
rect 68911 25936 68920 25948
rect 68868 25876 68920 25884
rect 68868 25872 68877 25876
rect 68911 25872 68920 25876
rect 68868 25814 68920 25820
rect 68954 26114 69006 26120
rect 68954 26058 68963 26062
rect 68997 26058 69006 26062
rect 68954 26050 69006 26058
rect 68954 25986 68963 25998
rect 68997 25986 69006 25998
rect 68954 25948 69006 25986
rect 68954 25914 68963 25948
rect 68997 25914 69006 25948
rect 68954 25876 69006 25914
rect 68954 25842 68963 25876
rect 68997 25842 69006 25876
rect 68954 25814 69006 25842
rect 69040 26092 69092 26120
rect 69040 26058 69049 26092
rect 69083 26058 69092 26092
rect 69040 26020 69092 26058
rect 69040 25986 69049 26020
rect 69083 25986 69092 26020
rect 69040 25948 69092 25986
rect 69040 25936 69049 25948
rect 69083 25936 69092 25948
rect 69040 25876 69092 25884
rect 69040 25872 69049 25876
rect 69083 25872 69092 25876
rect 69040 25814 69092 25820
rect 69148 26092 69206 26120
rect 69148 26058 69160 26092
rect 69194 26058 69206 26092
rect 69148 26020 69206 26058
rect 69148 25986 69160 26020
rect 69194 25986 69206 26020
rect 69148 25948 69206 25986
rect 69148 25914 69160 25948
rect 69194 25914 69206 25948
rect 69148 25876 69206 25914
rect 69148 25842 69160 25876
rect 69194 25842 69206 25876
rect 69148 25814 69206 25842
rect 68766 25640 68800 25814
rect 68879 25764 69081 25776
rect 68879 25730 68891 25764
rect 68925 25730 68963 25764
rect 68997 25730 69035 25764
rect 69069 25730 69081 25764
rect 68879 25710 69081 25730
rect 68879 25650 68893 25710
rect 69067 25650 69081 25710
rect 59960 25580 60000 25640
rect 59560 22750 60000 25580
rect 68760 25580 68800 25640
rect 69160 25640 69194 25814
rect 69304 25726 69314 26158
rect 69384 25726 69394 26158
rect 69160 25580 69200 25640
rect 68760 22750 69200 25580
rect -3880 20750 73600 22750
rect -3880 12870 -1870 20750
rect 75600 18750 77600 26630
rect 0 16892 77600 18750
rect 0 16750 4192 16892
rect 4186 16495 4192 16750
rect 4230 16750 4930 16892
rect 4230 16495 4236 16750
rect 4186 16483 4236 16495
rect 4924 16495 4930 16750
rect 4968 16750 13392 16892
rect 4968 16495 4974 16750
rect 4924 16483 4974 16495
rect 13386 16495 13392 16750
rect 13430 16750 14130 16892
rect 13430 16495 13436 16750
rect 13386 16483 13436 16495
rect 14124 16495 14130 16750
rect 14168 16750 22592 16892
rect 14168 16495 14174 16750
rect 14124 16483 14174 16495
rect 22586 16495 22592 16750
rect 22630 16750 23330 16892
rect 22630 16495 22636 16750
rect 22586 16483 22636 16495
rect 23324 16495 23330 16750
rect 23368 16750 31792 16892
rect 23368 16495 23374 16750
rect 23324 16483 23374 16495
rect 31786 16495 31792 16750
rect 31830 16750 32530 16892
rect 31830 16495 31836 16750
rect 31786 16483 31836 16495
rect 32524 16495 32530 16750
rect 32568 16750 40992 16892
rect 32568 16495 32574 16750
rect 32524 16483 32574 16495
rect 40986 16495 40992 16750
rect 41030 16750 41730 16892
rect 41030 16495 41036 16750
rect 40986 16483 41036 16495
rect 41724 16495 41730 16750
rect 41768 16750 50192 16892
rect 41768 16495 41774 16750
rect 41724 16483 41774 16495
rect 50186 16495 50192 16750
rect 50230 16750 50930 16892
rect 50230 16495 50236 16750
rect 50186 16483 50236 16495
rect 50924 16495 50930 16750
rect 50968 16750 59392 16892
rect 50968 16495 50974 16750
rect 50924 16483 50974 16495
rect 59386 16495 59392 16750
rect 59430 16750 60130 16892
rect 59430 16495 59436 16750
rect 59386 16483 59436 16495
rect 60124 16495 60130 16750
rect 60168 16750 68592 16892
rect 60168 16495 60174 16750
rect 60124 16483 60174 16495
rect 68586 16495 68592 16750
rect 68630 16750 69330 16892
rect 68630 16495 68636 16750
rect 68586 16483 68636 16495
rect 69324 16495 69330 16750
rect 69368 16750 77600 16892
rect 69368 16495 69374 16750
rect 69324 16483 69374 16495
rect 4479 16324 4681 16344
rect 4479 16290 4491 16324
rect 4525 16290 4563 16324
rect 4597 16290 4635 16324
rect 4669 16290 4681 16324
rect 4479 16278 4681 16290
rect 13679 16324 13881 16344
rect 13679 16290 13691 16324
rect 13725 16290 13763 16324
rect 13797 16290 13835 16324
rect 13869 16290 13881 16324
rect 13679 16278 13881 16290
rect 22879 16324 23081 16344
rect 22879 16290 22891 16324
rect 22925 16290 22963 16324
rect 22997 16290 23035 16324
rect 23069 16290 23081 16324
rect 22879 16278 23081 16290
rect 32079 16324 32281 16344
rect 32079 16290 32091 16324
rect 32125 16290 32163 16324
rect 32197 16290 32235 16324
rect 32269 16290 32281 16324
rect 32079 16278 32281 16290
rect 41279 16324 41481 16344
rect 41279 16290 41291 16324
rect 41325 16290 41363 16324
rect 41397 16290 41435 16324
rect 41469 16290 41481 16324
rect 41279 16278 41481 16290
rect 50479 16324 50681 16344
rect 50479 16290 50491 16324
rect 50525 16290 50563 16324
rect 50597 16290 50635 16324
rect 50669 16290 50681 16324
rect 50479 16278 50681 16290
rect 59679 16324 59881 16344
rect 59679 16290 59691 16324
rect 59725 16290 59763 16324
rect 59797 16290 59835 16324
rect 59869 16290 59881 16324
rect 59679 16278 59881 16290
rect 68879 16324 69081 16344
rect 68879 16290 68891 16324
rect 68925 16290 68963 16324
rect 68997 16290 69035 16324
rect 69069 16290 69081 16324
rect 68879 16278 69081 16290
rect 4166 15846 4176 16278
rect 4246 15846 4256 16278
rect 4354 16212 4412 16240
rect 4354 16178 4366 16212
rect 4400 16178 4412 16212
rect 4354 16140 4412 16178
rect 4354 16106 4366 16140
rect 4400 16106 4412 16140
rect 4354 16068 4412 16106
rect 4354 16034 4366 16068
rect 4400 16034 4412 16068
rect 4354 15996 4412 16034
rect 4354 15962 4366 15996
rect 4400 15962 4412 15996
rect 4354 15934 4412 15962
rect 4468 16212 4520 16240
rect 4468 16178 4477 16212
rect 4511 16178 4520 16212
rect 4468 16140 4520 16178
rect 4468 16106 4477 16140
rect 4511 16106 4520 16140
rect 4468 16068 4520 16106
rect 4468 16056 4477 16068
rect 4511 16056 4520 16068
rect 4468 15996 4520 16004
rect 4468 15992 4477 15996
rect 4511 15992 4520 15996
rect 4468 15934 4520 15940
rect 4554 16234 4606 16240
rect 4554 16178 4563 16182
rect 4597 16178 4606 16182
rect 4554 16170 4606 16178
rect 4554 16106 4563 16118
rect 4597 16106 4606 16118
rect 4554 16068 4606 16106
rect 4554 16034 4563 16068
rect 4597 16034 4606 16068
rect 4554 15996 4606 16034
rect 4554 15962 4563 15996
rect 4597 15962 4606 15996
rect 4554 15934 4606 15962
rect 4640 16212 4692 16240
rect 4640 16178 4649 16212
rect 4683 16178 4692 16212
rect 4640 16140 4692 16178
rect 4640 16106 4649 16140
rect 4683 16106 4692 16140
rect 4640 16068 4692 16106
rect 4640 16056 4649 16068
rect 4683 16056 4692 16068
rect 4640 15996 4692 16004
rect 4640 15992 4649 15996
rect 4683 15992 4692 15996
rect 4640 15934 4692 15940
rect 4748 16212 4806 16240
rect 4748 16178 4760 16212
rect 4794 16178 4806 16212
rect 4748 16140 4806 16178
rect 4748 16106 4760 16140
rect 4794 16106 4806 16140
rect 4748 16068 4806 16106
rect 4748 16034 4760 16068
rect 4794 16034 4806 16068
rect 4748 15996 4806 16034
rect 4748 15962 4760 15996
rect 4794 15962 4806 15996
rect 4748 15934 4806 15962
rect 4366 15760 4400 15934
rect 4479 15884 4681 15896
rect 4479 15850 4491 15884
rect 4525 15850 4563 15884
rect 4597 15850 4635 15884
rect 4669 15850 4681 15884
rect 4479 15830 4681 15850
rect 4479 15770 4493 15830
rect 4667 15770 4681 15830
rect 4360 15700 4400 15760
rect 4760 15760 4794 15934
rect 4904 15846 4914 16278
rect 4984 15846 4994 16278
rect 13366 15846 13376 16278
rect 13446 15846 13456 16278
rect 13554 16212 13612 16240
rect 13554 16178 13566 16212
rect 13600 16178 13612 16212
rect 13554 16140 13612 16178
rect 13554 16106 13566 16140
rect 13600 16106 13612 16140
rect 13554 16068 13612 16106
rect 13554 16034 13566 16068
rect 13600 16034 13612 16068
rect 13554 15996 13612 16034
rect 13554 15962 13566 15996
rect 13600 15962 13612 15996
rect 13554 15934 13612 15962
rect 13668 16212 13720 16240
rect 13668 16178 13677 16212
rect 13711 16178 13720 16212
rect 13668 16140 13720 16178
rect 13668 16106 13677 16140
rect 13711 16106 13720 16140
rect 13668 16068 13720 16106
rect 13668 16056 13677 16068
rect 13711 16056 13720 16068
rect 13668 15996 13720 16004
rect 13668 15992 13677 15996
rect 13711 15992 13720 15996
rect 13668 15934 13720 15940
rect 13754 16234 13806 16240
rect 13754 16178 13763 16182
rect 13797 16178 13806 16182
rect 13754 16170 13806 16178
rect 13754 16106 13763 16118
rect 13797 16106 13806 16118
rect 13754 16068 13806 16106
rect 13754 16034 13763 16068
rect 13797 16034 13806 16068
rect 13754 15996 13806 16034
rect 13754 15962 13763 15996
rect 13797 15962 13806 15996
rect 13754 15934 13806 15962
rect 13840 16212 13892 16240
rect 13840 16178 13849 16212
rect 13883 16178 13892 16212
rect 13840 16140 13892 16178
rect 13840 16106 13849 16140
rect 13883 16106 13892 16140
rect 13840 16068 13892 16106
rect 13840 16056 13849 16068
rect 13883 16056 13892 16068
rect 13840 15996 13892 16004
rect 13840 15992 13849 15996
rect 13883 15992 13892 15996
rect 13840 15934 13892 15940
rect 13948 16212 14006 16240
rect 13948 16178 13960 16212
rect 13994 16178 14006 16212
rect 13948 16140 14006 16178
rect 13948 16106 13960 16140
rect 13994 16106 14006 16140
rect 13948 16068 14006 16106
rect 13948 16034 13960 16068
rect 13994 16034 14006 16068
rect 13948 15996 14006 16034
rect 13948 15962 13960 15996
rect 13994 15962 14006 15996
rect 13948 15934 14006 15962
rect 13566 15760 13600 15934
rect 13679 15884 13881 15896
rect 13679 15850 13691 15884
rect 13725 15850 13763 15884
rect 13797 15850 13835 15884
rect 13869 15850 13881 15884
rect 13679 15830 13881 15850
rect 13679 15770 13693 15830
rect 13867 15770 13881 15830
rect 4760 15700 4800 15760
rect 4360 12870 4800 15700
rect 13560 15700 13600 15760
rect 13960 15760 13994 15934
rect 14104 15846 14114 16278
rect 14184 15846 14194 16278
rect 22566 15846 22576 16278
rect 22646 15846 22656 16278
rect 22754 16212 22812 16240
rect 22754 16178 22766 16212
rect 22800 16178 22812 16212
rect 22754 16140 22812 16178
rect 22754 16106 22766 16140
rect 22800 16106 22812 16140
rect 22754 16068 22812 16106
rect 22754 16034 22766 16068
rect 22800 16034 22812 16068
rect 22754 15996 22812 16034
rect 22754 15962 22766 15996
rect 22800 15962 22812 15996
rect 22754 15934 22812 15962
rect 22868 16212 22920 16240
rect 22868 16178 22877 16212
rect 22911 16178 22920 16212
rect 22868 16140 22920 16178
rect 22868 16106 22877 16140
rect 22911 16106 22920 16140
rect 22868 16068 22920 16106
rect 22868 16056 22877 16068
rect 22911 16056 22920 16068
rect 22868 15996 22920 16004
rect 22868 15992 22877 15996
rect 22911 15992 22920 15996
rect 22868 15934 22920 15940
rect 22954 16234 23006 16240
rect 22954 16178 22963 16182
rect 22997 16178 23006 16182
rect 22954 16170 23006 16178
rect 22954 16106 22963 16118
rect 22997 16106 23006 16118
rect 22954 16068 23006 16106
rect 22954 16034 22963 16068
rect 22997 16034 23006 16068
rect 22954 15996 23006 16034
rect 22954 15962 22963 15996
rect 22997 15962 23006 15996
rect 22954 15934 23006 15962
rect 23040 16212 23092 16240
rect 23040 16178 23049 16212
rect 23083 16178 23092 16212
rect 23040 16140 23092 16178
rect 23040 16106 23049 16140
rect 23083 16106 23092 16140
rect 23040 16068 23092 16106
rect 23040 16056 23049 16068
rect 23083 16056 23092 16068
rect 23040 15996 23092 16004
rect 23040 15992 23049 15996
rect 23083 15992 23092 15996
rect 23040 15934 23092 15940
rect 23148 16212 23206 16240
rect 23148 16178 23160 16212
rect 23194 16178 23206 16212
rect 23148 16140 23206 16178
rect 23148 16106 23160 16140
rect 23194 16106 23206 16140
rect 23148 16068 23206 16106
rect 23148 16034 23160 16068
rect 23194 16034 23206 16068
rect 23148 15996 23206 16034
rect 23148 15962 23160 15996
rect 23194 15962 23206 15996
rect 23148 15934 23206 15962
rect 22766 15760 22800 15934
rect 22879 15884 23081 15896
rect 22879 15850 22891 15884
rect 22925 15850 22963 15884
rect 22997 15850 23035 15884
rect 23069 15850 23081 15884
rect 22879 15830 23081 15850
rect 22879 15770 22893 15830
rect 23067 15770 23081 15830
rect 13960 15700 14000 15760
rect 13560 12870 14000 15700
rect 22760 15700 22800 15760
rect 23160 15760 23194 15934
rect 23304 15846 23314 16278
rect 23384 15846 23394 16278
rect 31766 15846 31776 16278
rect 31846 15846 31856 16278
rect 31954 16212 32012 16240
rect 31954 16178 31966 16212
rect 32000 16178 32012 16212
rect 31954 16140 32012 16178
rect 31954 16106 31966 16140
rect 32000 16106 32012 16140
rect 31954 16068 32012 16106
rect 31954 16034 31966 16068
rect 32000 16034 32012 16068
rect 31954 15996 32012 16034
rect 31954 15962 31966 15996
rect 32000 15962 32012 15996
rect 31954 15934 32012 15962
rect 32068 16212 32120 16240
rect 32068 16178 32077 16212
rect 32111 16178 32120 16212
rect 32068 16140 32120 16178
rect 32068 16106 32077 16140
rect 32111 16106 32120 16140
rect 32068 16068 32120 16106
rect 32068 16056 32077 16068
rect 32111 16056 32120 16068
rect 32068 15996 32120 16004
rect 32068 15992 32077 15996
rect 32111 15992 32120 15996
rect 32068 15934 32120 15940
rect 32154 16234 32206 16240
rect 32154 16178 32163 16182
rect 32197 16178 32206 16182
rect 32154 16170 32206 16178
rect 32154 16106 32163 16118
rect 32197 16106 32206 16118
rect 32154 16068 32206 16106
rect 32154 16034 32163 16068
rect 32197 16034 32206 16068
rect 32154 15996 32206 16034
rect 32154 15962 32163 15996
rect 32197 15962 32206 15996
rect 32154 15934 32206 15962
rect 32240 16212 32292 16240
rect 32240 16178 32249 16212
rect 32283 16178 32292 16212
rect 32240 16140 32292 16178
rect 32240 16106 32249 16140
rect 32283 16106 32292 16140
rect 32240 16068 32292 16106
rect 32240 16056 32249 16068
rect 32283 16056 32292 16068
rect 32240 15996 32292 16004
rect 32240 15992 32249 15996
rect 32283 15992 32292 15996
rect 32240 15934 32292 15940
rect 32348 16212 32406 16240
rect 32348 16178 32360 16212
rect 32394 16178 32406 16212
rect 32348 16140 32406 16178
rect 32348 16106 32360 16140
rect 32394 16106 32406 16140
rect 32348 16068 32406 16106
rect 32348 16034 32360 16068
rect 32394 16034 32406 16068
rect 32348 15996 32406 16034
rect 32348 15962 32360 15996
rect 32394 15962 32406 15996
rect 32348 15934 32406 15962
rect 31966 15760 32000 15934
rect 32079 15884 32281 15896
rect 32079 15850 32091 15884
rect 32125 15850 32163 15884
rect 32197 15850 32235 15884
rect 32269 15850 32281 15884
rect 32079 15830 32281 15850
rect 32079 15770 32093 15830
rect 32267 15770 32281 15830
rect 23160 15700 23200 15760
rect 22760 12870 23200 15700
rect 31960 15700 32000 15760
rect 32360 15760 32394 15934
rect 32504 15846 32514 16278
rect 32584 15846 32594 16278
rect 40966 15846 40976 16278
rect 41046 15846 41056 16278
rect 41154 16212 41212 16240
rect 41154 16178 41166 16212
rect 41200 16178 41212 16212
rect 41154 16140 41212 16178
rect 41154 16106 41166 16140
rect 41200 16106 41212 16140
rect 41154 16068 41212 16106
rect 41154 16034 41166 16068
rect 41200 16034 41212 16068
rect 41154 15996 41212 16034
rect 41154 15962 41166 15996
rect 41200 15962 41212 15996
rect 41154 15934 41212 15962
rect 41268 16212 41320 16240
rect 41268 16178 41277 16212
rect 41311 16178 41320 16212
rect 41268 16140 41320 16178
rect 41268 16106 41277 16140
rect 41311 16106 41320 16140
rect 41268 16068 41320 16106
rect 41268 16056 41277 16068
rect 41311 16056 41320 16068
rect 41268 15996 41320 16004
rect 41268 15992 41277 15996
rect 41311 15992 41320 15996
rect 41268 15934 41320 15940
rect 41354 16234 41406 16240
rect 41354 16178 41363 16182
rect 41397 16178 41406 16182
rect 41354 16170 41406 16178
rect 41354 16106 41363 16118
rect 41397 16106 41406 16118
rect 41354 16068 41406 16106
rect 41354 16034 41363 16068
rect 41397 16034 41406 16068
rect 41354 15996 41406 16034
rect 41354 15962 41363 15996
rect 41397 15962 41406 15996
rect 41354 15934 41406 15962
rect 41440 16212 41492 16240
rect 41440 16178 41449 16212
rect 41483 16178 41492 16212
rect 41440 16140 41492 16178
rect 41440 16106 41449 16140
rect 41483 16106 41492 16140
rect 41440 16068 41492 16106
rect 41440 16056 41449 16068
rect 41483 16056 41492 16068
rect 41440 15996 41492 16004
rect 41440 15992 41449 15996
rect 41483 15992 41492 15996
rect 41440 15934 41492 15940
rect 41548 16212 41606 16240
rect 41548 16178 41560 16212
rect 41594 16178 41606 16212
rect 41548 16140 41606 16178
rect 41548 16106 41560 16140
rect 41594 16106 41606 16140
rect 41548 16068 41606 16106
rect 41548 16034 41560 16068
rect 41594 16034 41606 16068
rect 41548 15996 41606 16034
rect 41548 15962 41560 15996
rect 41594 15962 41606 15996
rect 41548 15934 41606 15962
rect 41166 15760 41200 15934
rect 41279 15884 41481 15896
rect 41279 15850 41291 15884
rect 41325 15850 41363 15884
rect 41397 15850 41435 15884
rect 41469 15850 41481 15884
rect 41279 15830 41481 15850
rect 41279 15770 41293 15830
rect 41467 15770 41481 15830
rect 32360 15700 32400 15760
rect 31960 12870 32400 15700
rect 41160 15700 41200 15760
rect 41560 15760 41594 15934
rect 41704 15846 41714 16278
rect 41784 15846 41794 16278
rect 50166 15846 50176 16278
rect 50246 15846 50256 16278
rect 50354 16212 50412 16240
rect 50354 16178 50366 16212
rect 50400 16178 50412 16212
rect 50354 16140 50412 16178
rect 50354 16106 50366 16140
rect 50400 16106 50412 16140
rect 50354 16068 50412 16106
rect 50354 16034 50366 16068
rect 50400 16034 50412 16068
rect 50354 15996 50412 16034
rect 50354 15962 50366 15996
rect 50400 15962 50412 15996
rect 50354 15934 50412 15962
rect 50468 16212 50520 16240
rect 50468 16178 50477 16212
rect 50511 16178 50520 16212
rect 50468 16140 50520 16178
rect 50468 16106 50477 16140
rect 50511 16106 50520 16140
rect 50468 16068 50520 16106
rect 50468 16056 50477 16068
rect 50511 16056 50520 16068
rect 50468 15996 50520 16004
rect 50468 15992 50477 15996
rect 50511 15992 50520 15996
rect 50468 15934 50520 15940
rect 50554 16234 50606 16240
rect 50554 16178 50563 16182
rect 50597 16178 50606 16182
rect 50554 16170 50606 16178
rect 50554 16106 50563 16118
rect 50597 16106 50606 16118
rect 50554 16068 50606 16106
rect 50554 16034 50563 16068
rect 50597 16034 50606 16068
rect 50554 15996 50606 16034
rect 50554 15962 50563 15996
rect 50597 15962 50606 15996
rect 50554 15934 50606 15962
rect 50640 16212 50692 16240
rect 50640 16178 50649 16212
rect 50683 16178 50692 16212
rect 50640 16140 50692 16178
rect 50640 16106 50649 16140
rect 50683 16106 50692 16140
rect 50640 16068 50692 16106
rect 50640 16056 50649 16068
rect 50683 16056 50692 16068
rect 50640 15996 50692 16004
rect 50640 15992 50649 15996
rect 50683 15992 50692 15996
rect 50640 15934 50692 15940
rect 50748 16212 50806 16240
rect 50748 16178 50760 16212
rect 50794 16178 50806 16212
rect 50748 16140 50806 16178
rect 50748 16106 50760 16140
rect 50794 16106 50806 16140
rect 50748 16068 50806 16106
rect 50748 16034 50760 16068
rect 50794 16034 50806 16068
rect 50748 15996 50806 16034
rect 50748 15962 50760 15996
rect 50794 15962 50806 15996
rect 50748 15934 50806 15962
rect 50366 15760 50400 15934
rect 50479 15884 50681 15896
rect 50479 15850 50491 15884
rect 50525 15850 50563 15884
rect 50597 15850 50635 15884
rect 50669 15850 50681 15884
rect 50479 15830 50681 15850
rect 50479 15770 50493 15830
rect 50667 15770 50681 15830
rect 41560 15700 41600 15760
rect 41160 12870 41600 15700
rect 50360 15700 50400 15760
rect 50760 15760 50794 15934
rect 50904 15846 50914 16278
rect 50984 15846 50994 16278
rect 59366 15846 59376 16278
rect 59446 15846 59456 16278
rect 59554 16212 59612 16240
rect 59554 16178 59566 16212
rect 59600 16178 59612 16212
rect 59554 16140 59612 16178
rect 59554 16106 59566 16140
rect 59600 16106 59612 16140
rect 59554 16068 59612 16106
rect 59554 16034 59566 16068
rect 59600 16034 59612 16068
rect 59554 15996 59612 16034
rect 59554 15962 59566 15996
rect 59600 15962 59612 15996
rect 59554 15934 59612 15962
rect 59668 16212 59720 16240
rect 59668 16178 59677 16212
rect 59711 16178 59720 16212
rect 59668 16140 59720 16178
rect 59668 16106 59677 16140
rect 59711 16106 59720 16140
rect 59668 16068 59720 16106
rect 59668 16056 59677 16068
rect 59711 16056 59720 16068
rect 59668 15996 59720 16004
rect 59668 15992 59677 15996
rect 59711 15992 59720 15996
rect 59668 15934 59720 15940
rect 59754 16234 59806 16240
rect 59754 16178 59763 16182
rect 59797 16178 59806 16182
rect 59754 16170 59806 16178
rect 59754 16106 59763 16118
rect 59797 16106 59806 16118
rect 59754 16068 59806 16106
rect 59754 16034 59763 16068
rect 59797 16034 59806 16068
rect 59754 15996 59806 16034
rect 59754 15962 59763 15996
rect 59797 15962 59806 15996
rect 59754 15934 59806 15962
rect 59840 16212 59892 16240
rect 59840 16178 59849 16212
rect 59883 16178 59892 16212
rect 59840 16140 59892 16178
rect 59840 16106 59849 16140
rect 59883 16106 59892 16140
rect 59840 16068 59892 16106
rect 59840 16056 59849 16068
rect 59883 16056 59892 16068
rect 59840 15996 59892 16004
rect 59840 15992 59849 15996
rect 59883 15992 59892 15996
rect 59840 15934 59892 15940
rect 59948 16212 60006 16240
rect 59948 16178 59960 16212
rect 59994 16178 60006 16212
rect 59948 16140 60006 16178
rect 59948 16106 59960 16140
rect 59994 16106 60006 16140
rect 59948 16068 60006 16106
rect 59948 16034 59960 16068
rect 59994 16034 60006 16068
rect 59948 15996 60006 16034
rect 59948 15962 59960 15996
rect 59994 15962 60006 15996
rect 59948 15934 60006 15962
rect 59566 15760 59600 15934
rect 59679 15884 59881 15896
rect 59679 15850 59691 15884
rect 59725 15850 59763 15884
rect 59797 15850 59835 15884
rect 59869 15850 59881 15884
rect 59679 15830 59881 15850
rect 59679 15770 59693 15830
rect 59867 15770 59881 15830
rect 50760 15700 50800 15760
rect 50360 12870 50800 15700
rect 59560 15700 59600 15760
rect 59960 15760 59994 15934
rect 60104 15846 60114 16278
rect 60184 15846 60194 16278
rect 68566 15846 68576 16278
rect 68646 15846 68656 16278
rect 68754 16212 68812 16240
rect 68754 16178 68766 16212
rect 68800 16178 68812 16212
rect 68754 16140 68812 16178
rect 68754 16106 68766 16140
rect 68800 16106 68812 16140
rect 68754 16068 68812 16106
rect 68754 16034 68766 16068
rect 68800 16034 68812 16068
rect 68754 15996 68812 16034
rect 68754 15962 68766 15996
rect 68800 15962 68812 15996
rect 68754 15934 68812 15962
rect 68868 16212 68920 16240
rect 68868 16178 68877 16212
rect 68911 16178 68920 16212
rect 68868 16140 68920 16178
rect 68868 16106 68877 16140
rect 68911 16106 68920 16140
rect 68868 16068 68920 16106
rect 68868 16056 68877 16068
rect 68911 16056 68920 16068
rect 68868 15996 68920 16004
rect 68868 15992 68877 15996
rect 68911 15992 68920 15996
rect 68868 15934 68920 15940
rect 68954 16234 69006 16240
rect 68954 16178 68963 16182
rect 68997 16178 69006 16182
rect 68954 16170 69006 16178
rect 68954 16106 68963 16118
rect 68997 16106 69006 16118
rect 68954 16068 69006 16106
rect 68954 16034 68963 16068
rect 68997 16034 69006 16068
rect 68954 15996 69006 16034
rect 68954 15962 68963 15996
rect 68997 15962 69006 15996
rect 68954 15934 69006 15962
rect 69040 16212 69092 16240
rect 69040 16178 69049 16212
rect 69083 16178 69092 16212
rect 69040 16140 69092 16178
rect 69040 16106 69049 16140
rect 69083 16106 69092 16140
rect 69040 16068 69092 16106
rect 69040 16056 69049 16068
rect 69083 16056 69092 16068
rect 69040 15996 69092 16004
rect 69040 15992 69049 15996
rect 69083 15992 69092 15996
rect 69040 15934 69092 15940
rect 69148 16212 69206 16240
rect 69148 16178 69160 16212
rect 69194 16178 69206 16212
rect 69148 16140 69206 16178
rect 69148 16106 69160 16140
rect 69194 16106 69206 16140
rect 69148 16068 69206 16106
rect 69148 16034 69160 16068
rect 69194 16034 69206 16068
rect 69148 15996 69206 16034
rect 69148 15962 69160 15996
rect 69194 15962 69206 15996
rect 69148 15934 69206 15962
rect 68766 15760 68800 15934
rect 68879 15884 69081 15896
rect 68879 15850 68891 15884
rect 68925 15850 68963 15884
rect 68997 15850 69035 15884
rect 69069 15850 69081 15884
rect 68879 15830 69081 15850
rect 68879 15770 68893 15830
rect 69067 15770 69081 15830
rect 59960 15700 60000 15760
rect 59560 12870 60000 15700
rect 68760 15700 68800 15760
rect 69160 15760 69194 15934
rect 69304 15846 69314 16278
rect 69384 15846 69394 16278
rect 69160 15700 69200 15760
rect 68760 12870 69200 15700
rect -3880 10870 73600 12870
rect -3880 5380 -1870 10870
rect 75600 8870 77600 16750
rect -610 7012 77600 8870
rect -610 6870 4192 7012
rect -610 5840 -550 6870
rect -510 6620 -220 6640
rect -510 6560 -490 6620
rect -240 6560 -220 6620
rect 4186 6615 4192 6870
rect 4230 6870 4930 7012
rect 4230 6615 4236 6870
rect 4186 6603 4236 6615
rect 4924 6615 4930 6870
rect 4968 6870 13392 7012
rect 4968 6615 4974 6870
rect 4924 6603 4974 6615
rect 13386 6615 13392 6870
rect 13430 6870 14130 7012
rect 13430 6615 13436 6870
rect 13386 6603 13436 6615
rect 14124 6615 14130 6870
rect 14168 6870 22592 7012
rect 14168 6615 14174 6870
rect 14124 6603 14174 6615
rect 22586 6615 22592 6870
rect 22630 6870 23330 7012
rect 22630 6615 22636 6870
rect 22586 6603 22636 6615
rect 23324 6615 23330 6870
rect 23368 6870 31792 7012
rect 23368 6615 23374 6870
rect 23324 6603 23374 6615
rect 31786 6615 31792 6870
rect 31830 6870 32530 7012
rect 31830 6615 31836 6870
rect 31786 6603 31836 6615
rect 32524 6615 32530 6870
rect 32568 6870 40992 7012
rect 32568 6615 32574 6870
rect 32524 6603 32574 6615
rect 40986 6615 40992 6870
rect 41030 6870 41730 7012
rect 41030 6615 41036 6870
rect 40986 6603 41036 6615
rect 41724 6615 41730 6870
rect 41768 6870 50192 7012
rect 41768 6615 41774 6870
rect 41724 6603 41774 6615
rect 50186 6615 50192 6870
rect 50230 6870 50930 7012
rect 50230 6615 50236 6870
rect 50186 6603 50236 6615
rect 50924 6615 50930 6870
rect 50968 6870 59392 7012
rect 50968 6615 50974 6870
rect 50924 6603 50974 6615
rect 59386 6615 59392 6870
rect 59430 6870 60130 7012
rect 59430 6615 59436 6870
rect 59386 6603 59436 6615
rect 60124 6615 60130 6870
rect 60168 6870 68592 7012
rect 60168 6615 60174 6870
rect 60124 6603 60174 6615
rect 68586 6615 68592 6870
rect 68630 6870 69330 7012
rect 68630 6615 68636 6870
rect 68586 6603 68636 6615
rect 69324 6615 69330 6870
rect 69368 6870 77600 7012
rect 69368 6615 69374 6870
rect 69324 6603 69374 6615
rect -510 6540 -220 6560
rect -430 6464 -384 6476
rect -430 5888 -424 6464
rect -390 5888 -384 6464
rect -430 5876 -384 5888
rect -342 6464 -296 6476
rect -342 5888 -336 6464
rect -302 5888 -296 6464
rect 4479 6444 4681 6464
rect 4479 6410 4491 6444
rect 4525 6410 4563 6444
rect 4597 6410 4635 6444
rect 4669 6410 4681 6444
rect 4479 6398 4681 6410
rect 13679 6444 13881 6464
rect 13679 6410 13691 6444
rect 13725 6410 13763 6444
rect 13797 6410 13835 6444
rect 13869 6410 13881 6444
rect 13679 6398 13881 6410
rect 22879 6444 23081 6464
rect 22879 6410 22891 6444
rect 22925 6410 22963 6444
rect 22997 6410 23035 6444
rect 23069 6410 23081 6444
rect 22879 6398 23081 6410
rect 32079 6444 32281 6464
rect 32079 6410 32091 6444
rect 32125 6410 32163 6444
rect 32197 6410 32235 6444
rect 32269 6410 32281 6444
rect 32079 6398 32281 6410
rect 41279 6444 41481 6464
rect 41279 6410 41291 6444
rect 41325 6410 41363 6444
rect 41397 6410 41435 6444
rect 41469 6410 41481 6444
rect 41279 6398 41481 6410
rect 50479 6444 50681 6464
rect 50479 6410 50491 6444
rect 50525 6410 50563 6444
rect 50597 6410 50635 6444
rect 50669 6410 50681 6444
rect 50479 6398 50681 6410
rect 59679 6444 59881 6464
rect 59679 6410 59691 6444
rect 59725 6410 59763 6444
rect 59797 6410 59835 6444
rect 59869 6410 59881 6444
rect 59679 6398 59881 6410
rect 68879 6444 69081 6464
rect 68879 6410 68891 6444
rect 68925 6410 68963 6444
rect 68997 6410 69035 6444
rect 69069 6410 69081 6444
rect 68879 6398 69081 6410
rect 4166 5966 4176 6398
rect 4246 5966 4256 6398
rect 4354 6332 4412 6360
rect 4354 6298 4366 6332
rect 4400 6298 4412 6332
rect 4354 6260 4412 6298
rect 4354 6226 4366 6260
rect 4400 6226 4412 6260
rect 4354 6188 4412 6226
rect 4354 6154 4366 6188
rect 4400 6154 4412 6188
rect 4354 6116 4412 6154
rect 4354 6082 4366 6116
rect 4400 6082 4412 6116
rect 4354 6054 4412 6082
rect 4468 6332 4520 6360
rect 4468 6298 4477 6332
rect 4511 6298 4520 6332
rect 4468 6260 4520 6298
rect 4468 6226 4477 6260
rect 4511 6226 4520 6260
rect 4468 6188 4520 6226
rect 4468 6176 4477 6188
rect 4511 6176 4520 6188
rect 4468 6116 4520 6124
rect 4468 6112 4477 6116
rect 4511 6112 4520 6116
rect 4468 6054 4520 6060
rect 4554 6354 4606 6360
rect 4554 6298 4563 6302
rect 4597 6298 4606 6302
rect 4554 6290 4606 6298
rect 4554 6226 4563 6238
rect 4597 6226 4606 6238
rect 4554 6188 4606 6226
rect 4554 6154 4563 6188
rect 4597 6154 4606 6188
rect 4554 6116 4606 6154
rect 4554 6082 4563 6116
rect 4597 6082 4606 6116
rect 4554 6054 4606 6082
rect 4640 6332 4692 6360
rect 4640 6298 4649 6332
rect 4683 6298 4692 6332
rect 4640 6260 4692 6298
rect 4640 6226 4649 6260
rect 4683 6226 4692 6260
rect 4640 6188 4692 6226
rect 4640 6176 4649 6188
rect 4683 6176 4692 6188
rect 4640 6116 4692 6124
rect 4640 6112 4649 6116
rect 4683 6112 4692 6116
rect 4640 6054 4692 6060
rect 4748 6332 4806 6360
rect 4748 6298 4760 6332
rect 4794 6298 4806 6332
rect 4748 6260 4806 6298
rect 4748 6226 4760 6260
rect 4794 6226 4806 6260
rect 4748 6188 4806 6226
rect 4748 6154 4760 6188
rect 4794 6154 4806 6188
rect 4748 6116 4806 6154
rect 4748 6082 4760 6116
rect 4794 6082 4806 6116
rect 4748 6054 4806 6082
rect -342 5876 -296 5888
rect 4366 5880 4400 6054
rect 4479 6004 4681 6016
rect 4479 5970 4491 6004
rect 4525 5970 4563 6004
rect 4597 5970 4635 6004
rect 4669 5970 4681 6004
rect 4479 5950 4681 5970
rect 4479 5890 4493 5950
rect 4667 5890 4681 5950
rect -610 5800 -600 5840
rect -560 5830 -550 5840
rect -240 5830 -160 5840
rect -560 5800 -430 5830
rect -610 5790 -430 5800
rect -610 5780 -550 5790
rect -240 5770 -230 5830
rect -170 5770 -160 5830
rect -240 5760 -160 5770
rect 4360 5820 4400 5880
rect 4760 5880 4794 6054
rect 4904 5966 4914 6398
rect 4984 5966 4994 6398
rect 13366 5966 13376 6398
rect 13446 5966 13456 6398
rect 13554 6332 13612 6360
rect 13554 6298 13566 6332
rect 13600 6298 13612 6332
rect 13554 6260 13612 6298
rect 13554 6226 13566 6260
rect 13600 6226 13612 6260
rect 13554 6188 13612 6226
rect 13554 6154 13566 6188
rect 13600 6154 13612 6188
rect 13554 6116 13612 6154
rect 13554 6082 13566 6116
rect 13600 6082 13612 6116
rect 13554 6054 13612 6082
rect 13668 6332 13720 6360
rect 13668 6298 13677 6332
rect 13711 6298 13720 6332
rect 13668 6260 13720 6298
rect 13668 6226 13677 6260
rect 13711 6226 13720 6260
rect 13668 6188 13720 6226
rect 13668 6176 13677 6188
rect 13711 6176 13720 6188
rect 13668 6116 13720 6124
rect 13668 6112 13677 6116
rect 13711 6112 13720 6116
rect 13668 6054 13720 6060
rect 13754 6354 13806 6360
rect 13754 6298 13763 6302
rect 13797 6298 13806 6302
rect 13754 6290 13806 6298
rect 13754 6226 13763 6238
rect 13797 6226 13806 6238
rect 13754 6188 13806 6226
rect 13754 6154 13763 6188
rect 13797 6154 13806 6188
rect 13754 6116 13806 6154
rect 13754 6082 13763 6116
rect 13797 6082 13806 6116
rect 13754 6054 13806 6082
rect 13840 6332 13892 6360
rect 13840 6298 13849 6332
rect 13883 6298 13892 6332
rect 13840 6260 13892 6298
rect 13840 6226 13849 6260
rect 13883 6226 13892 6260
rect 13840 6188 13892 6226
rect 13840 6176 13849 6188
rect 13883 6176 13892 6188
rect 13840 6116 13892 6124
rect 13840 6112 13849 6116
rect 13883 6112 13892 6116
rect 13840 6054 13892 6060
rect 13948 6332 14006 6360
rect 13948 6298 13960 6332
rect 13994 6298 14006 6332
rect 13948 6260 14006 6298
rect 13948 6226 13960 6260
rect 13994 6226 14006 6260
rect 13948 6188 14006 6226
rect 13948 6154 13960 6188
rect 13994 6154 14006 6188
rect 13948 6116 14006 6154
rect 13948 6082 13960 6116
rect 13994 6082 14006 6116
rect 13948 6054 14006 6082
rect 13566 5880 13600 6054
rect 13679 6004 13881 6016
rect 13679 5970 13691 6004
rect 13725 5970 13763 6004
rect 13797 5970 13835 6004
rect 13869 5970 13881 6004
rect 13679 5950 13881 5970
rect 13679 5890 13693 5950
rect 13867 5890 13881 5950
rect 4760 5820 4800 5880
rect -430 5734 -384 5746
rect -430 5458 -424 5734
rect -390 5458 -384 5734
rect -430 5446 -384 5458
rect -342 5734 -296 5746
rect -342 5458 -336 5734
rect -302 5458 -296 5734
rect -342 5446 -296 5458
rect -3880 5370 0 5380
rect -3880 5320 -440 5370
rect -390 5320 -330 5370
rect -280 5320 0 5370
rect -3880 5300 0 5320
rect -3880 2990 -1870 5300
rect 4360 2990 4800 5820
rect 13560 5820 13600 5880
rect 13960 5880 13994 6054
rect 14104 5966 14114 6398
rect 14184 5966 14194 6398
rect 22566 5966 22576 6398
rect 22646 5966 22656 6398
rect 22754 6332 22812 6360
rect 22754 6298 22766 6332
rect 22800 6298 22812 6332
rect 22754 6260 22812 6298
rect 22754 6226 22766 6260
rect 22800 6226 22812 6260
rect 22754 6188 22812 6226
rect 22754 6154 22766 6188
rect 22800 6154 22812 6188
rect 22754 6116 22812 6154
rect 22754 6082 22766 6116
rect 22800 6082 22812 6116
rect 22754 6054 22812 6082
rect 22868 6332 22920 6360
rect 22868 6298 22877 6332
rect 22911 6298 22920 6332
rect 22868 6260 22920 6298
rect 22868 6226 22877 6260
rect 22911 6226 22920 6260
rect 22868 6188 22920 6226
rect 22868 6176 22877 6188
rect 22911 6176 22920 6188
rect 22868 6116 22920 6124
rect 22868 6112 22877 6116
rect 22911 6112 22920 6116
rect 22868 6054 22920 6060
rect 22954 6354 23006 6360
rect 22954 6298 22963 6302
rect 22997 6298 23006 6302
rect 22954 6290 23006 6298
rect 22954 6226 22963 6238
rect 22997 6226 23006 6238
rect 22954 6188 23006 6226
rect 22954 6154 22963 6188
rect 22997 6154 23006 6188
rect 22954 6116 23006 6154
rect 22954 6082 22963 6116
rect 22997 6082 23006 6116
rect 22954 6054 23006 6082
rect 23040 6332 23092 6360
rect 23040 6298 23049 6332
rect 23083 6298 23092 6332
rect 23040 6260 23092 6298
rect 23040 6226 23049 6260
rect 23083 6226 23092 6260
rect 23040 6188 23092 6226
rect 23040 6176 23049 6188
rect 23083 6176 23092 6188
rect 23040 6116 23092 6124
rect 23040 6112 23049 6116
rect 23083 6112 23092 6116
rect 23040 6054 23092 6060
rect 23148 6332 23206 6360
rect 23148 6298 23160 6332
rect 23194 6298 23206 6332
rect 23148 6260 23206 6298
rect 23148 6226 23160 6260
rect 23194 6226 23206 6260
rect 23148 6188 23206 6226
rect 23148 6154 23160 6188
rect 23194 6154 23206 6188
rect 23148 6116 23206 6154
rect 23148 6082 23160 6116
rect 23194 6082 23206 6116
rect 23148 6054 23206 6082
rect 22766 5880 22800 6054
rect 22879 6004 23081 6016
rect 22879 5970 22891 6004
rect 22925 5970 22963 6004
rect 22997 5970 23035 6004
rect 23069 5970 23081 6004
rect 22879 5950 23081 5970
rect 22879 5890 22893 5950
rect 23067 5890 23081 5950
rect 13960 5820 14000 5880
rect 13560 2990 14000 5820
rect 22760 5820 22800 5880
rect 23160 5880 23194 6054
rect 23304 5966 23314 6398
rect 23384 5966 23394 6398
rect 31766 5966 31776 6398
rect 31846 5966 31856 6398
rect 31954 6332 32012 6360
rect 31954 6298 31966 6332
rect 32000 6298 32012 6332
rect 31954 6260 32012 6298
rect 31954 6226 31966 6260
rect 32000 6226 32012 6260
rect 31954 6188 32012 6226
rect 31954 6154 31966 6188
rect 32000 6154 32012 6188
rect 31954 6116 32012 6154
rect 31954 6082 31966 6116
rect 32000 6082 32012 6116
rect 31954 6054 32012 6082
rect 32068 6332 32120 6360
rect 32068 6298 32077 6332
rect 32111 6298 32120 6332
rect 32068 6260 32120 6298
rect 32068 6226 32077 6260
rect 32111 6226 32120 6260
rect 32068 6188 32120 6226
rect 32068 6176 32077 6188
rect 32111 6176 32120 6188
rect 32068 6116 32120 6124
rect 32068 6112 32077 6116
rect 32111 6112 32120 6116
rect 32068 6054 32120 6060
rect 32154 6354 32206 6360
rect 32154 6298 32163 6302
rect 32197 6298 32206 6302
rect 32154 6290 32206 6298
rect 32154 6226 32163 6238
rect 32197 6226 32206 6238
rect 32154 6188 32206 6226
rect 32154 6154 32163 6188
rect 32197 6154 32206 6188
rect 32154 6116 32206 6154
rect 32154 6082 32163 6116
rect 32197 6082 32206 6116
rect 32154 6054 32206 6082
rect 32240 6332 32292 6360
rect 32240 6298 32249 6332
rect 32283 6298 32292 6332
rect 32240 6260 32292 6298
rect 32240 6226 32249 6260
rect 32283 6226 32292 6260
rect 32240 6188 32292 6226
rect 32240 6176 32249 6188
rect 32283 6176 32292 6188
rect 32240 6116 32292 6124
rect 32240 6112 32249 6116
rect 32283 6112 32292 6116
rect 32240 6054 32292 6060
rect 32348 6332 32406 6360
rect 32348 6298 32360 6332
rect 32394 6298 32406 6332
rect 32348 6260 32406 6298
rect 32348 6226 32360 6260
rect 32394 6226 32406 6260
rect 32348 6188 32406 6226
rect 32348 6154 32360 6188
rect 32394 6154 32406 6188
rect 32348 6116 32406 6154
rect 32348 6082 32360 6116
rect 32394 6082 32406 6116
rect 32348 6054 32406 6082
rect 31966 5880 32000 6054
rect 32079 6004 32281 6016
rect 32079 5970 32091 6004
rect 32125 5970 32163 6004
rect 32197 5970 32235 6004
rect 32269 5970 32281 6004
rect 32079 5950 32281 5970
rect 32079 5890 32093 5950
rect 32267 5890 32281 5950
rect 23160 5820 23200 5880
rect 22760 2990 23200 5820
rect 31960 5820 32000 5880
rect 32360 5880 32394 6054
rect 32504 5966 32514 6398
rect 32584 5966 32594 6398
rect 40966 5966 40976 6398
rect 41046 5966 41056 6398
rect 41154 6332 41212 6360
rect 41154 6298 41166 6332
rect 41200 6298 41212 6332
rect 41154 6260 41212 6298
rect 41154 6226 41166 6260
rect 41200 6226 41212 6260
rect 41154 6188 41212 6226
rect 41154 6154 41166 6188
rect 41200 6154 41212 6188
rect 41154 6116 41212 6154
rect 41154 6082 41166 6116
rect 41200 6082 41212 6116
rect 41154 6054 41212 6082
rect 41268 6332 41320 6360
rect 41268 6298 41277 6332
rect 41311 6298 41320 6332
rect 41268 6260 41320 6298
rect 41268 6226 41277 6260
rect 41311 6226 41320 6260
rect 41268 6188 41320 6226
rect 41268 6176 41277 6188
rect 41311 6176 41320 6188
rect 41268 6116 41320 6124
rect 41268 6112 41277 6116
rect 41311 6112 41320 6116
rect 41268 6054 41320 6060
rect 41354 6354 41406 6360
rect 41354 6298 41363 6302
rect 41397 6298 41406 6302
rect 41354 6290 41406 6298
rect 41354 6226 41363 6238
rect 41397 6226 41406 6238
rect 41354 6188 41406 6226
rect 41354 6154 41363 6188
rect 41397 6154 41406 6188
rect 41354 6116 41406 6154
rect 41354 6082 41363 6116
rect 41397 6082 41406 6116
rect 41354 6054 41406 6082
rect 41440 6332 41492 6360
rect 41440 6298 41449 6332
rect 41483 6298 41492 6332
rect 41440 6260 41492 6298
rect 41440 6226 41449 6260
rect 41483 6226 41492 6260
rect 41440 6188 41492 6226
rect 41440 6176 41449 6188
rect 41483 6176 41492 6188
rect 41440 6116 41492 6124
rect 41440 6112 41449 6116
rect 41483 6112 41492 6116
rect 41440 6054 41492 6060
rect 41548 6332 41606 6360
rect 41548 6298 41560 6332
rect 41594 6298 41606 6332
rect 41548 6260 41606 6298
rect 41548 6226 41560 6260
rect 41594 6226 41606 6260
rect 41548 6188 41606 6226
rect 41548 6154 41560 6188
rect 41594 6154 41606 6188
rect 41548 6116 41606 6154
rect 41548 6082 41560 6116
rect 41594 6082 41606 6116
rect 41548 6054 41606 6082
rect 41166 5880 41200 6054
rect 41279 6004 41481 6016
rect 41279 5970 41291 6004
rect 41325 5970 41363 6004
rect 41397 5970 41435 6004
rect 41469 5970 41481 6004
rect 41279 5950 41481 5970
rect 41279 5890 41293 5950
rect 41467 5890 41481 5950
rect 32360 5820 32400 5880
rect 31960 2990 32400 5820
rect 41160 5820 41200 5880
rect 41560 5880 41594 6054
rect 41704 5966 41714 6398
rect 41784 5966 41794 6398
rect 50166 5966 50176 6398
rect 50246 5966 50256 6398
rect 50354 6332 50412 6360
rect 50354 6298 50366 6332
rect 50400 6298 50412 6332
rect 50354 6260 50412 6298
rect 50354 6226 50366 6260
rect 50400 6226 50412 6260
rect 50354 6188 50412 6226
rect 50354 6154 50366 6188
rect 50400 6154 50412 6188
rect 50354 6116 50412 6154
rect 50354 6082 50366 6116
rect 50400 6082 50412 6116
rect 50354 6054 50412 6082
rect 50468 6332 50520 6360
rect 50468 6298 50477 6332
rect 50511 6298 50520 6332
rect 50468 6260 50520 6298
rect 50468 6226 50477 6260
rect 50511 6226 50520 6260
rect 50468 6188 50520 6226
rect 50468 6176 50477 6188
rect 50511 6176 50520 6188
rect 50468 6116 50520 6124
rect 50468 6112 50477 6116
rect 50511 6112 50520 6116
rect 50468 6054 50520 6060
rect 50554 6354 50606 6360
rect 50554 6298 50563 6302
rect 50597 6298 50606 6302
rect 50554 6290 50606 6298
rect 50554 6226 50563 6238
rect 50597 6226 50606 6238
rect 50554 6188 50606 6226
rect 50554 6154 50563 6188
rect 50597 6154 50606 6188
rect 50554 6116 50606 6154
rect 50554 6082 50563 6116
rect 50597 6082 50606 6116
rect 50554 6054 50606 6082
rect 50640 6332 50692 6360
rect 50640 6298 50649 6332
rect 50683 6298 50692 6332
rect 50640 6260 50692 6298
rect 50640 6226 50649 6260
rect 50683 6226 50692 6260
rect 50640 6188 50692 6226
rect 50640 6176 50649 6188
rect 50683 6176 50692 6188
rect 50640 6116 50692 6124
rect 50640 6112 50649 6116
rect 50683 6112 50692 6116
rect 50640 6054 50692 6060
rect 50748 6332 50806 6360
rect 50748 6298 50760 6332
rect 50794 6298 50806 6332
rect 50748 6260 50806 6298
rect 50748 6226 50760 6260
rect 50794 6226 50806 6260
rect 50748 6188 50806 6226
rect 50748 6154 50760 6188
rect 50794 6154 50806 6188
rect 50748 6116 50806 6154
rect 50748 6082 50760 6116
rect 50794 6082 50806 6116
rect 50748 6054 50806 6082
rect 50366 5880 50400 6054
rect 50479 6004 50681 6016
rect 50479 5970 50491 6004
rect 50525 5970 50563 6004
rect 50597 5970 50635 6004
rect 50669 5970 50681 6004
rect 50479 5950 50681 5970
rect 50479 5890 50493 5950
rect 50667 5890 50681 5950
rect 41560 5820 41600 5880
rect 41160 2990 41600 5820
rect 50360 5820 50400 5880
rect 50760 5880 50794 6054
rect 50904 5966 50914 6398
rect 50984 5966 50994 6398
rect 59366 5966 59376 6398
rect 59446 5966 59456 6398
rect 59554 6332 59612 6360
rect 59554 6298 59566 6332
rect 59600 6298 59612 6332
rect 59554 6260 59612 6298
rect 59554 6226 59566 6260
rect 59600 6226 59612 6260
rect 59554 6188 59612 6226
rect 59554 6154 59566 6188
rect 59600 6154 59612 6188
rect 59554 6116 59612 6154
rect 59554 6082 59566 6116
rect 59600 6082 59612 6116
rect 59554 6054 59612 6082
rect 59668 6332 59720 6360
rect 59668 6298 59677 6332
rect 59711 6298 59720 6332
rect 59668 6260 59720 6298
rect 59668 6226 59677 6260
rect 59711 6226 59720 6260
rect 59668 6188 59720 6226
rect 59668 6176 59677 6188
rect 59711 6176 59720 6188
rect 59668 6116 59720 6124
rect 59668 6112 59677 6116
rect 59711 6112 59720 6116
rect 59668 6054 59720 6060
rect 59754 6354 59806 6360
rect 59754 6298 59763 6302
rect 59797 6298 59806 6302
rect 59754 6290 59806 6298
rect 59754 6226 59763 6238
rect 59797 6226 59806 6238
rect 59754 6188 59806 6226
rect 59754 6154 59763 6188
rect 59797 6154 59806 6188
rect 59754 6116 59806 6154
rect 59754 6082 59763 6116
rect 59797 6082 59806 6116
rect 59754 6054 59806 6082
rect 59840 6332 59892 6360
rect 59840 6298 59849 6332
rect 59883 6298 59892 6332
rect 59840 6260 59892 6298
rect 59840 6226 59849 6260
rect 59883 6226 59892 6260
rect 59840 6188 59892 6226
rect 59840 6176 59849 6188
rect 59883 6176 59892 6188
rect 59840 6116 59892 6124
rect 59840 6112 59849 6116
rect 59883 6112 59892 6116
rect 59840 6054 59892 6060
rect 59948 6332 60006 6360
rect 59948 6298 59960 6332
rect 59994 6298 60006 6332
rect 59948 6260 60006 6298
rect 59948 6226 59960 6260
rect 59994 6226 60006 6260
rect 59948 6188 60006 6226
rect 59948 6154 59960 6188
rect 59994 6154 60006 6188
rect 59948 6116 60006 6154
rect 59948 6082 59960 6116
rect 59994 6082 60006 6116
rect 59948 6054 60006 6082
rect 59566 5880 59600 6054
rect 59679 6004 59881 6016
rect 59679 5970 59691 6004
rect 59725 5970 59763 6004
rect 59797 5970 59835 6004
rect 59869 5970 59881 6004
rect 59679 5950 59881 5970
rect 59679 5890 59693 5950
rect 59867 5890 59881 5950
rect 50760 5820 50800 5880
rect 50360 2990 50800 5820
rect 59560 5820 59600 5880
rect 59960 5880 59994 6054
rect 60104 5966 60114 6398
rect 60184 5966 60194 6398
rect 68566 5966 68576 6398
rect 68646 5966 68656 6398
rect 68754 6332 68812 6360
rect 68754 6298 68766 6332
rect 68800 6298 68812 6332
rect 68754 6260 68812 6298
rect 68754 6226 68766 6260
rect 68800 6226 68812 6260
rect 68754 6188 68812 6226
rect 68754 6154 68766 6188
rect 68800 6154 68812 6188
rect 68754 6116 68812 6154
rect 68754 6082 68766 6116
rect 68800 6082 68812 6116
rect 68754 6054 68812 6082
rect 68868 6332 68920 6360
rect 68868 6298 68877 6332
rect 68911 6298 68920 6332
rect 68868 6260 68920 6298
rect 68868 6226 68877 6260
rect 68911 6226 68920 6260
rect 68868 6188 68920 6226
rect 68868 6176 68877 6188
rect 68911 6176 68920 6188
rect 68868 6116 68920 6124
rect 68868 6112 68877 6116
rect 68911 6112 68920 6116
rect 68868 6054 68920 6060
rect 68954 6354 69006 6360
rect 68954 6298 68963 6302
rect 68997 6298 69006 6302
rect 68954 6290 69006 6298
rect 68954 6226 68963 6238
rect 68997 6226 69006 6238
rect 68954 6188 69006 6226
rect 68954 6154 68963 6188
rect 68997 6154 69006 6188
rect 68954 6116 69006 6154
rect 68954 6082 68963 6116
rect 68997 6082 69006 6116
rect 68954 6054 69006 6082
rect 69040 6332 69092 6360
rect 69040 6298 69049 6332
rect 69083 6298 69092 6332
rect 69040 6260 69092 6298
rect 69040 6226 69049 6260
rect 69083 6226 69092 6260
rect 69040 6188 69092 6226
rect 69040 6176 69049 6188
rect 69083 6176 69092 6188
rect 69040 6116 69092 6124
rect 69040 6112 69049 6116
rect 69083 6112 69092 6116
rect 69040 6054 69092 6060
rect 69148 6332 69206 6360
rect 69148 6298 69160 6332
rect 69194 6298 69206 6332
rect 69148 6260 69206 6298
rect 69148 6226 69160 6260
rect 69194 6226 69206 6260
rect 69148 6188 69206 6226
rect 69148 6154 69160 6188
rect 69194 6154 69206 6188
rect 69148 6116 69206 6154
rect 69148 6082 69160 6116
rect 69194 6082 69206 6116
rect 69148 6054 69206 6082
rect 68766 5880 68800 6054
rect 68879 6004 69081 6016
rect 68879 5970 68891 6004
rect 68925 5970 68963 6004
rect 68997 5970 69035 6004
rect 69069 5970 69081 6004
rect 68879 5950 69081 5970
rect 68879 5890 68893 5950
rect 69067 5890 69081 5950
rect 59960 5820 60000 5880
rect 59560 2990 60000 5820
rect 68760 5820 68800 5880
rect 69160 5880 69194 6054
rect 69304 5966 69314 6398
rect 69384 5966 69394 6398
rect 69160 5820 69200 5880
rect 68760 2990 69200 5820
rect -3880 990 73600 2990
rect -3880 -10 -1870 990
<< via1 >>
rect -490 95530 -240 95540
rect -490 95490 -480 95530
rect -480 95490 -440 95530
rect -440 95490 -400 95530
rect -400 95490 -360 95530
rect -360 95490 -310 95530
rect -310 95490 -270 95530
rect -270 95490 -240 95530
rect -490 95480 -240 95490
rect 4176 95301 4246 95318
rect 4176 94904 4192 95301
rect 4192 94904 4230 95301
rect 4230 94904 4246 95301
rect 4176 94886 4246 94904
rect 4468 95074 4477 95096
rect 4477 95074 4511 95096
rect 4511 95074 4520 95096
rect 4468 95044 4520 95074
rect 4468 95002 4477 95032
rect 4477 95002 4511 95032
rect 4511 95002 4520 95032
rect 4468 94980 4520 95002
rect 4554 95252 4606 95274
rect 4554 95222 4563 95252
rect 4563 95222 4597 95252
rect 4597 95222 4606 95252
rect 4554 95180 4606 95210
rect 4554 95158 4563 95180
rect 4563 95158 4597 95180
rect 4597 95158 4606 95180
rect 4640 95074 4649 95096
rect 4649 95074 4683 95096
rect 4683 95074 4692 95096
rect 4640 95044 4692 95074
rect 4640 95002 4649 95032
rect 4649 95002 4683 95032
rect 4683 95002 4692 95032
rect 4640 94980 4692 95002
rect 4493 94810 4667 94870
rect -230 94740 -170 94750
rect -230 94700 -220 94740
rect -220 94700 -180 94740
rect -180 94700 -170 94740
rect -230 94690 -170 94700
rect 4914 95301 4984 95318
rect 4914 94904 4930 95301
rect 4930 94904 4968 95301
rect 4968 94904 4984 95301
rect 4914 94886 4984 94904
rect -490 85650 -240 85660
rect -490 85610 -480 85650
rect -480 85610 -440 85650
rect -440 85610 -400 85650
rect -400 85610 -360 85650
rect -360 85610 -310 85650
rect -310 85610 -270 85650
rect -270 85610 -240 85650
rect -490 85600 -240 85610
rect 4176 85421 4246 85438
rect 4176 85024 4192 85421
rect 4192 85024 4230 85421
rect 4230 85024 4246 85421
rect 4176 85006 4246 85024
rect 4468 85194 4477 85216
rect 4477 85194 4511 85216
rect 4511 85194 4520 85216
rect 4468 85164 4520 85194
rect 4468 85122 4477 85152
rect 4477 85122 4511 85152
rect 4511 85122 4520 85152
rect 4468 85100 4520 85122
rect 4554 85372 4606 85394
rect 4554 85342 4563 85372
rect 4563 85342 4597 85372
rect 4597 85342 4606 85372
rect 4554 85300 4606 85330
rect 4554 85278 4563 85300
rect 4563 85278 4597 85300
rect 4597 85278 4606 85300
rect 4640 85194 4649 85216
rect 4649 85194 4683 85216
rect 4683 85194 4692 85216
rect 4640 85164 4692 85194
rect 4640 85122 4649 85152
rect 4649 85122 4683 85152
rect 4683 85122 4692 85152
rect 4640 85100 4692 85122
rect 4493 84930 4667 84990
rect -230 84860 -170 84870
rect -230 84820 -220 84860
rect -220 84820 -180 84860
rect -180 84820 -170 84860
rect -230 84810 -170 84820
rect 4914 85421 4984 85438
rect 4914 85024 4930 85421
rect 4930 85024 4968 85421
rect 4968 85024 4984 85421
rect 4914 85006 4984 85024
rect 13376 85421 13446 85438
rect 13376 85024 13392 85421
rect 13392 85024 13430 85421
rect 13430 85024 13446 85421
rect 13376 85006 13446 85024
rect 13668 85194 13677 85216
rect 13677 85194 13711 85216
rect 13711 85194 13720 85216
rect 13668 85164 13720 85194
rect 13668 85122 13677 85152
rect 13677 85122 13711 85152
rect 13711 85122 13720 85152
rect 13668 85100 13720 85122
rect 13754 85372 13806 85394
rect 13754 85342 13763 85372
rect 13763 85342 13797 85372
rect 13797 85342 13806 85372
rect 13754 85300 13806 85330
rect 13754 85278 13763 85300
rect 13763 85278 13797 85300
rect 13797 85278 13806 85300
rect 13840 85194 13849 85216
rect 13849 85194 13883 85216
rect 13883 85194 13892 85216
rect 13840 85164 13892 85194
rect 13840 85122 13849 85152
rect 13849 85122 13883 85152
rect 13883 85122 13892 85152
rect 13840 85100 13892 85122
rect 13693 84930 13867 84990
rect 14114 85421 14184 85438
rect 14114 85024 14130 85421
rect 14130 85024 14168 85421
rect 14168 85024 14184 85421
rect 14114 85006 14184 85024
rect -490 75770 -240 75780
rect -490 75730 -480 75770
rect -480 75730 -440 75770
rect -440 75730 -400 75770
rect -400 75730 -360 75770
rect -360 75730 -310 75770
rect -310 75730 -270 75770
rect -270 75730 -240 75770
rect -490 75720 -240 75730
rect 4176 75541 4246 75558
rect 4176 75144 4192 75541
rect 4192 75144 4230 75541
rect 4230 75144 4246 75541
rect 4176 75126 4246 75144
rect 4468 75314 4477 75336
rect 4477 75314 4511 75336
rect 4511 75314 4520 75336
rect 4468 75284 4520 75314
rect 4468 75242 4477 75272
rect 4477 75242 4511 75272
rect 4511 75242 4520 75272
rect 4468 75220 4520 75242
rect 4554 75492 4606 75514
rect 4554 75462 4563 75492
rect 4563 75462 4597 75492
rect 4597 75462 4606 75492
rect 4554 75420 4606 75450
rect 4554 75398 4563 75420
rect 4563 75398 4597 75420
rect 4597 75398 4606 75420
rect 4640 75314 4649 75336
rect 4649 75314 4683 75336
rect 4683 75314 4692 75336
rect 4640 75284 4692 75314
rect 4640 75242 4649 75272
rect 4649 75242 4683 75272
rect 4683 75242 4692 75272
rect 4640 75220 4692 75242
rect 4493 75050 4667 75110
rect -230 74980 -170 74990
rect -230 74940 -220 74980
rect -220 74940 -180 74980
rect -180 74940 -170 74980
rect -230 74930 -170 74940
rect 4914 75541 4984 75558
rect 4914 75144 4930 75541
rect 4930 75144 4968 75541
rect 4968 75144 4984 75541
rect 4914 75126 4984 75144
rect 13376 75541 13446 75558
rect 13376 75144 13392 75541
rect 13392 75144 13430 75541
rect 13430 75144 13446 75541
rect 13376 75126 13446 75144
rect 13668 75314 13677 75336
rect 13677 75314 13711 75336
rect 13711 75314 13720 75336
rect 13668 75284 13720 75314
rect 13668 75242 13677 75272
rect 13677 75242 13711 75272
rect 13711 75242 13720 75272
rect 13668 75220 13720 75242
rect 13754 75492 13806 75514
rect 13754 75462 13763 75492
rect 13763 75462 13797 75492
rect 13797 75462 13806 75492
rect 13754 75420 13806 75450
rect 13754 75398 13763 75420
rect 13763 75398 13797 75420
rect 13797 75398 13806 75420
rect 13840 75314 13849 75336
rect 13849 75314 13883 75336
rect 13883 75314 13892 75336
rect 13840 75284 13892 75314
rect 13840 75242 13849 75272
rect 13849 75242 13883 75272
rect 13883 75242 13892 75272
rect 13840 75220 13892 75242
rect 13693 75050 13867 75110
rect 14114 75541 14184 75558
rect 14114 75144 14130 75541
rect 14130 75144 14168 75541
rect 14168 75144 14184 75541
rect 14114 75126 14184 75144
rect 22576 75541 22646 75558
rect 22576 75144 22592 75541
rect 22592 75144 22630 75541
rect 22630 75144 22646 75541
rect 22576 75126 22646 75144
rect 22868 75314 22877 75336
rect 22877 75314 22911 75336
rect 22911 75314 22920 75336
rect 22868 75284 22920 75314
rect 22868 75242 22877 75272
rect 22877 75242 22911 75272
rect 22911 75242 22920 75272
rect 22868 75220 22920 75242
rect 22954 75492 23006 75514
rect 22954 75462 22963 75492
rect 22963 75462 22997 75492
rect 22997 75462 23006 75492
rect 22954 75420 23006 75450
rect 22954 75398 22963 75420
rect 22963 75398 22997 75420
rect 22997 75398 23006 75420
rect 23040 75314 23049 75336
rect 23049 75314 23083 75336
rect 23083 75314 23092 75336
rect 23040 75284 23092 75314
rect 23040 75242 23049 75272
rect 23049 75242 23083 75272
rect 23083 75242 23092 75272
rect 23040 75220 23092 75242
rect 22893 75050 23067 75110
rect 23314 75541 23384 75558
rect 23314 75144 23330 75541
rect 23330 75144 23368 75541
rect 23368 75144 23384 75541
rect 23314 75126 23384 75144
rect 31776 75541 31846 75558
rect 31776 75144 31792 75541
rect 31792 75144 31830 75541
rect 31830 75144 31846 75541
rect 31776 75126 31846 75144
rect 32068 75314 32077 75336
rect 32077 75314 32111 75336
rect 32111 75314 32120 75336
rect 32068 75284 32120 75314
rect 32068 75242 32077 75272
rect 32077 75242 32111 75272
rect 32111 75242 32120 75272
rect 32068 75220 32120 75242
rect 32154 75492 32206 75514
rect 32154 75462 32163 75492
rect 32163 75462 32197 75492
rect 32197 75462 32206 75492
rect 32154 75420 32206 75450
rect 32154 75398 32163 75420
rect 32163 75398 32197 75420
rect 32197 75398 32206 75420
rect 32240 75314 32249 75336
rect 32249 75314 32283 75336
rect 32283 75314 32292 75336
rect 32240 75284 32292 75314
rect 32240 75242 32249 75272
rect 32249 75242 32283 75272
rect 32283 75242 32292 75272
rect 32240 75220 32292 75242
rect 32093 75050 32267 75110
rect 32514 75541 32584 75558
rect 32514 75144 32530 75541
rect 32530 75144 32568 75541
rect 32568 75144 32584 75541
rect 32514 75126 32584 75144
rect -490 65890 -240 65900
rect -490 65850 -480 65890
rect -480 65850 -440 65890
rect -440 65850 -400 65890
rect -400 65850 -360 65890
rect -360 65850 -310 65890
rect -310 65850 -270 65890
rect -270 65850 -240 65890
rect -490 65840 -240 65850
rect 4176 65661 4246 65678
rect 4176 65264 4192 65661
rect 4192 65264 4230 65661
rect 4230 65264 4246 65661
rect 4176 65246 4246 65264
rect 4468 65434 4477 65456
rect 4477 65434 4511 65456
rect 4511 65434 4520 65456
rect 4468 65404 4520 65434
rect 4468 65362 4477 65392
rect 4477 65362 4511 65392
rect 4511 65362 4520 65392
rect 4468 65340 4520 65362
rect 4554 65612 4606 65634
rect 4554 65582 4563 65612
rect 4563 65582 4597 65612
rect 4597 65582 4606 65612
rect 4554 65540 4606 65570
rect 4554 65518 4563 65540
rect 4563 65518 4597 65540
rect 4597 65518 4606 65540
rect 4640 65434 4649 65456
rect 4649 65434 4683 65456
rect 4683 65434 4692 65456
rect 4640 65404 4692 65434
rect 4640 65362 4649 65392
rect 4649 65362 4683 65392
rect 4683 65362 4692 65392
rect 4640 65340 4692 65362
rect 4493 65170 4667 65230
rect -230 65100 -170 65110
rect -230 65060 -220 65100
rect -220 65060 -180 65100
rect -180 65060 -170 65100
rect -230 65050 -170 65060
rect 4914 65661 4984 65678
rect 4914 65264 4930 65661
rect 4930 65264 4968 65661
rect 4968 65264 4984 65661
rect 4914 65246 4984 65264
rect 13376 65661 13446 65678
rect 13376 65264 13392 65661
rect 13392 65264 13430 65661
rect 13430 65264 13446 65661
rect 13376 65246 13446 65264
rect 13668 65434 13677 65456
rect 13677 65434 13711 65456
rect 13711 65434 13720 65456
rect 13668 65404 13720 65434
rect 13668 65362 13677 65392
rect 13677 65362 13711 65392
rect 13711 65362 13720 65392
rect 13668 65340 13720 65362
rect 13754 65612 13806 65634
rect 13754 65582 13763 65612
rect 13763 65582 13797 65612
rect 13797 65582 13806 65612
rect 13754 65540 13806 65570
rect 13754 65518 13763 65540
rect 13763 65518 13797 65540
rect 13797 65518 13806 65540
rect 13840 65434 13849 65456
rect 13849 65434 13883 65456
rect 13883 65434 13892 65456
rect 13840 65404 13892 65434
rect 13840 65362 13849 65392
rect 13849 65362 13883 65392
rect 13883 65362 13892 65392
rect 13840 65340 13892 65362
rect 13693 65170 13867 65230
rect 14114 65661 14184 65678
rect 14114 65264 14130 65661
rect 14130 65264 14168 65661
rect 14168 65264 14184 65661
rect 14114 65246 14184 65264
rect 22576 65661 22646 65678
rect 22576 65264 22592 65661
rect 22592 65264 22630 65661
rect 22630 65264 22646 65661
rect 22576 65246 22646 65264
rect 22868 65434 22877 65456
rect 22877 65434 22911 65456
rect 22911 65434 22920 65456
rect 22868 65404 22920 65434
rect 22868 65362 22877 65392
rect 22877 65362 22911 65392
rect 22911 65362 22920 65392
rect 22868 65340 22920 65362
rect 22954 65612 23006 65634
rect 22954 65582 22963 65612
rect 22963 65582 22997 65612
rect 22997 65582 23006 65612
rect 22954 65540 23006 65570
rect 22954 65518 22963 65540
rect 22963 65518 22997 65540
rect 22997 65518 23006 65540
rect 23040 65434 23049 65456
rect 23049 65434 23083 65456
rect 23083 65434 23092 65456
rect 23040 65404 23092 65434
rect 23040 65362 23049 65392
rect 23049 65362 23083 65392
rect 23083 65362 23092 65392
rect 23040 65340 23092 65362
rect 22893 65170 23067 65230
rect 23314 65661 23384 65678
rect 23314 65264 23330 65661
rect 23330 65264 23368 65661
rect 23368 65264 23384 65661
rect 23314 65246 23384 65264
rect 31776 65661 31846 65678
rect 31776 65264 31792 65661
rect 31792 65264 31830 65661
rect 31830 65264 31846 65661
rect 31776 65246 31846 65264
rect 32068 65434 32077 65456
rect 32077 65434 32111 65456
rect 32111 65434 32120 65456
rect 32068 65404 32120 65434
rect 32068 65362 32077 65392
rect 32077 65362 32111 65392
rect 32111 65362 32120 65392
rect 32068 65340 32120 65362
rect 32154 65612 32206 65634
rect 32154 65582 32163 65612
rect 32163 65582 32197 65612
rect 32197 65582 32206 65612
rect 32154 65540 32206 65570
rect 32154 65518 32163 65540
rect 32163 65518 32197 65540
rect 32197 65518 32206 65540
rect 32240 65434 32249 65456
rect 32249 65434 32283 65456
rect 32283 65434 32292 65456
rect 32240 65404 32292 65434
rect 32240 65362 32249 65392
rect 32249 65362 32283 65392
rect 32283 65362 32292 65392
rect 32240 65340 32292 65362
rect 32093 65170 32267 65230
rect 32514 65661 32584 65678
rect 32514 65264 32530 65661
rect 32530 65264 32568 65661
rect 32568 65264 32584 65661
rect 32514 65246 32584 65264
rect 40976 65661 41046 65678
rect 40976 65264 40992 65661
rect 40992 65264 41030 65661
rect 41030 65264 41046 65661
rect 40976 65246 41046 65264
rect 41268 65434 41277 65456
rect 41277 65434 41311 65456
rect 41311 65434 41320 65456
rect 41268 65404 41320 65434
rect 41268 65362 41277 65392
rect 41277 65362 41311 65392
rect 41311 65362 41320 65392
rect 41268 65340 41320 65362
rect 41354 65612 41406 65634
rect 41354 65582 41363 65612
rect 41363 65582 41397 65612
rect 41397 65582 41406 65612
rect 41354 65540 41406 65570
rect 41354 65518 41363 65540
rect 41363 65518 41397 65540
rect 41397 65518 41406 65540
rect 41440 65434 41449 65456
rect 41449 65434 41483 65456
rect 41483 65434 41492 65456
rect 41440 65404 41492 65434
rect 41440 65362 41449 65392
rect 41449 65362 41483 65392
rect 41483 65362 41492 65392
rect 41440 65340 41492 65362
rect 41293 65170 41467 65230
rect 41714 65661 41784 65678
rect 41714 65264 41730 65661
rect 41730 65264 41768 65661
rect 41768 65264 41784 65661
rect 41714 65246 41784 65264
rect 50176 65661 50246 65678
rect 50176 65264 50192 65661
rect 50192 65264 50230 65661
rect 50230 65264 50246 65661
rect 50176 65246 50246 65264
rect 50468 65434 50477 65456
rect 50477 65434 50511 65456
rect 50511 65434 50520 65456
rect 50468 65404 50520 65434
rect 50468 65362 50477 65392
rect 50477 65362 50511 65392
rect 50511 65362 50520 65392
rect 50468 65340 50520 65362
rect 50554 65612 50606 65634
rect 50554 65582 50563 65612
rect 50563 65582 50597 65612
rect 50597 65582 50606 65612
rect 50554 65540 50606 65570
rect 50554 65518 50563 65540
rect 50563 65518 50597 65540
rect 50597 65518 50606 65540
rect 50640 65434 50649 65456
rect 50649 65434 50683 65456
rect 50683 65434 50692 65456
rect 50640 65404 50692 65434
rect 50640 65362 50649 65392
rect 50649 65362 50683 65392
rect 50683 65362 50692 65392
rect 50640 65340 50692 65362
rect 50493 65170 50667 65230
rect 50914 65661 50984 65678
rect 50914 65264 50930 65661
rect 50930 65264 50968 65661
rect 50968 65264 50984 65661
rect 50914 65246 50984 65264
rect 59376 65661 59446 65678
rect 59376 65264 59392 65661
rect 59392 65264 59430 65661
rect 59430 65264 59446 65661
rect 59376 65246 59446 65264
rect 59668 65434 59677 65456
rect 59677 65434 59711 65456
rect 59711 65434 59720 65456
rect 59668 65404 59720 65434
rect 59668 65362 59677 65392
rect 59677 65362 59711 65392
rect 59711 65362 59720 65392
rect 59668 65340 59720 65362
rect 59754 65612 59806 65634
rect 59754 65582 59763 65612
rect 59763 65582 59797 65612
rect 59797 65582 59806 65612
rect 59754 65540 59806 65570
rect 59754 65518 59763 65540
rect 59763 65518 59797 65540
rect 59797 65518 59806 65540
rect 59840 65434 59849 65456
rect 59849 65434 59883 65456
rect 59883 65434 59892 65456
rect 59840 65404 59892 65434
rect 59840 65362 59849 65392
rect 59849 65362 59883 65392
rect 59883 65362 59892 65392
rect 59840 65340 59892 65362
rect 59693 65170 59867 65230
rect 60114 65661 60184 65678
rect 60114 65264 60130 65661
rect 60130 65264 60168 65661
rect 60168 65264 60184 65661
rect 60114 65246 60184 65264
rect 68576 65661 68646 65678
rect 68576 65264 68592 65661
rect 68592 65264 68630 65661
rect 68630 65264 68646 65661
rect 68576 65246 68646 65264
rect 68868 65434 68877 65456
rect 68877 65434 68911 65456
rect 68911 65434 68920 65456
rect 68868 65404 68920 65434
rect 68868 65362 68877 65392
rect 68877 65362 68911 65392
rect 68911 65362 68920 65392
rect 68868 65340 68920 65362
rect 68954 65612 69006 65634
rect 68954 65582 68963 65612
rect 68963 65582 68997 65612
rect 68997 65582 69006 65612
rect 68954 65540 69006 65570
rect 68954 65518 68963 65540
rect 68963 65518 68997 65540
rect 68997 65518 69006 65540
rect 69040 65434 69049 65456
rect 69049 65434 69083 65456
rect 69083 65434 69092 65456
rect 69040 65404 69092 65434
rect 69040 65362 69049 65392
rect 69049 65362 69083 65392
rect 69083 65362 69092 65392
rect 69040 65340 69092 65362
rect 68893 65170 69067 65230
rect 69314 65661 69384 65678
rect 69314 65264 69330 65661
rect 69330 65264 69368 65661
rect 69368 65264 69384 65661
rect 69314 65246 69384 65264
rect 4176 55781 4246 55798
rect 4176 55384 4192 55781
rect 4192 55384 4230 55781
rect 4230 55384 4246 55781
rect 4176 55366 4246 55384
rect 4468 55554 4477 55576
rect 4477 55554 4511 55576
rect 4511 55554 4520 55576
rect 4468 55524 4520 55554
rect 4468 55482 4477 55512
rect 4477 55482 4511 55512
rect 4511 55482 4520 55512
rect 4468 55460 4520 55482
rect 4554 55732 4606 55754
rect 4554 55702 4563 55732
rect 4563 55702 4597 55732
rect 4597 55702 4606 55732
rect 4554 55660 4606 55690
rect 4554 55638 4563 55660
rect 4563 55638 4597 55660
rect 4597 55638 4606 55660
rect 4640 55554 4649 55576
rect 4649 55554 4683 55576
rect 4683 55554 4692 55576
rect 4640 55524 4692 55554
rect 4640 55482 4649 55512
rect 4649 55482 4683 55512
rect 4683 55482 4692 55512
rect 4640 55460 4692 55482
rect 4493 55290 4667 55350
rect 4914 55781 4984 55798
rect 4914 55384 4930 55781
rect 4930 55384 4968 55781
rect 4968 55384 4984 55781
rect 4914 55366 4984 55384
rect 13376 55781 13446 55798
rect 13376 55384 13392 55781
rect 13392 55384 13430 55781
rect 13430 55384 13446 55781
rect 13376 55366 13446 55384
rect 13668 55554 13677 55576
rect 13677 55554 13711 55576
rect 13711 55554 13720 55576
rect 13668 55524 13720 55554
rect 13668 55482 13677 55512
rect 13677 55482 13711 55512
rect 13711 55482 13720 55512
rect 13668 55460 13720 55482
rect 13754 55732 13806 55754
rect 13754 55702 13763 55732
rect 13763 55702 13797 55732
rect 13797 55702 13806 55732
rect 13754 55660 13806 55690
rect 13754 55638 13763 55660
rect 13763 55638 13797 55660
rect 13797 55638 13806 55660
rect 13840 55554 13849 55576
rect 13849 55554 13883 55576
rect 13883 55554 13892 55576
rect 13840 55524 13892 55554
rect 13840 55482 13849 55512
rect 13849 55482 13883 55512
rect 13883 55482 13892 55512
rect 13840 55460 13892 55482
rect 13693 55290 13867 55350
rect 14114 55781 14184 55798
rect 14114 55384 14130 55781
rect 14130 55384 14168 55781
rect 14168 55384 14184 55781
rect 14114 55366 14184 55384
rect 22576 55781 22646 55798
rect 22576 55384 22592 55781
rect 22592 55384 22630 55781
rect 22630 55384 22646 55781
rect 22576 55366 22646 55384
rect 22868 55554 22877 55576
rect 22877 55554 22911 55576
rect 22911 55554 22920 55576
rect 22868 55524 22920 55554
rect 22868 55482 22877 55512
rect 22877 55482 22911 55512
rect 22911 55482 22920 55512
rect 22868 55460 22920 55482
rect 22954 55732 23006 55754
rect 22954 55702 22963 55732
rect 22963 55702 22997 55732
rect 22997 55702 23006 55732
rect 22954 55660 23006 55690
rect 22954 55638 22963 55660
rect 22963 55638 22997 55660
rect 22997 55638 23006 55660
rect 23040 55554 23049 55576
rect 23049 55554 23083 55576
rect 23083 55554 23092 55576
rect 23040 55524 23092 55554
rect 23040 55482 23049 55512
rect 23049 55482 23083 55512
rect 23083 55482 23092 55512
rect 23040 55460 23092 55482
rect 22893 55290 23067 55350
rect 23314 55781 23384 55798
rect 23314 55384 23330 55781
rect 23330 55384 23368 55781
rect 23368 55384 23384 55781
rect 23314 55366 23384 55384
rect 31776 55781 31846 55798
rect 31776 55384 31792 55781
rect 31792 55384 31830 55781
rect 31830 55384 31846 55781
rect 31776 55366 31846 55384
rect 32068 55554 32077 55576
rect 32077 55554 32111 55576
rect 32111 55554 32120 55576
rect 32068 55524 32120 55554
rect 32068 55482 32077 55512
rect 32077 55482 32111 55512
rect 32111 55482 32120 55512
rect 32068 55460 32120 55482
rect 32154 55732 32206 55754
rect 32154 55702 32163 55732
rect 32163 55702 32197 55732
rect 32197 55702 32206 55732
rect 32154 55660 32206 55690
rect 32154 55638 32163 55660
rect 32163 55638 32197 55660
rect 32197 55638 32206 55660
rect 32240 55554 32249 55576
rect 32249 55554 32283 55576
rect 32283 55554 32292 55576
rect 32240 55524 32292 55554
rect 32240 55482 32249 55512
rect 32249 55482 32283 55512
rect 32283 55482 32292 55512
rect 32240 55460 32292 55482
rect 32093 55290 32267 55350
rect 32514 55781 32584 55798
rect 32514 55384 32530 55781
rect 32530 55384 32568 55781
rect 32568 55384 32584 55781
rect 32514 55366 32584 55384
rect 40976 55781 41046 55798
rect 40976 55384 40992 55781
rect 40992 55384 41030 55781
rect 41030 55384 41046 55781
rect 40976 55366 41046 55384
rect 41268 55554 41277 55576
rect 41277 55554 41311 55576
rect 41311 55554 41320 55576
rect 41268 55524 41320 55554
rect 41268 55482 41277 55512
rect 41277 55482 41311 55512
rect 41311 55482 41320 55512
rect 41268 55460 41320 55482
rect 41354 55732 41406 55754
rect 41354 55702 41363 55732
rect 41363 55702 41397 55732
rect 41397 55702 41406 55732
rect 41354 55660 41406 55690
rect 41354 55638 41363 55660
rect 41363 55638 41397 55660
rect 41397 55638 41406 55660
rect 41440 55554 41449 55576
rect 41449 55554 41483 55576
rect 41483 55554 41492 55576
rect 41440 55524 41492 55554
rect 41440 55482 41449 55512
rect 41449 55482 41483 55512
rect 41483 55482 41492 55512
rect 41440 55460 41492 55482
rect 41293 55290 41467 55350
rect 41714 55781 41784 55798
rect 41714 55384 41730 55781
rect 41730 55384 41768 55781
rect 41768 55384 41784 55781
rect 41714 55366 41784 55384
rect 50176 55781 50246 55798
rect 50176 55384 50192 55781
rect 50192 55384 50230 55781
rect 50230 55384 50246 55781
rect 50176 55366 50246 55384
rect 50468 55554 50477 55576
rect 50477 55554 50511 55576
rect 50511 55554 50520 55576
rect 50468 55524 50520 55554
rect 50468 55482 50477 55512
rect 50477 55482 50511 55512
rect 50511 55482 50520 55512
rect 50468 55460 50520 55482
rect 50554 55732 50606 55754
rect 50554 55702 50563 55732
rect 50563 55702 50597 55732
rect 50597 55702 50606 55732
rect 50554 55660 50606 55690
rect 50554 55638 50563 55660
rect 50563 55638 50597 55660
rect 50597 55638 50606 55660
rect 50640 55554 50649 55576
rect 50649 55554 50683 55576
rect 50683 55554 50692 55576
rect 50640 55524 50692 55554
rect 50640 55482 50649 55512
rect 50649 55482 50683 55512
rect 50683 55482 50692 55512
rect 50640 55460 50692 55482
rect 50493 55290 50667 55350
rect 50914 55781 50984 55798
rect 50914 55384 50930 55781
rect 50930 55384 50968 55781
rect 50968 55384 50984 55781
rect 50914 55366 50984 55384
rect 59376 55781 59446 55798
rect 59376 55384 59392 55781
rect 59392 55384 59430 55781
rect 59430 55384 59446 55781
rect 59376 55366 59446 55384
rect 59668 55554 59677 55576
rect 59677 55554 59711 55576
rect 59711 55554 59720 55576
rect 59668 55524 59720 55554
rect 59668 55482 59677 55512
rect 59677 55482 59711 55512
rect 59711 55482 59720 55512
rect 59668 55460 59720 55482
rect 59754 55732 59806 55754
rect 59754 55702 59763 55732
rect 59763 55702 59797 55732
rect 59797 55702 59806 55732
rect 59754 55660 59806 55690
rect 59754 55638 59763 55660
rect 59763 55638 59797 55660
rect 59797 55638 59806 55660
rect 59840 55554 59849 55576
rect 59849 55554 59883 55576
rect 59883 55554 59892 55576
rect 59840 55524 59892 55554
rect 59840 55482 59849 55512
rect 59849 55482 59883 55512
rect 59883 55482 59892 55512
rect 59840 55460 59892 55482
rect 59693 55290 59867 55350
rect 60114 55781 60184 55798
rect 60114 55384 60130 55781
rect 60130 55384 60168 55781
rect 60168 55384 60184 55781
rect 60114 55366 60184 55384
rect 68576 55781 68646 55798
rect 68576 55384 68592 55781
rect 68592 55384 68630 55781
rect 68630 55384 68646 55781
rect 68576 55366 68646 55384
rect 68868 55554 68877 55576
rect 68877 55554 68911 55576
rect 68911 55554 68920 55576
rect 68868 55524 68920 55554
rect 68868 55482 68877 55512
rect 68877 55482 68911 55512
rect 68911 55482 68920 55512
rect 68868 55460 68920 55482
rect 68954 55732 69006 55754
rect 68954 55702 68963 55732
rect 68963 55702 68997 55732
rect 68997 55702 69006 55732
rect 68954 55660 69006 55690
rect 68954 55638 68963 55660
rect 68963 55638 68997 55660
rect 68997 55638 69006 55660
rect 69040 55554 69049 55576
rect 69049 55554 69083 55576
rect 69083 55554 69092 55576
rect 69040 55524 69092 55554
rect 69040 55482 69049 55512
rect 69049 55482 69083 55512
rect 69083 55482 69092 55512
rect 69040 55460 69092 55482
rect 68893 55290 69067 55350
rect 69314 55781 69384 55798
rect 69314 55384 69330 55781
rect 69330 55384 69368 55781
rect 69368 55384 69384 55781
rect 69314 55366 69384 55384
rect -490 46130 -240 46140
rect -490 46090 -480 46130
rect -480 46090 -440 46130
rect -440 46090 -400 46130
rect -400 46090 -360 46130
rect -360 46090 -310 46130
rect -310 46090 -270 46130
rect -270 46090 -240 46130
rect -490 46080 -240 46090
rect 4176 45901 4246 45918
rect 4176 45504 4192 45901
rect 4192 45504 4230 45901
rect 4230 45504 4246 45901
rect 4176 45486 4246 45504
rect 4468 45674 4477 45696
rect 4477 45674 4511 45696
rect 4511 45674 4520 45696
rect 4468 45644 4520 45674
rect 4468 45602 4477 45632
rect 4477 45602 4511 45632
rect 4511 45602 4520 45632
rect 4468 45580 4520 45602
rect 4554 45852 4606 45874
rect 4554 45822 4563 45852
rect 4563 45822 4597 45852
rect 4597 45822 4606 45852
rect 4554 45780 4606 45810
rect 4554 45758 4563 45780
rect 4563 45758 4597 45780
rect 4597 45758 4606 45780
rect 4640 45674 4649 45696
rect 4649 45674 4683 45696
rect 4683 45674 4692 45696
rect 4640 45644 4692 45674
rect 4640 45602 4649 45632
rect 4649 45602 4683 45632
rect 4683 45602 4692 45632
rect 4640 45580 4692 45602
rect 4493 45410 4667 45470
rect -230 45340 -170 45350
rect -230 45300 -220 45340
rect -220 45300 -180 45340
rect -180 45300 -170 45340
rect -230 45290 -170 45300
rect 4914 45901 4984 45918
rect 4914 45504 4930 45901
rect 4930 45504 4968 45901
rect 4968 45504 4984 45901
rect 4914 45486 4984 45504
rect 13376 45901 13446 45918
rect 13376 45504 13392 45901
rect 13392 45504 13430 45901
rect 13430 45504 13446 45901
rect 13376 45486 13446 45504
rect 13668 45674 13677 45696
rect 13677 45674 13711 45696
rect 13711 45674 13720 45696
rect 13668 45644 13720 45674
rect 13668 45602 13677 45632
rect 13677 45602 13711 45632
rect 13711 45602 13720 45632
rect 13668 45580 13720 45602
rect 13754 45852 13806 45874
rect 13754 45822 13763 45852
rect 13763 45822 13797 45852
rect 13797 45822 13806 45852
rect 13754 45780 13806 45810
rect 13754 45758 13763 45780
rect 13763 45758 13797 45780
rect 13797 45758 13806 45780
rect 13840 45674 13849 45696
rect 13849 45674 13883 45696
rect 13883 45674 13892 45696
rect 13840 45644 13892 45674
rect 13840 45602 13849 45632
rect 13849 45602 13883 45632
rect 13883 45602 13892 45632
rect 13840 45580 13892 45602
rect 13693 45410 13867 45470
rect 14114 45901 14184 45918
rect 14114 45504 14130 45901
rect 14130 45504 14168 45901
rect 14168 45504 14184 45901
rect 14114 45486 14184 45504
rect 22576 45901 22646 45918
rect 22576 45504 22592 45901
rect 22592 45504 22630 45901
rect 22630 45504 22646 45901
rect 22576 45486 22646 45504
rect 22868 45674 22877 45696
rect 22877 45674 22911 45696
rect 22911 45674 22920 45696
rect 22868 45644 22920 45674
rect 22868 45602 22877 45632
rect 22877 45602 22911 45632
rect 22911 45602 22920 45632
rect 22868 45580 22920 45602
rect 22954 45852 23006 45874
rect 22954 45822 22963 45852
rect 22963 45822 22997 45852
rect 22997 45822 23006 45852
rect 22954 45780 23006 45810
rect 22954 45758 22963 45780
rect 22963 45758 22997 45780
rect 22997 45758 23006 45780
rect 23040 45674 23049 45696
rect 23049 45674 23083 45696
rect 23083 45674 23092 45696
rect 23040 45644 23092 45674
rect 23040 45602 23049 45632
rect 23049 45602 23083 45632
rect 23083 45602 23092 45632
rect 23040 45580 23092 45602
rect 22893 45410 23067 45470
rect 23314 45901 23384 45918
rect 23314 45504 23330 45901
rect 23330 45504 23368 45901
rect 23368 45504 23384 45901
rect 23314 45486 23384 45504
rect 31776 45901 31846 45918
rect 31776 45504 31792 45901
rect 31792 45504 31830 45901
rect 31830 45504 31846 45901
rect 31776 45486 31846 45504
rect 32068 45674 32077 45696
rect 32077 45674 32111 45696
rect 32111 45674 32120 45696
rect 32068 45644 32120 45674
rect 32068 45602 32077 45632
rect 32077 45602 32111 45632
rect 32111 45602 32120 45632
rect 32068 45580 32120 45602
rect 32154 45852 32206 45874
rect 32154 45822 32163 45852
rect 32163 45822 32197 45852
rect 32197 45822 32206 45852
rect 32154 45780 32206 45810
rect 32154 45758 32163 45780
rect 32163 45758 32197 45780
rect 32197 45758 32206 45780
rect 32240 45674 32249 45696
rect 32249 45674 32283 45696
rect 32283 45674 32292 45696
rect 32240 45644 32292 45674
rect 32240 45602 32249 45632
rect 32249 45602 32283 45632
rect 32283 45602 32292 45632
rect 32240 45580 32292 45602
rect 32093 45410 32267 45470
rect 32514 45901 32584 45918
rect 32514 45504 32530 45901
rect 32530 45504 32568 45901
rect 32568 45504 32584 45901
rect 32514 45486 32584 45504
rect 40976 45901 41046 45918
rect 40976 45504 40992 45901
rect 40992 45504 41030 45901
rect 41030 45504 41046 45901
rect 40976 45486 41046 45504
rect 41268 45674 41277 45696
rect 41277 45674 41311 45696
rect 41311 45674 41320 45696
rect 41268 45644 41320 45674
rect 41268 45602 41277 45632
rect 41277 45602 41311 45632
rect 41311 45602 41320 45632
rect 41268 45580 41320 45602
rect 41354 45852 41406 45874
rect 41354 45822 41363 45852
rect 41363 45822 41397 45852
rect 41397 45822 41406 45852
rect 41354 45780 41406 45810
rect 41354 45758 41363 45780
rect 41363 45758 41397 45780
rect 41397 45758 41406 45780
rect 41440 45674 41449 45696
rect 41449 45674 41483 45696
rect 41483 45674 41492 45696
rect 41440 45644 41492 45674
rect 41440 45602 41449 45632
rect 41449 45602 41483 45632
rect 41483 45602 41492 45632
rect 41440 45580 41492 45602
rect 41293 45410 41467 45470
rect 41714 45901 41784 45918
rect 41714 45504 41730 45901
rect 41730 45504 41768 45901
rect 41768 45504 41784 45901
rect 41714 45486 41784 45504
rect 50176 45901 50246 45918
rect 50176 45504 50192 45901
rect 50192 45504 50230 45901
rect 50230 45504 50246 45901
rect 50176 45486 50246 45504
rect 50468 45674 50477 45696
rect 50477 45674 50511 45696
rect 50511 45674 50520 45696
rect 50468 45644 50520 45674
rect 50468 45602 50477 45632
rect 50477 45602 50511 45632
rect 50511 45602 50520 45632
rect 50468 45580 50520 45602
rect 50554 45852 50606 45874
rect 50554 45822 50563 45852
rect 50563 45822 50597 45852
rect 50597 45822 50606 45852
rect 50554 45780 50606 45810
rect 50554 45758 50563 45780
rect 50563 45758 50597 45780
rect 50597 45758 50606 45780
rect 50640 45674 50649 45696
rect 50649 45674 50683 45696
rect 50683 45674 50692 45696
rect 50640 45644 50692 45674
rect 50640 45602 50649 45632
rect 50649 45602 50683 45632
rect 50683 45602 50692 45632
rect 50640 45580 50692 45602
rect 50493 45410 50667 45470
rect 50914 45901 50984 45918
rect 50914 45504 50930 45901
rect 50930 45504 50968 45901
rect 50968 45504 50984 45901
rect 50914 45486 50984 45504
rect 59376 45901 59446 45918
rect 59376 45504 59392 45901
rect 59392 45504 59430 45901
rect 59430 45504 59446 45901
rect 59376 45486 59446 45504
rect 59668 45674 59677 45696
rect 59677 45674 59711 45696
rect 59711 45674 59720 45696
rect 59668 45644 59720 45674
rect 59668 45602 59677 45632
rect 59677 45602 59711 45632
rect 59711 45602 59720 45632
rect 59668 45580 59720 45602
rect 59754 45852 59806 45874
rect 59754 45822 59763 45852
rect 59763 45822 59797 45852
rect 59797 45822 59806 45852
rect 59754 45780 59806 45810
rect 59754 45758 59763 45780
rect 59763 45758 59797 45780
rect 59797 45758 59806 45780
rect 59840 45674 59849 45696
rect 59849 45674 59883 45696
rect 59883 45674 59892 45696
rect 59840 45644 59892 45674
rect 59840 45602 59849 45632
rect 59849 45602 59883 45632
rect 59883 45602 59892 45632
rect 59840 45580 59892 45602
rect 59693 45410 59867 45470
rect 60114 45901 60184 45918
rect 60114 45504 60130 45901
rect 60130 45504 60168 45901
rect 60168 45504 60184 45901
rect 60114 45486 60184 45504
rect 68576 45901 68646 45918
rect 68576 45504 68592 45901
rect 68592 45504 68630 45901
rect 68630 45504 68646 45901
rect 68576 45486 68646 45504
rect 68868 45674 68877 45696
rect 68877 45674 68911 45696
rect 68911 45674 68920 45696
rect 68868 45644 68920 45674
rect 68868 45602 68877 45632
rect 68877 45602 68911 45632
rect 68911 45602 68920 45632
rect 68868 45580 68920 45602
rect 68954 45852 69006 45874
rect 68954 45822 68963 45852
rect 68963 45822 68997 45852
rect 68997 45822 69006 45852
rect 68954 45780 69006 45810
rect 68954 45758 68963 45780
rect 68963 45758 68997 45780
rect 68997 45758 69006 45780
rect 69040 45674 69049 45696
rect 69049 45674 69083 45696
rect 69083 45674 69092 45696
rect 69040 45644 69092 45674
rect 69040 45602 69049 45632
rect 69049 45602 69083 45632
rect 69083 45602 69092 45632
rect 69040 45580 69092 45602
rect 68893 45410 69067 45470
rect 69314 45901 69384 45918
rect 69314 45504 69330 45901
rect 69330 45504 69368 45901
rect 69368 45504 69384 45901
rect 69314 45486 69384 45504
rect 4176 36021 4246 36038
rect 4176 35624 4192 36021
rect 4192 35624 4230 36021
rect 4230 35624 4246 36021
rect 4176 35606 4246 35624
rect 4468 35794 4477 35816
rect 4477 35794 4511 35816
rect 4511 35794 4520 35816
rect 4468 35764 4520 35794
rect 4468 35722 4477 35752
rect 4477 35722 4511 35752
rect 4511 35722 4520 35752
rect 4468 35700 4520 35722
rect 4554 35972 4606 35994
rect 4554 35942 4563 35972
rect 4563 35942 4597 35972
rect 4597 35942 4606 35972
rect 4554 35900 4606 35930
rect 4554 35878 4563 35900
rect 4563 35878 4597 35900
rect 4597 35878 4606 35900
rect 4640 35794 4649 35816
rect 4649 35794 4683 35816
rect 4683 35794 4692 35816
rect 4640 35764 4692 35794
rect 4640 35722 4649 35752
rect 4649 35722 4683 35752
rect 4683 35722 4692 35752
rect 4640 35700 4692 35722
rect 4493 35530 4667 35590
rect 4914 36021 4984 36038
rect 4914 35624 4930 36021
rect 4930 35624 4968 36021
rect 4968 35624 4984 36021
rect 4914 35606 4984 35624
rect 13376 36021 13446 36038
rect 13376 35624 13392 36021
rect 13392 35624 13430 36021
rect 13430 35624 13446 36021
rect 13376 35606 13446 35624
rect 13668 35794 13677 35816
rect 13677 35794 13711 35816
rect 13711 35794 13720 35816
rect 13668 35764 13720 35794
rect 13668 35722 13677 35752
rect 13677 35722 13711 35752
rect 13711 35722 13720 35752
rect 13668 35700 13720 35722
rect 13754 35972 13806 35994
rect 13754 35942 13763 35972
rect 13763 35942 13797 35972
rect 13797 35942 13806 35972
rect 13754 35900 13806 35930
rect 13754 35878 13763 35900
rect 13763 35878 13797 35900
rect 13797 35878 13806 35900
rect 13840 35794 13849 35816
rect 13849 35794 13883 35816
rect 13883 35794 13892 35816
rect 13840 35764 13892 35794
rect 13840 35722 13849 35752
rect 13849 35722 13883 35752
rect 13883 35722 13892 35752
rect 13840 35700 13892 35722
rect 13693 35530 13867 35590
rect 14114 36021 14184 36038
rect 14114 35624 14130 36021
rect 14130 35624 14168 36021
rect 14168 35624 14184 36021
rect 14114 35606 14184 35624
rect 22576 36021 22646 36038
rect 22576 35624 22592 36021
rect 22592 35624 22630 36021
rect 22630 35624 22646 36021
rect 22576 35606 22646 35624
rect 22868 35794 22877 35816
rect 22877 35794 22911 35816
rect 22911 35794 22920 35816
rect 22868 35764 22920 35794
rect 22868 35722 22877 35752
rect 22877 35722 22911 35752
rect 22911 35722 22920 35752
rect 22868 35700 22920 35722
rect 22954 35972 23006 35994
rect 22954 35942 22963 35972
rect 22963 35942 22997 35972
rect 22997 35942 23006 35972
rect 22954 35900 23006 35930
rect 22954 35878 22963 35900
rect 22963 35878 22997 35900
rect 22997 35878 23006 35900
rect 23040 35794 23049 35816
rect 23049 35794 23083 35816
rect 23083 35794 23092 35816
rect 23040 35764 23092 35794
rect 23040 35722 23049 35752
rect 23049 35722 23083 35752
rect 23083 35722 23092 35752
rect 23040 35700 23092 35722
rect 22893 35530 23067 35590
rect 23314 36021 23384 36038
rect 23314 35624 23330 36021
rect 23330 35624 23368 36021
rect 23368 35624 23384 36021
rect 23314 35606 23384 35624
rect 31776 36021 31846 36038
rect 31776 35624 31792 36021
rect 31792 35624 31830 36021
rect 31830 35624 31846 36021
rect 31776 35606 31846 35624
rect 32068 35794 32077 35816
rect 32077 35794 32111 35816
rect 32111 35794 32120 35816
rect 32068 35764 32120 35794
rect 32068 35722 32077 35752
rect 32077 35722 32111 35752
rect 32111 35722 32120 35752
rect 32068 35700 32120 35722
rect 32154 35972 32206 35994
rect 32154 35942 32163 35972
rect 32163 35942 32197 35972
rect 32197 35942 32206 35972
rect 32154 35900 32206 35930
rect 32154 35878 32163 35900
rect 32163 35878 32197 35900
rect 32197 35878 32206 35900
rect 32240 35794 32249 35816
rect 32249 35794 32283 35816
rect 32283 35794 32292 35816
rect 32240 35764 32292 35794
rect 32240 35722 32249 35752
rect 32249 35722 32283 35752
rect 32283 35722 32292 35752
rect 32240 35700 32292 35722
rect 32093 35530 32267 35590
rect 32514 36021 32584 36038
rect 32514 35624 32530 36021
rect 32530 35624 32568 36021
rect 32568 35624 32584 36021
rect 32514 35606 32584 35624
rect 40976 36021 41046 36038
rect 40976 35624 40992 36021
rect 40992 35624 41030 36021
rect 41030 35624 41046 36021
rect 40976 35606 41046 35624
rect 41268 35794 41277 35816
rect 41277 35794 41311 35816
rect 41311 35794 41320 35816
rect 41268 35764 41320 35794
rect 41268 35722 41277 35752
rect 41277 35722 41311 35752
rect 41311 35722 41320 35752
rect 41268 35700 41320 35722
rect 41354 35972 41406 35994
rect 41354 35942 41363 35972
rect 41363 35942 41397 35972
rect 41397 35942 41406 35972
rect 41354 35900 41406 35930
rect 41354 35878 41363 35900
rect 41363 35878 41397 35900
rect 41397 35878 41406 35900
rect 41440 35794 41449 35816
rect 41449 35794 41483 35816
rect 41483 35794 41492 35816
rect 41440 35764 41492 35794
rect 41440 35722 41449 35752
rect 41449 35722 41483 35752
rect 41483 35722 41492 35752
rect 41440 35700 41492 35722
rect 41293 35530 41467 35590
rect 41714 36021 41784 36038
rect 41714 35624 41730 36021
rect 41730 35624 41768 36021
rect 41768 35624 41784 36021
rect 41714 35606 41784 35624
rect 50176 36021 50246 36038
rect 50176 35624 50192 36021
rect 50192 35624 50230 36021
rect 50230 35624 50246 36021
rect 50176 35606 50246 35624
rect 50468 35794 50477 35816
rect 50477 35794 50511 35816
rect 50511 35794 50520 35816
rect 50468 35764 50520 35794
rect 50468 35722 50477 35752
rect 50477 35722 50511 35752
rect 50511 35722 50520 35752
rect 50468 35700 50520 35722
rect 50554 35972 50606 35994
rect 50554 35942 50563 35972
rect 50563 35942 50597 35972
rect 50597 35942 50606 35972
rect 50554 35900 50606 35930
rect 50554 35878 50563 35900
rect 50563 35878 50597 35900
rect 50597 35878 50606 35900
rect 50640 35794 50649 35816
rect 50649 35794 50683 35816
rect 50683 35794 50692 35816
rect 50640 35764 50692 35794
rect 50640 35722 50649 35752
rect 50649 35722 50683 35752
rect 50683 35722 50692 35752
rect 50640 35700 50692 35722
rect 50493 35530 50667 35590
rect 50914 36021 50984 36038
rect 50914 35624 50930 36021
rect 50930 35624 50968 36021
rect 50968 35624 50984 36021
rect 50914 35606 50984 35624
rect 59376 36021 59446 36038
rect 59376 35624 59392 36021
rect 59392 35624 59430 36021
rect 59430 35624 59446 36021
rect 59376 35606 59446 35624
rect 59668 35794 59677 35816
rect 59677 35794 59711 35816
rect 59711 35794 59720 35816
rect 59668 35764 59720 35794
rect 59668 35722 59677 35752
rect 59677 35722 59711 35752
rect 59711 35722 59720 35752
rect 59668 35700 59720 35722
rect 59754 35972 59806 35994
rect 59754 35942 59763 35972
rect 59763 35942 59797 35972
rect 59797 35942 59806 35972
rect 59754 35900 59806 35930
rect 59754 35878 59763 35900
rect 59763 35878 59797 35900
rect 59797 35878 59806 35900
rect 59840 35794 59849 35816
rect 59849 35794 59883 35816
rect 59883 35794 59892 35816
rect 59840 35764 59892 35794
rect 59840 35722 59849 35752
rect 59849 35722 59883 35752
rect 59883 35722 59892 35752
rect 59840 35700 59892 35722
rect 59693 35530 59867 35590
rect 60114 36021 60184 36038
rect 60114 35624 60130 36021
rect 60130 35624 60168 36021
rect 60168 35624 60184 36021
rect 60114 35606 60184 35624
rect 68576 36021 68646 36038
rect 68576 35624 68592 36021
rect 68592 35624 68630 36021
rect 68630 35624 68646 36021
rect 68576 35606 68646 35624
rect 68868 35794 68877 35816
rect 68877 35794 68911 35816
rect 68911 35794 68920 35816
rect 68868 35764 68920 35794
rect 68868 35722 68877 35752
rect 68877 35722 68911 35752
rect 68911 35722 68920 35752
rect 68868 35700 68920 35722
rect 68954 35972 69006 35994
rect 68954 35942 68963 35972
rect 68963 35942 68997 35972
rect 68997 35942 69006 35972
rect 68954 35900 69006 35930
rect 68954 35878 68963 35900
rect 68963 35878 68997 35900
rect 68997 35878 69006 35900
rect 69040 35794 69049 35816
rect 69049 35794 69083 35816
rect 69083 35794 69092 35816
rect 69040 35764 69092 35794
rect 69040 35722 69049 35752
rect 69049 35722 69083 35752
rect 69083 35722 69092 35752
rect 69040 35700 69092 35722
rect 68893 35530 69067 35590
rect 69314 36021 69384 36038
rect 69314 35624 69330 36021
rect 69330 35624 69368 36021
rect 69368 35624 69384 36021
rect 69314 35606 69384 35624
rect 4176 26141 4246 26158
rect 4176 25744 4192 26141
rect 4192 25744 4230 26141
rect 4230 25744 4246 26141
rect 4176 25726 4246 25744
rect 4468 25914 4477 25936
rect 4477 25914 4511 25936
rect 4511 25914 4520 25936
rect 4468 25884 4520 25914
rect 4468 25842 4477 25872
rect 4477 25842 4511 25872
rect 4511 25842 4520 25872
rect 4468 25820 4520 25842
rect 4554 26092 4606 26114
rect 4554 26062 4563 26092
rect 4563 26062 4597 26092
rect 4597 26062 4606 26092
rect 4554 26020 4606 26050
rect 4554 25998 4563 26020
rect 4563 25998 4597 26020
rect 4597 25998 4606 26020
rect 4640 25914 4649 25936
rect 4649 25914 4683 25936
rect 4683 25914 4692 25936
rect 4640 25884 4692 25914
rect 4640 25842 4649 25872
rect 4649 25842 4683 25872
rect 4683 25842 4692 25872
rect 4640 25820 4692 25842
rect 4493 25650 4667 25710
rect 4914 26141 4984 26158
rect 4914 25744 4930 26141
rect 4930 25744 4968 26141
rect 4968 25744 4984 26141
rect 4914 25726 4984 25744
rect 13376 26141 13446 26158
rect 13376 25744 13392 26141
rect 13392 25744 13430 26141
rect 13430 25744 13446 26141
rect 13376 25726 13446 25744
rect 13668 25914 13677 25936
rect 13677 25914 13711 25936
rect 13711 25914 13720 25936
rect 13668 25884 13720 25914
rect 13668 25842 13677 25872
rect 13677 25842 13711 25872
rect 13711 25842 13720 25872
rect 13668 25820 13720 25842
rect 13754 26092 13806 26114
rect 13754 26062 13763 26092
rect 13763 26062 13797 26092
rect 13797 26062 13806 26092
rect 13754 26020 13806 26050
rect 13754 25998 13763 26020
rect 13763 25998 13797 26020
rect 13797 25998 13806 26020
rect 13840 25914 13849 25936
rect 13849 25914 13883 25936
rect 13883 25914 13892 25936
rect 13840 25884 13892 25914
rect 13840 25842 13849 25872
rect 13849 25842 13883 25872
rect 13883 25842 13892 25872
rect 13840 25820 13892 25842
rect 13693 25650 13867 25710
rect 14114 26141 14184 26158
rect 14114 25744 14130 26141
rect 14130 25744 14168 26141
rect 14168 25744 14184 26141
rect 14114 25726 14184 25744
rect 22576 26141 22646 26158
rect 22576 25744 22592 26141
rect 22592 25744 22630 26141
rect 22630 25744 22646 26141
rect 22576 25726 22646 25744
rect 22868 25914 22877 25936
rect 22877 25914 22911 25936
rect 22911 25914 22920 25936
rect 22868 25884 22920 25914
rect 22868 25842 22877 25872
rect 22877 25842 22911 25872
rect 22911 25842 22920 25872
rect 22868 25820 22920 25842
rect 22954 26092 23006 26114
rect 22954 26062 22963 26092
rect 22963 26062 22997 26092
rect 22997 26062 23006 26092
rect 22954 26020 23006 26050
rect 22954 25998 22963 26020
rect 22963 25998 22997 26020
rect 22997 25998 23006 26020
rect 23040 25914 23049 25936
rect 23049 25914 23083 25936
rect 23083 25914 23092 25936
rect 23040 25884 23092 25914
rect 23040 25842 23049 25872
rect 23049 25842 23083 25872
rect 23083 25842 23092 25872
rect 23040 25820 23092 25842
rect 22893 25650 23067 25710
rect 23314 26141 23384 26158
rect 23314 25744 23330 26141
rect 23330 25744 23368 26141
rect 23368 25744 23384 26141
rect 23314 25726 23384 25744
rect 31776 26141 31846 26158
rect 31776 25744 31792 26141
rect 31792 25744 31830 26141
rect 31830 25744 31846 26141
rect 31776 25726 31846 25744
rect 32068 25914 32077 25936
rect 32077 25914 32111 25936
rect 32111 25914 32120 25936
rect 32068 25884 32120 25914
rect 32068 25842 32077 25872
rect 32077 25842 32111 25872
rect 32111 25842 32120 25872
rect 32068 25820 32120 25842
rect 32154 26092 32206 26114
rect 32154 26062 32163 26092
rect 32163 26062 32197 26092
rect 32197 26062 32206 26092
rect 32154 26020 32206 26050
rect 32154 25998 32163 26020
rect 32163 25998 32197 26020
rect 32197 25998 32206 26020
rect 32240 25914 32249 25936
rect 32249 25914 32283 25936
rect 32283 25914 32292 25936
rect 32240 25884 32292 25914
rect 32240 25842 32249 25872
rect 32249 25842 32283 25872
rect 32283 25842 32292 25872
rect 32240 25820 32292 25842
rect 32093 25650 32267 25710
rect 32514 26141 32584 26158
rect 32514 25744 32530 26141
rect 32530 25744 32568 26141
rect 32568 25744 32584 26141
rect 32514 25726 32584 25744
rect 40976 26141 41046 26158
rect 40976 25744 40992 26141
rect 40992 25744 41030 26141
rect 41030 25744 41046 26141
rect 40976 25726 41046 25744
rect 41268 25914 41277 25936
rect 41277 25914 41311 25936
rect 41311 25914 41320 25936
rect 41268 25884 41320 25914
rect 41268 25842 41277 25872
rect 41277 25842 41311 25872
rect 41311 25842 41320 25872
rect 41268 25820 41320 25842
rect 41354 26092 41406 26114
rect 41354 26062 41363 26092
rect 41363 26062 41397 26092
rect 41397 26062 41406 26092
rect 41354 26020 41406 26050
rect 41354 25998 41363 26020
rect 41363 25998 41397 26020
rect 41397 25998 41406 26020
rect 41440 25914 41449 25936
rect 41449 25914 41483 25936
rect 41483 25914 41492 25936
rect 41440 25884 41492 25914
rect 41440 25842 41449 25872
rect 41449 25842 41483 25872
rect 41483 25842 41492 25872
rect 41440 25820 41492 25842
rect 41293 25650 41467 25710
rect 41714 26141 41784 26158
rect 41714 25744 41730 26141
rect 41730 25744 41768 26141
rect 41768 25744 41784 26141
rect 41714 25726 41784 25744
rect 50176 26141 50246 26158
rect 50176 25744 50192 26141
rect 50192 25744 50230 26141
rect 50230 25744 50246 26141
rect 50176 25726 50246 25744
rect 50468 25914 50477 25936
rect 50477 25914 50511 25936
rect 50511 25914 50520 25936
rect 50468 25884 50520 25914
rect 50468 25842 50477 25872
rect 50477 25842 50511 25872
rect 50511 25842 50520 25872
rect 50468 25820 50520 25842
rect 50554 26092 50606 26114
rect 50554 26062 50563 26092
rect 50563 26062 50597 26092
rect 50597 26062 50606 26092
rect 50554 26020 50606 26050
rect 50554 25998 50563 26020
rect 50563 25998 50597 26020
rect 50597 25998 50606 26020
rect 50640 25914 50649 25936
rect 50649 25914 50683 25936
rect 50683 25914 50692 25936
rect 50640 25884 50692 25914
rect 50640 25842 50649 25872
rect 50649 25842 50683 25872
rect 50683 25842 50692 25872
rect 50640 25820 50692 25842
rect 50493 25650 50667 25710
rect 50914 26141 50984 26158
rect 50914 25744 50930 26141
rect 50930 25744 50968 26141
rect 50968 25744 50984 26141
rect 50914 25726 50984 25744
rect 59376 26141 59446 26158
rect 59376 25744 59392 26141
rect 59392 25744 59430 26141
rect 59430 25744 59446 26141
rect 59376 25726 59446 25744
rect 59668 25914 59677 25936
rect 59677 25914 59711 25936
rect 59711 25914 59720 25936
rect 59668 25884 59720 25914
rect 59668 25842 59677 25872
rect 59677 25842 59711 25872
rect 59711 25842 59720 25872
rect 59668 25820 59720 25842
rect 59754 26092 59806 26114
rect 59754 26062 59763 26092
rect 59763 26062 59797 26092
rect 59797 26062 59806 26092
rect 59754 26020 59806 26050
rect 59754 25998 59763 26020
rect 59763 25998 59797 26020
rect 59797 25998 59806 26020
rect 59840 25914 59849 25936
rect 59849 25914 59883 25936
rect 59883 25914 59892 25936
rect 59840 25884 59892 25914
rect 59840 25842 59849 25872
rect 59849 25842 59883 25872
rect 59883 25842 59892 25872
rect 59840 25820 59892 25842
rect 59693 25650 59867 25710
rect 60114 26141 60184 26158
rect 60114 25744 60130 26141
rect 60130 25744 60168 26141
rect 60168 25744 60184 26141
rect 60114 25726 60184 25744
rect 68576 26141 68646 26158
rect 68576 25744 68592 26141
rect 68592 25744 68630 26141
rect 68630 25744 68646 26141
rect 68576 25726 68646 25744
rect 68868 25914 68877 25936
rect 68877 25914 68911 25936
rect 68911 25914 68920 25936
rect 68868 25884 68920 25914
rect 68868 25842 68877 25872
rect 68877 25842 68911 25872
rect 68911 25842 68920 25872
rect 68868 25820 68920 25842
rect 68954 26092 69006 26114
rect 68954 26062 68963 26092
rect 68963 26062 68997 26092
rect 68997 26062 69006 26092
rect 68954 26020 69006 26050
rect 68954 25998 68963 26020
rect 68963 25998 68997 26020
rect 68997 25998 69006 26020
rect 69040 25914 69049 25936
rect 69049 25914 69083 25936
rect 69083 25914 69092 25936
rect 69040 25884 69092 25914
rect 69040 25842 69049 25872
rect 69049 25842 69083 25872
rect 69083 25842 69092 25872
rect 69040 25820 69092 25842
rect 68893 25650 69067 25710
rect 69314 26141 69384 26158
rect 69314 25744 69330 26141
rect 69330 25744 69368 26141
rect 69368 25744 69384 26141
rect 69314 25726 69384 25744
rect 4176 16261 4246 16278
rect 4176 15864 4192 16261
rect 4192 15864 4230 16261
rect 4230 15864 4246 16261
rect 4176 15846 4246 15864
rect 4468 16034 4477 16056
rect 4477 16034 4511 16056
rect 4511 16034 4520 16056
rect 4468 16004 4520 16034
rect 4468 15962 4477 15992
rect 4477 15962 4511 15992
rect 4511 15962 4520 15992
rect 4468 15940 4520 15962
rect 4554 16212 4606 16234
rect 4554 16182 4563 16212
rect 4563 16182 4597 16212
rect 4597 16182 4606 16212
rect 4554 16140 4606 16170
rect 4554 16118 4563 16140
rect 4563 16118 4597 16140
rect 4597 16118 4606 16140
rect 4640 16034 4649 16056
rect 4649 16034 4683 16056
rect 4683 16034 4692 16056
rect 4640 16004 4692 16034
rect 4640 15962 4649 15992
rect 4649 15962 4683 15992
rect 4683 15962 4692 15992
rect 4640 15940 4692 15962
rect 4493 15770 4667 15830
rect 4914 16261 4984 16278
rect 4914 15864 4930 16261
rect 4930 15864 4968 16261
rect 4968 15864 4984 16261
rect 4914 15846 4984 15864
rect 13376 16261 13446 16278
rect 13376 15864 13392 16261
rect 13392 15864 13430 16261
rect 13430 15864 13446 16261
rect 13376 15846 13446 15864
rect 13668 16034 13677 16056
rect 13677 16034 13711 16056
rect 13711 16034 13720 16056
rect 13668 16004 13720 16034
rect 13668 15962 13677 15992
rect 13677 15962 13711 15992
rect 13711 15962 13720 15992
rect 13668 15940 13720 15962
rect 13754 16212 13806 16234
rect 13754 16182 13763 16212
rect 13763 16182 13797 16212
rect 13797 16182 13806 16212
rect 13754 16140 13806 16170
rect 13754 16118 13763 16140
rect 13763 16118 13797 16140
rect 13797 16118 13806 16140
rect 13840 16034 13849 16056
rect 13849 16034 13883 16056
rect 13883 16034 13892 16056
rect 13840 16004 13892 16034
rect 13840 15962 13849 15992
rect 13849 15962 13883 15992
rect 13883 15962 13892 15992
rect 13840 15940 13892 15962
rect 13693 15770 13867 15830
rect 14114 16261 14184 16278
rect 14114 15864 14130 16261
rect 14130 15864 14168 16261
rect 14168 15864 14184 16261
rect 14114 15846 14184 15864
rect 22576 16261 22646 16278
rect 22576 15864 22592 16261
rect 22592 15864 22630 16261
rect 22630 15864 22646 16261
rect 22576 15846 22646 15864
rect 22868 16034 22877 16056
rect 22877 16034 22911 16056
rect 22911 16034 22920 16056
rect 22868 16004 22920 16034
rect 22868 15962 22877 15992
rect 22877 15962 22911 15992
rect 22911 15962 22920 15992
rect 22868 15940 22920 15962
rect 22954 16212 23006 16234
rect 22954 16182 22963 16212
rect 22963 16182 22997 16212
rect 22997 16182 23006 16212
rect 22954 16140 23006 16170
rect 22954 16118 22963 16140
rect 22963 16118 22997 16140
rect 22997 16118 23006 16140
rect 23040 16034 23049 16056
rect 23049 16034 23083 16056
rect 23083 16034 23092 16056
rect 23040 16004 23092 16034
rect 23040 15962 23049 15992
rect 23049 15962 23083 15992
rect 23083 15962 23092 15992
rect 23040 15940 23092 15962
rect 22893 15770 23067 15830
rect 23314 16261 23384 16278
rect 23314 15864 23330 16261
rect 23330 15864 23368 16261
rect 23368 15864 23384 16261
rect 23314 15846 23384 15864
rect 31776 16261 31846 16278
rect 31776 15864 31792 16261
rect 31792 15864 31830 16261
rect 31830 15864 31846 16261
rect 31776 15846 31846 15864
rect 32068 16034 32077 16056
rect 32077 16034 32111 16056
rect 32111 16034 32120 16056
rect 32068 16004 32120 16034
rect 32068 15962 32077 15992
rect 32077 15962 32111 15992
rect 32111 15962 32120 15992
rect 32068 15940 32120 15962
rect 32154 16212 32206 16234
rect 32154 16182 32163 16212
rect 32163 16182 32197 16212
rect 32197 16182 32206 16212
rect 32154 16140 32206 16170
rect 32154 16118 32163 16140
rect 32163 16118 32197 16140
rect 32197 16118 32206 16140
rect 32240 16034 32249 16056
rect 32249 16034 32283 16056
rect 32283 16034 32292 16056
rect 32240 16004 32292 16034
rect 32240 15962 32249 15992
rect 32249 15962 32283 15992
rect 32283 15962 32292 15992
rect 32240 15940 32292 15962
rect 32093 15770 32267 15830
rect 32514 16261 32584 16278
rect 32514 15864 32530 16261
rect 32530 15864 32568 16261
rect 32568 15864 32584 16261
rect 32514 15846 32584 15864
rect 40976 16261 41046 16278
rect 40976 15864 40992 16261
rect 40992 15864 41030 16261
rect 41030 15864 41046 16261
rect 40976 15846 41046 15864
rect 41268 16034 41277 16056
rect 41277 16034 41311 16056
rect 41311 16034 41320 16056
rect 41268 16004 41320 16034
rect 41268 15962 41277 15992
rect 41277 15962 41311 15992
rect 41311 15962 41320 15992
rect 41268 15940 41320 15962
rect 41354 16212 41406 16234
rect 41354 16182 41363 16212
rect 41363 16182 41397 16212
rect 41397 16182 41406 16212
rect 41354 16140 41406 16170
rect 41354 16118 41363 16140
rect 41363 16118 41397 16140
rect 41397 16118 41406 16140
rect 41440 16034 41449 16056
rect 41449 16034 41483 16056
rect 41483 16034 41492 16056
rect 41440 16004 41492 16034
rect 41440 15962 41449 15992
rect 41449 15962 41483 15992
rect 41483 15962 41492 15992
rect 41440 15940 41492 15962
rect 41293 15770 41467 15830
rect 41714 16261 41784 16278
rect 41714 15864 41730 16261
rect 41730 15864 41768 16261
rect 41768 15864 41784 16261
rect 41714 15846 41784 15864
rect 50176 16261 50246 16278
rect 50176 15864 50192 16261
rect 50192 15864 50230 16261
rect 50230 15864 50246 16261
rect 50176 15846 50246 15864
rect 50468 16034 50477 16056
rect 50477 16034 50511 16056
rect 50511 16034 50520 16056
rect 50468 16004 50520 16034
rect 50468 15962 50477 15992
rect 50477 15962 50511 15992
rect 50511 15962 50520 15992
rect 50468 15940 50520 15962
rect 50554 16212 50606 16234
rect 50554 16182 50563 16212
rect 50563 16182 50597 16212
rect 50597 16182 50606 16212
rect 50554 16140 50606 16170
rect 50554 16118 50563 16140
rect 50563 16118 50597 16140
rect 50597 16118 50606 16140
rect 50640 16034 50649 16056
rect 50649 16034 50683 16056
rect 50683 16034 50692 16056
rect 50640 16004 50692 16034
rect 50640 15962 50649 15992
rect 50649 15962 50683 15992
rect 50683 15962 50692 15992
rect 50640 15940 50692 15962
rect 50493 15770 50667 15830
rect 50914 16261 50984 16278
rect 50914 15864 50930 16261
rect 50930 15864 50968 16261
rect 50968 15864 50984 16261
rect 50914 15846 50984 15864
rect 59376 16261 59446 16278
rect 59376 15864 59392 16261
rect 59392 15864 59430 16261
rect 59430 15864 59446 16261
rect 59376 15846 59446 15864
rect 59668 16034 59677 16056
rect 59677 16034 59711 16056
rect 59711 16034 59720 16056
rect 59668 16004 59720 16034
rect 59668 15962 59677 15992
rect 59677 15962 59711 15992
rect 59711 15962 59720 15992
rect 59668 15940 59720 15962
rect 59754 16212 59806 16234
rect 59754 16182 59763 16212
rect 59763 16182 59797 16212
rect 59797 16182 59806 16212
rect 59754 16140 59806 16170
rect 59754 16118 59763 16140
rect 59763 16118 59797 16140
rect 59797 16118 59806 16140
rect 59840 16034 59849 16056
rect 59849 16034 59883 16056
rect 59883 16034 59892 16056
rect 59840 16004 59892 16034
rect 59840 15962 59849 15992
rect 59849 15962 59883 15992
rect 59883 15962 59892 15992
rect 59840 15940 59892 15962
rect 59693 15770 59867 15830
rect 60114 16261 60184 16278
rect 60114 15864 60130 16261
rect 60130 15864 60168 16261
rect 60168 15864 60184 16261
rect 60114 15846 60184 15864
rect 68576 16261 68646 16278
rect 68576 15864 68592 16261
rect 68592 15864 68630 16261
rect 68630 15864 68646 16261
rect 68576 15846 68646 15864
rect 68868 16034 68877 16056
rect 68877 16034 68911 16056
rect 68911 16034 68920 16056
rect 68868 16004 68920 16034
rect 68868 15962 68877 15992
rect 68877 15962 68911 15992
rect 68911 15962 68920 15992
rect 68868 15940 68920 15962
rect 68954 16212 69006 16234
rect 68954 16182 68963 16212
rect 68963 16182 68997 16212
rect 68997 16182 69006 16212
rect 68954 16140 69006 16170
rect 68954 16118 68963 16140
rect 68963 16118 68997 16140
rect 68997 16118 69006 16140
rect 69040 16034 69049 16056
rect 69049 16034 69083 16056
rect 69083 16034 69092 16056
rect 69040 16004 69092 16034
rect 69040 15962 69049 15992
rect 69049 15962 69083 15992
rect 69083 15962 69092 15992
rect 69040 15940 69092 15962
rect 68893 15770 69067 15830
rect 69314 16261 69384 16278
rect 69314 15864 69330 16261
rect 69330 15864 69368 16261
rect 69368 15864 69384 16261
rect 69314 15846 69384 15864
rect -490 6610 -240 6620
rect -490 6570 -480 6610
rect -480 6570 -440 6610
rect -440 6570 -400 6610
rect -400 6570 -360 6610
rect -360 6570 -310 6610
rect -310 6570 -270 6610
rect -270 6570 -240 6610
rect -490 6560 -240 6570
rect 4176 6381 4246 6398
rect 4176 5984 4192 6381
rect 4192 5984 4230 6381
rect 4230 5984 4246 6381
rect 4176 5966 4246 5984
rect 4468 6154 4477 6176
rect 4477 6154 4511 6176
rect 4511 6154 4520 6176
rect 4468 6124 4520 6154
rect 4468 6082 4477 6112
rect 4477 6082 4511 6112
rect 4511 6082 4520 6112
rect 4468 6060 4520 6082
rect 4554 6332 4606 6354
rect 4554 6302 4563 6332
rect 4563 6302 4597 6332
rect 4597 6302 4606 6332
rect 4554 6260 4606 6290
rect 4554 6238 4563 6260
rect 4563 6238 4597 6260
rect 4597 6238 4606 6260
rect 4640 6154 4649 6176
rect 4649 6154 4683 6176
rect 4683 6154 4692 6176
rect 4640 6124 4692 6154
rect 4640 6082 4649 6112
rect 4649 6082 4683 6112
rect 4683 6082 4692 6112
rect 4640 6060 4692 6082
rect 4493 5890 4667 5950
rect -230 5820 -170 5830
rect -230 5780 -220 5820
rect -220 5780 -180 5820
rect -180 5780 -170 5820
rect -230 5770 -170 5780
rect 4914 6381 4984 6398
rect 4914 5984 4930 6381
rect 4930 5984 4968 6381
rect 4968 5984 4984 6381
rect 4914 5966 4984 5984
rect 13376 6381 13446 6398
rect 13376 5984 13392 6381
rect 13392 5984 13430 6381
rect 13430 5984 13446 6381
rect 13376 5966 13446 5984
rect 13668 6154 13677 6176
rect 13677 6154 13711 6176
rect 13711 6154 13720 6176
rect 13668 6124 13720 6154
rect 13668 6082 13677 6112
rect 13677 6082 13711 6112
rect 13711 6082 13720 6112
rect 13668 6060 13720 6082
rect 13754 6332 13806 6354
rect 13754 6302 13763 6332
rect 13763 6302 13797 6332
rect 13797 6302 13806 6332
rect 13754 6260 13806 6290
rect 13754 6238 13763 6260
rect 13763 6238 13797 6260
rect 13797 6238 13806 6260
rect 13840 6154 13849 6176
rect 13849 6154 13883 6176
rect 13883 6154 13892 6176
rect 13840 6124 13892 6154
rect 13840 6082 13849 6112
rect 13849 6082 13883 6112
rect 13883 6082 13892 6112
rect 13840 6060 13892 6082
rect 13693 5890 13867 5950
rect 14114 6381 14184 6398
rect 14114 5984 14130 6381
rect 14130 5984 14168 6381
rect 14168 5984 14184 6381
rect 14114 5966 14184 5984
rect 22576 6381 22646 6398
rect 22576 5984 22592 6381
rect 22592 5984 22630 6381
rect 22630 5984 22646 6381
rect 22576 5966 22646 5984
rect 22868 6154 22877 6176
rect 22877 6154 22911 6176
rect 22911 6154 22920 6176
rect 22868 6124 22920 6154
rect 22868 6082 22877 6112
rect 22877 6082 22911 6112
rect 22911 6082 22920 6112
rect 22868 6060 22920 6082
rect 22954 6332 23006 6354
rect 22954 6302 22963 6332
rect 22963 6302 22997 6332
rect 22997 6302 23006 6332
rect 22954 6260 23006 6290
rect 22954 6238 22963 6260
rect 22963 6238 22997 6260
rect 22997 6238 23006 6260
rect 23040 6154 23049 6176
rect 23049 6154 23083 6176
rect 23083 6154 23092 6176
rect 23040 6124 23092 6154
rect 23040 6082 23049 6112
rect 23049 6082 23083 6112
rect 23083 6082 23092 6112
rect 23040 6060 23092 6082
rect 22893 5890 23067 5950
rect 23314 6381 23384 6398
rect 23314 5984 23330 6381
rect 23330 5984 23368 6381
rect 23368 5984 23384 6381
rect 23314 5966 23384 5984
rect 31776 6381 31846 6398
rect 31776 5984 31792 6381
rect 31792 5984 31830 6381
rect 31830 5984 31846 6381
rect 31776 5966 31846 5984
rect 32068 6154 32077 6176
rect 32077 6154 32111 6176
rect 32111 6154 32120 6176
rect 32068 6124 32120 6154
rect 32068 6082 32077 6112
rect 32077 6082 32111 6112
rect 32111 6082 32120 6112
rect 32068 6060 32120 6082
rect 32154 6332 32206 6354
rect 32154 6302 32163 6332
rect 32163 6302 32197 6332
rect 32197 6302 32206 6332
rect 32154 6260 32206 6290
rect 32154 6238 32163 6260
rect 32163 6238 32197 6260
rect 32197 6238 32206 6260
rect 32240 6154 32249 6176
rect 32249 6154 32283 6176
rect 32283 6154 32292 6176
rect 32240 6124 32292 6154
rect 32240 6082 32249 6112
rect 32249 6082 32283 6112
rect 32283 6082 32292 6112
rect 32240 6060 32292 6082
rect 32093 5890 32267 5950
rect 32514 6381 32584 6398
rect 32514 5984 32530 6381
rect 32530 5984 32568 6381
rect 32568 5984 32584 6381
rect 32514 5966 32584 5984
rect 40976 6381 41046 6398
rect 40976 5984 40992 6381
rect 40992 5984 41030 6381
rect 41030 5984 41046 6381
rect 40976 5966 41046 5984
rect 41268 6154 41277 6176
rect 41277 6154 41311 6176
rect 41311 6154 41320 6176
rect 41268 6124 41320 6154
rect 41268 6082 41277 6112
rect 41277 6082 41311 6112
rect 41311 6082 41320 6112
rect 41268 6060 41320 6082
rect 41354 6332 41406 6354
rect 41354 6302 41363 6332
rect 41363 6302 41397 6332
rect 41397 6302 41406 6332
rect 41354 6260 41406 6290
rect 41354 6238 41363 6260
rect 41363 6238 41397 6260
rect 41397 6238 41406 6260
rect 41440 6154 41449 6176
rect 41449 6154 41483 6176
rect 41483 6154 41492 6176
rect 41440 6124 41492 6154
rect 41440 6082 41449 6112
rect 41449 6082 41483 6112
rect 41483 6082 41492 6112
rect 41440 6060 41492 6082
rect 41293 5890 41467 5950
rect 41714 6381 41784 6398
rect 41714 5984 41730 6381
rect 41730 5984 41768 6381
rect 41768 5984 41784 6381
rect 41714 5966 41784 5984
rect 50176 6381 50246 6398
rect 50176 5984 50192 6381
rect 50192 5984 50230 6381
rect 50230 5984 50246 6381
rect 50176 5966 50246 5984
rect 50468 6154 50477 6176
rect 50477 6154 50511 6176
rect 50511 6154 50520 6176
rect 50468 6124 50520 6154
rect 50468 6082 50477 6112
rect 50477 6082 50511 6112
rect 50511 6082 50520 6112
rect 50468 6060 50520 6082
rect 50554 6332 50606 6354
rect 50554 6302 50563 6332
rect 50563 6302 50597 6332
rect 50597 6302 50606 6332
rect 50554 6260 50606 6290
rect 50554 6238 50563 6260
rect 50563 6238 50597 6260
rect 50597 6238 50606 6260
rect 50640 6154 50649 6176
rect 50649 6154 50683 6176
rect 50683 6154 50692 6176
rect 50640 6124 50692 6154
rect 50640 6082 50649 6112
rect 50649 6082 50683 6112
rect 50683 6082 50692 6112
rect 50640 6060 50692 6082
rect 50493 5890 50667 5950
rect 50914 6381 50984 6398
rect 50914 5984 50930 6381
rect 50930 5984 50968 6381
rect 50968 5984 50984 6381
rect 50914 5966 50984 5984
rect 59376 6381 59446 6398
rect 59376 5984 59392 6381
rect 59392 5984 59430 6381
rect 59430 5984 59446 6381
rect 59376 5966 59446 5984
rect 59668 6154 59677 6176
rect 59677 6154 59711 6176
rect 59711 6154 59720 6176
rect 59668 6124 59720 6154
rect 59668 6082 59677 6112
rect 59677 6082 59711 6112
rect 59711 6082 59720 6112
rect 59668 6060 59720 6082
rect 59754 6332 59806 6354
rect 59754 6302 59763 6332
rect 59763 6302 59797 6332
rect 59797 6302 59806 6332
rect 59754 6260 59806 6290
rect 59754 6238 59763 6260
rect 59763 6238 59797 6260
rect 59797 6238 59806 6260
rect 59840 6154 59849 6176
rect 59849 6154 59883 6176
rect 59883 6154 59892 6176
rect 59840 6124 59892 6154
rect 59840 6082 59849 6112
rect 59849 6082 59883 6112
rect 59883 6082 59892 6112
rect 59840 6060 59892 6082
rect 59693 5890 59867 5950
rect 60114 6381 60184 6398
rect 60114 5984 60130 6381
rect 60130 5984 60168 6381
rect 60168 5984 60184 6381
rect 60114 5966 60184 5984
rect 68576 6381 68646 6398
rect 68576 5984 68592 6381
rect 68592 5984 68630 6381
rect 68630 5984 68646 6381
rect 68576 5966 68646 5984
rect 68868 6154 68877 6176
rect 68877 6154 68911 6176
rect 68911 6154 68920 6176
rect 68868 6124 68920 6154
rect 68868 6082 68877 6112
rect 68877 6082 68911 6112
rect 68911 6082 68920 6112
rect 68868 6060 68920 6082
rect 68954 6332 69006 6354
rect 68954 6302 68963 6332
rect 68963 6302 68997 6332
rect 68997 6302 69006 6332
rect 68954 6260 69006 6290
rect 68954 6238 68963 6260
rect 68963 6238 68997 6260
rect 68997 6238 69006 6260
rect 69040 6154 69049 6176
rect 69049 6154 69083 6176
rect 69083 6154 69092 6176
rect 69040 6124 69092 6154
rect 69040 6082 69049 6112
rect 69049 6082 69083 6112
rect 69083 6082 69092 6112
rect 69040 6060 69092 6082
rect 68893 5890 69067 5950
rect 69314 6381 69384 6398
rect 69314 5984 69330 6381
rect 69330 5984 69368 6381
rect 69368 5984 69384 6381
rect 69314 5966 69384 5984
<< metal2 >>
rect -6880 98790 -4880 110790
rect -6880 95560 -4870 98790
rect -6880 95540 -220 95560
rect -6880 95480 -490 95540
rect -240 95480 -220 95540
rect -6880 95460 -220 95480
rect -6880 85680 -4870 95460
rect 4176 95318 4246 95328
rect 4170 94886 4176 95280
rect 4914 95318 4984 95328
rect 4246 95274 4832 95280
rect 4246 95222 4554 95274
rect 4606 95222 4832 95274
rect 4246 95210 4832 95222
rect 4246 95158 4554 95210
rect 4606 95158 4832 95210
rect 4246 95152 4832 95158
rect 4246 94886 4250 95152
rect 4328 95096 4914 95102
rect 4328 95044 4468 95096
rect 4520 95044 4640 95096
rect 4692 95044 4914 95096
rect 4328 95032 4914 95044
rect 4328 94980 4468 95032
rect 4520 94980 4640 95032
rect 4692 94980 4914 95032
rect 4328 94974 4914 94980
rect -240 94750 0 94760
rect -240 94690 -230 94750
rect -170 94690 0 94750
rect -240 94680 0 94690
rect -160 94410 0 94680
rect 4170 94630 4250 94886
rect 4910 94886 4914 94974
rect 4984 94886 4990 95102
rect 4160 94610 4250 94630
rect 4160 94540 4170 94610
rect 4240 94540 4250 94610
rect 4160 94530 4250 94540
rect 4490 94870 4670 94880
rect 4490 94810 4493 94870
rect 4667 94810 4670 94870
rect 4490 94410 4670 94810
rect 4910 94630 4990 94886
rect 4910 94610 5000 94630
rect 4910 94540 4920 94610
rect 4990 94540 5000 94610
rect 4910 94530 5000 94540
rect -160 92410 82600 94410
rect -6880 85660 -220 85680
rect -6880 85600 -490 85660
rect -240 85600 -220 85660
rect -6880 85580 -220 85600
rect -6880 75800 -4870 85580
rect 4176 85438 4246 85448
rect 4170 85006 4176 85400
rect 4914 85438 4984 85448
rect 4246 85394 4832 85400
rect 4246 85342 4554 85394
rect 4606 85342 4832 85394
rect 4246 85330 4832 85342
rect 4246 85278 4554 85330
rect 4606 85278 4832 85330
rect 4246 85272 4832 85278
rect 4246 85006 4250 85272
rect 4328 85216 4914 85222
rect 4328 85164 4468 85216
rect 4520 85164 4640 85216
rect 4692 85164 4914 85216
rect 4328 85152 4914 85164
rect 4328 85100 4468 85152
rect 4520 85100 4640 85152
rect 4692 85100 4914 85152
rect 4328 85094 4914 85100
rect -240 84870 0 84880
rect -240 84810 -230 84870
rect -170 84810 0 84870
rect -240 84800 0 84810
rect -160 84530 0 84800
rect 4170 84750 4250 85006
rect 4910 85006 4914 85094
rect 13376 85438 13446 85448
rect 4984 85006 4990 85222
rect 4160 84730 4250 84750
rect 4160 84660 4170 84730
rect 4240 84660 4250 84730
rect 4160 84650 4250 84660
rect 4490 84990 4670 85000
rect 4490 84930 4493 84990
rect 4667 84930 4670 84990
rect 4490 84530 4670 84930
rect 4910 84750 4990 85006
rect 13370 85006 13376 85400
rect 14114 85438 14184 85448
rect 13446 85394 14032 85400
rect 13446 85342 13754 85394
rect 13806 85342 14032 85394
rect 13446 85330 14032 85342
rect 13446 85278 13754 85330
rect 13806 85278 14032 85330
rect 13446 85272 14032 85278
rect 13446 85006 13450 85272
rect 13528 85216 14114 85222
rect 13528 85164 13668 85216
rect 13720 85164 13840 85216
rect 13892 85164 14114 85216
rect 13528 85152 14114 85164
rect 13528 85100 13668 85152
rect 13720 85100 13840 85152
rect 13892 85100 14114 85152
rect 13528 85094 14114 85100
rect 13370 84750 13450 85006
rect 14110 85006 14114 85094
rect 14184 85006 14190 85222
rect 4910 84730 5000 84750
rect 4910 84660 4920 84730
rect 4990 84660 5000 84730
rect 4910 84650 5000 84660
rect 13360 84730 13450 84750
rect 13360 84660 13370 84730
rect 13440 84660 13450 84730
rect 13360 84650 13450 84660
rect 13690 84990 13870 85000
rect 13690 84930 13693 84990
rect 13867 84930 13870 84990
rect 13690 84530 13870 84930
rect 14110 84750 14190 85006
rect 14110 84730 14200 84750
rect 14110 84660 14120 84730
rect 14190 84660 14200 84730
rect 14110 84650 14200 84660
rect -160 82530 82600 84530
rect -6880 75780 -220 75800
rect -6880 75720 -490 75780
rect -240 75720 -220 75780
rect -6880 75700 -220 75720
rect -6880 65920 -4870 75700
rect 4176 75558 4246 75568
rect 4170 75126 4176 75520
rect 4914 75558 4984 75568
rect 4246 75514 4832 75520
rect 4246 75462 4554 75514
rect 4606 75462 4832 75514
rect 4246 75450 4832 75462
rect 4246 75398 4554 75450
rect 4606 75398 4832 75450
rect 4246 75392 4832 75398
rect 4246 75126 4250 75392
rect 4328 75336 4914 75342
rect 4328 75284 4468 75336
rect 4520 75284 4640 75336
rect 4692 75284 4914 75336
rect 4328 75272 4914 75284
rect 4328 75220 4468 75272
rect 4520 75220 4640 75272
rect 4692 75220 4914 75272
rect 4328 75214 4914 75220
rect -240 74990 0 75000
rect -240 74930 -230 74990
rect -170 74930 0 74990
rect -240 74920 0 74930
rect -160 74650 0 74920
rect 4170 74870 4250 75126
rect 4910 75126 4914 75214
rect 13376 75558 13446 75568
rect 4984 75126 4990 75342
rect 4160 74850 4250 74870
rect 4160 74780 4170 74850
rect 4240 74780 4250 74850
rect 4160 74770 4250 74780
rect 4490 75110 4670 75120
rect 4490 75050 4493 75110
rect 4667 75050 4670 75110
rect 4490 74650 4670 75050
rect 4910 74870 4990 75126
rect 13370 75126 13376 75520
rect 14114 75558 14184 75568
rect 13446 75514 14032 75520
rect 13446 75462 13754 75514
rect 13806 75462 14032 75514
rect 13446 75450 14032 75462
rect 13446 75398 13754 75450
rect 13806 75398 14032 75450
rect 13446 75392 14032 75398
rect 13446 75126 13450 75392
rect 13528 75336 14114 75342
rect 13528 75284 13668 75336
rect 13720 75284 13840 75336
rect 13892 75284 14114 75336
rect 13528 75272 14114 75284
rect 13528 75220 13668 75272
rect 13720 75220 13840 75272
rect 13892 75220 14114 75272
rect 13528 75214 14114 75220
rect 13370 74870 13450 75126
rect 14110 75126 14114 75214
rect 22576 75558 22646 75568
rect 14184 75126 14190 75342
rect 4910 74850 5000 74870
rect 4910 74780 4920 74850
rect 4990 74780 5000 74850
rect 4910 74770 5000 74780
rect 13360 74850 13450 74870
rect 13360 74780 13370 74850
rect 13440 74780 13450 74850
rect 13360 74770 13450 74780
rect 13690 75110 13870 75120
rect 13690 75050 13693 75110
rect 13867 75050 13870 75110
rect 13690 74650 13870 75050
rect 14110 74870 14190 75126
rect 22570 75126 22576 75520
rect 23314 75558 23384 75568
rect 22646 75514 23232 75520
rect 22646 75462 22954 75514
rect 23006 75462 23232 75514
rect 22646 75450 23232 75462
rect 22646 75398 22954 75450
rect 23006 75398 23232 75450
rect 22646 75392 23232 75398
rect 22646 75126 22650 75392
rect 22728 75336 23314 75342
rect 22728 75284 22868 75336
rect 22920 75284 23040 75336
rect 23092 75284 23314 75336
rect 22728 75272 23314 75284
rect 22728 75220 22868 75272
rect 22920 75220 23040 75272
rect 23092 75220 23314 75272
rect 22728 75214 23314 75220
rect 22570 74870 22650 75126
rect 23310 75126 23314 75214
rect 31776 75558 31846 75568
rect 23384 75126 23390 75342
rect 14110 74850 14200 74870
rect 14110 74780 14120 74850
rect 14190 74780 14200 74850
rect 14110 74770 14200 74780
rect 22560 74850 22650 74870
rect 22560 74780 22570 74850
rect 22640 74780 22650 74850
rect 22560 74770 22650 74780
rect 22890 75110 23070 75120
rect 22890 75050 22893 75110
rect 23067 75050 23070 75110
rect 22890 74650 23070 75050
rect 23310 74870 23390 75126
rect 31770 75126 31776 75520
rect 32514 75558 32584 75568
rect 31846 75514 32432 75520
rect 31846 75462 32154 75514
rect 32206 75462 32432 75514
rect 31846 75450 32432 75462
rect 31846 75398 32154 75450
rect 32206 75398 32432 75450
rect 31846 75392 32432 75398
rect 31846 75126 31850 75392
rect 31928 75336 32514 75342
rect 31928 75284 32068 75336
rect 32120 75284 32240 75336
rect 32292 75284 32514 75336
rect 31928 75272 32514 75284
rect 31928 75220 32068 75272
rect 32120 75220 32240 75272
rect 32292 75220 32514 75272
rect 31928 75214 32514 75220
rect 31770 74870 31850 75126
rect 32510 75126 32514 75214
rect 32584 75126 32590 75342
rect 23310 74850 23400 74870
rect 23310 74780 23320 74850
rect 23390 74780 23400 74850
rect 23310 74770 23400 74780
rect 31760 74850 31850 74870
rect 31760 74780 31770 74850
rect 31840 74780 31850 74850
rect 31760 74770 31850 74780
rect 32090 75110 32270 75120
rect 32090 75050 32093 75110
rect 32267 75050 32270 75110
rect 32090 74650 32270 75050
rect 32510 74870 32590 75126
rect 32510 74850 32600 74870
rect 32510 74780 32520 74850
rect 32590 74780 32600 74850
rect 32510 74770 32600 74780
rect -160 72650 82600 74650
rect -6880 65900 -220 65920
rect -6880 65840 -490 65900
rect -240 65840 -220 65900
rect -6880 65820 -220 65840
rect -6880 46160 -4870 65820
rect 4176 65678 4246 65688
rect 4170 65246 4176 65640
rect 4914 65678 4984 65688
rect 4246 65634 4832 65640
rect 4246 65582 4554 65634
rect 4606 65582 4832 65634
rect 4246 65570 4832 65582
rect 4246 65518 4554 65570
rect 4606 65518 4832 65570
rect 4246 65512 4832 65518
rect 4246 65246 4250 65512
rect 4328 65456 4914 65462
rect 4328 65404 4468 65456
rect 4520 65404 4640 65456
rect 4692 65404 4914 65456
rect 4328 65392 4914 65404
rect 4328 65340 4468 65392
rect 4520 65340 4640 65392
rect 4692 65340 4914 65392
rect 4328 65334 4914 65340
rect -240 65110 0 65120
rect -240 65050 -230 65110
rect -170 65050 0 65110
rect -240 65040 0 65050
rect -160 64770 0 65040
rect 4170 64990 4250 65246
rect 4910 65246 4914 65334
rect 13376 65678 13446 65688
rect 4984 65246 4990 65462
rect 4160 64970 4250 64990
rect 4160 64900 4170 64970
rect 4240 64900 4250 64970
rect 4160 64890 4250 64900
rect 4490 65230 4670 65240
rect 4490 65170 4493 65230
rect 4667 65170 4670 65230
rect 4490 64770 4670 65170
rect 4910 64990 4990 65246
rect 13370 65246 13376 65640
rect 14114 65678 14184 65688
rect 13446 65634 14032 65640
rect 13446 65582 13754 65634
rect 13806 65582 14032 65634
rect 13446 65570 14032 65582
rect 13446 65518 13754 65570
rect 13806 65518 14032 65570
rect 13446 65512 14032 65518
rect 13446 65246 13450 65512
rect 13528 65456 14114 65462
rect 13528 65404 13668 65456
rect 13720 65404 13840 65456
rect 13892 65404 14114 65456
rect 13528 65392 14114 65404
rect 13528 65340 13668 65392
rect 13720 65340 13840 65392
rect 13892 65340 14114 65392
rect 13528 65334 14114 65340
rect 13370 64990 13450 65246
rect 14110 65246 14114 65334
rect 22576 65678 22646 65688
rect 14184 65246 14190 65462
rect 4910 64970 5000 64990
rect 4910 64900 4920 64970
rect 4990 64900 5000 64970
rect 4910 64890 5000 64900
rect 13360 64970 13450 64990
rect 13360 64900 13370 64970
rect 13440 64900 13450 64970
rect 13360 64890 13450 64900
rect 13690 65230 13870 65240
rect 13690 65170 13693 65230
rect 13867 65170 13870 65230
rect 13690 64770 13870 65170
rect 14110 64990 14190 65246
rect 22570 65246 22576 65640
rect 23314 65678 23384 65688
rect 22646 65634 23232 65640
rect 22646 65582 22954 65634
rect 23006 65582 23232 65634
rect 22646 65570 23232 65582
rect 22646 65518 22954 65570
rect 23006 65518 23232 65570
rect 22646 65512 23232 65518
rect 22646 65246 22650 65512
rect 22728 65456 23314 65462
rect 22728 65404 22868 65456
rect 22920 65404 23040 65456
rect 23092 65404 23314 65456
rect 22728 65392 23314 65404
rect 22728 65340 22868 65392
rect 22920 65340 23040 65392
rect 23092 65340 23314 65392
rect 22728 65334 23314 65340
rect 22570 64990 22650 65246
rect 23310 65246 23314 65334
rect 31776 65678 31846 65688
rect 23384 65246 23390 65462
rect 14110 64970 14200 64990
rect 14110 64900 14120 64970
rect 14190 64900 14200 64970
rect 14110 64890 14200 64900
rect 22560 64970 22650 64990
rect 22560 64900 22570 64970
rect 22640 64900 22650 64970
rect 22560 64890 22650 64900
rect 22890 65230 23070 65240
rect 22890 65170 22893 65230
rect 23067 65170 23070 65230
rect 22890 64770 23070 65170
rect 23310 64990 23390 65246
rect 31770 65246 31776 65640
rect 32514 65678 32584 65688
rect 31846 65634 32432 65640
rect 31846 65582 32154 65634
rect 32206 65582 32432 65634
rect 31846 65570 32432 65582
rect 31846 65518 32154 65570
rect 32206 65518 32432 65570
rect 31846 65512 32432 65518
rect 31846 65246 31850 65512
rect 31928 65456 32514 65462
rect 31928 65404 32068 65456
rect 32120 65404 32240 65456
rect 32292 65404 32514 65456
rect 31928 65392 32514 65404
rect 31928 65340 32068 65392
rect 32120 65340 32240 65392
rect 32292 65340 32514 65392
rect 31928 65334 32514 65340
rect 31770 64990 31850 65246
rect 32510 65246 32514 65334
rect 40976 65678 41046 65688
rect 32584 65246 32590 65462
rect 23310 64970 23400 64990
rect 23310 64900 23320 64970
rect 23390 64900 23400 64970
rect 23310 64890 23400 64900
rect 31760 64970 31850 64990
rect 31760 64900 31770 64970
rect 31840 64900 31850 64970
rect 31760 64890 31850 64900
rect 32090 65230 32270 65240
rect 32090 65170 32093 65230
rect 32267 65170 32270 65230
rect 32090 64770 32270 65170
rect 32510 64990 32590 65246
rect 40970 65246 40976 65640
rect 41714 65678 41784 65688
rect 41046 65634 41632 65640
rect 41046 65582 41354 65634
rect 41406 65582 41632 65634
rect 41046 65570 41632 65582
rect 41046 65518 41354 65570
rect 41406 65518 41632 65570
rect 41046 65512 41632 65518
rect 41046 65246 41050 65512
rect 41128 65456 41714 65462
rect 41128 65404 41268 65456
rect 41320 65404 41440 65456
rect 41492 65404 41714 65456
rect 41128 65392 41714 65404
rect 41128 65340 41268 65392
rect 41320 65340 41440 65392
rect 41492 65340 41714 65392
rect 41128 65334 41714 65340
rect 40970 64990 41050 65246
rect 41710 65246 41714 65334
rect 50176 65678 50246 65688
rect 41784 65246 41790 65462
rect 32510 64970 32600 64990
rect 32510 64900 32520 64970
rect 32590 64900 32600 64970
rect 32510 64890 32600 64900
rect 40960 64970 41050 64990
rect 40960 64900 40970 64970
rect 41040 64900 41050 64970
rect 40960 64890 41050 64900
rect 41290 65230 41470 65240
rect 41290 65170 41293 65230
rect 41467 65170 41470 65230
rect 41290 64770 41470 65170
rect 41710 64990 41790 65246
rect 50170 65246 50176 65640
rect 50914 65678 50984 65688
rect 50246 65634 50832 65640
rect 50246 65582 50554 65634
rect 50606 65582 50832 65634
rect 50246 65570 50832 65582
rect 50246 65518 50554 65570
rect 50606 65518 50832 65570
rect 50246 65512 50832 65518
rect 50246 65246 50250 65512
rect 50328 65456 50914 65462
rect 50328 65404 50468 65456
rect 50520 65404 50640 65456
rect 50692 65404 50914 65456
rect 50328 65392 50914 65404
rect 50328 65340 50468 65392
rect 50520 65340 50640 65392
rect 50692 65340 50914 65392
rect 50328 65334 50914 65340
rect 50170 64990 50250 65246
rect 50910 65246 50914 65334
rect 59376 65678 59446 65688
rect 50984 65246 50990 65462
rect 41710 64970 41800 64990
rect 41710 64900 41720 64970
rect 41790 64900 41800 64970
rect 41710 64890 41800 64900
rect 50160 64970 50250 64990
rect 50160 64900 50170 64970
rect 50240 64900 50250 64970
rect 50160 64890 50250 64900
rect 50490 65230 50670 65240
rect 50490 65170 50493 65230
rect 50667 65170 50670 65230
rect 50490 64770 50670 65170
rect 50910 64990 50990 65246
rect 59370 65246 59376 65640
rect 60114 65678 60184 65688
rect 59446 65634 60032 65640
rect 59446 65582 59754 65634
rect 59806 65582 60032 65634
rect 59446 65570 60032 65582
rect 59446 65518 59754 65570
rect 59806 65518 60032 65570
rect 59446 65512 60032 65518
rect 59446 65246 59450 65512
rect 59528 65456 60114 65462
rect 59528 65404 59668 65456
rect 59720 65404 59840 65456
rect 59892 65404 60114 65456
rect 59528 65392 60114 65404
rect 59528 65340 59668 65392
rect 59720 65340 59840 65392
rect 59892 65340 60114 65392
rect 59528 65334 60114 65340
rect 59370 64990 59450 65246
rect 60110 65246 60114 65334
rect 68576 65678 68646 65688
rect 60184 65246 60190 65462
rect 50910 64970 51000 64990
rect 50910 64900 50920 64970
rect 50990 64900 51000 64970
rect 50910 64890 51000 64900
rect 59360 64970 59450 64990
rect 59360 64900 59370 64970
rect 59440 64900 59450 64970
rect 59360 64890 59450 64900
rect 59690 65230 59870 65240
rect 59690 65170 59693 65230
rect 59867 65170 59870 65230
rect 59690 64770 59870 65170
rect 60110 64990 60190 65246
rect 68570 65246 68576 65640
rect 69314 65678 69384 65688
rect 68646 65634 69232 65640
rect 68646 65582 68954 65634
rect 69006 65582 69232 65634
rect 68646 65570 69232 65582
rect 68646 65518 68954 65570
rect 69006 65518 69232 65570
rect 68646 65512 69232 65518
rect 68646 65246 68650 65512
rect 68728 65456 69314 65462
rect 68728 65404 68868 65456
rect 68920 65404 69040 65456
rect 69092 65404 69314 65456
rect 68728 65392 69314 65404
rect 68728 65340 68868 65392
rect 68920 65340 69040 65392
rect 69092 65340 69314 65392
rect 68728 65334 69314 65340
rect 68570 64990 68650 65246
rect 69310 65246 69314 65334
rect 69384 65246 69390 65462
rect 60110 64970 60200 64990
rect 60110 64900 60120 64970
rect 60190 64900 60200 64970
rect 60110 64890 60200 64900
rect 68560 64970 68650 64990
rect 68560 64900 68570 64970
rect 68640 64900 68650 64970
rect 68560 64890 68650 64900
rect 68890 65230 69070 65240
rect 68890 65170 68893 65230
rect 69067 65170 69070 65230
rect 68890 64770 69070 65170
rect 69310 64990 69390 65246
rect 69310 64970 69400 64990
rect 69310 64900 69320 64970
rect 69390 64900 69400 64970
rect 69310 64890 69400 64900
rect -160 62770 82600 64770
rect 4176 55798 4246 55808
rect 4170 55366 4176 55760
rect 4914 55798 4984 55808
rect 4246 55754 4832 55760
rect 4246 55702 4554 55754
rect 4606 55702 4832 55754
rect 4246 55690 4832 55702
rect 4246 55638 4554 55690
rect 4606 55638 4832 55690
rect 4246 55632 4832 55638
rect 4246 55366 4250 55632
rect 4328 55576 4914 55582
rect 4328 55524 4468 55576
rect 4520 55524 4640 55576
rect 4692 55524 4914 55576
rect 4328 55512 4914 55524
rect 4328 55460 4468 55512
rect 4520 55460 4640 55512
rect 4692 55460 4914 55512
rect 4328 55454 4914 55460
rect 4170 55110 4250 55366
rect 4910 55366 4914 55454
rect 13376 55798 13446 55808
rect 4984 55366 4990 55582
rect 4160 55090 4250 55110
rect 4160 55020 4170 55090
rect 4240 55020 4250 55090
rect 4160 55010 4250 55020
rect 4490 55350 4670 55360
rect 4490 55290 4493 55350
rect 4667 55290 4670 55350
rect 4490 54890 4670 55290
rect 4910 55110 4990 55366
rect 13370 55366 13376 55760
rect 14114 55798 14184 55808
rect 13446 55754 14032 55760
rect 13446 55702 13754 55754
rect 13806 55702 14032 55754
rect 13446 55690 14032 55702
rect 13446 55638 13754 55690
rect 13806 55638 14032 55690
rect 13446 55632 14032 55638
rect 13446 55366 13450 55632
rect 13528 55576 14114 55582
rect 13528 55524 13668 55576
rect 13720 55524 13840 55576
rect 13892 55524 14114 55576
rect 13528 55512 14114 55524
rect 13528 55460 13668 55512
rect 13720 55460 13840 55512
rect 13892 55460 14114 55512
rect 13528 55454 14114 55460
rect 13370 55110 13450 55366
rect 14110 55366 14114 55454
rect 22576 55798 22646 55808
rect 14184 55366 14190 55582
rect 4910 55090 5000 55110
rect 4910 55020 4920 55090
rect 4990 55020 5000 55090
rect 4910 55010 5000 55020
rect 13360 55090 13450 55110
rect 13360 55020 13370 55090
rect 13440 55020 13450 55090
rect 13360 55010 13450 55020
rect 13690 55350 13870 55360
rect 13690 55290 13693 55350
rect 13867 55290 13870 55350
rect 13690 54890 13870 55290
rect 14110 55110 14190 55366
rect 22570 55366 22576 55760
rect 23314 55798 23384 55808
rect 22646 55754 23232 55760
rect 22646 55702 22954 55754
rect 23006 55702 23232 55754
rect 22646 55690 23232 55702
rect 22646 55638 22954 55690
rect 23006 55638 23232 55690
rect 22646 55632 23232 55638
rect 22646 55366 22650 55632
rect 22728 55576 23314 55582
rect 22728 55524 22868 55576
rect 22920 55524 23040 55576
rect 23092 55524 23314 55576
rect 22728 55512 23314 55524
rect 22728 55460 22868 55512
rect 22920 55460 23040 55512
rect 23092 55460 23314 55512
rect 22728 55454 23314 55460
rect 22570 55110 22650 55366
rect 23310 55366 23314 55454
rect 31776 55798 31846 55808
rect 23384 55366 23390 55582
rect 14110 55090 14200 55110
rect 14110 55020 14120 55090
rect 14190 55020 14200 55090
rect 14110 55010 14200 55020
rect 22560 55090 22650 55110
rect 22560 55020 22570 55090
rect 22640 55020 22650 55090
rect 22560 55010 22650 55020
rect 22890 55350 23070 55360
rect 22890 55290 22893 55350
rect 23067 55290 23070 55350
rect 22890 54890 23070 55290
rect 23310 55110 23390 55366
rect 31770 55366 31776 55760
rect 32514 55798 32584 55808
rect 31846 55754 32432 55760
rect 31846 55702 32154 55754
rect 32206 55702 32432 55754
rect 31846 55690 32432 55702
rect 31846 55638 32154 55690
rect 32206 55638 32432 55690
rect 31846 55632 32432 55638
rect 31846 55366 31850 55632
rect 31928 55576 32514 55582
rect 31928 55524 32068 55576
rect 32120 55524 32240 55576
rect 32292 55524 32514 55576
rect 31928 55512 32514 55524
rect 31928 55460 32068 55512
rect 32120 55460 32240 55512
rect 32292 55460 32514 55512
rect 31928 55454 32514 55460
rect 31770 55110 31850 55366
rect 32510 55366 32514 55454
rect 40976 55798 41046 55808
rect 32584 55366 32590 55582
rect 23310 55090 23400 55110
rect 23310 55020 23320 55090
rect 23390 55020 23400 55090
rect 23310 55010 23400 55020
rect 31760 55090 31850 55110
rect 31760 55020 31770 55090
rect 31840 55020 31850 55090
rect 31760 55010 31850 55020
rect 32090 55350 32270 55360
rect 32090 55290 32093 55350
rect 32267 55290 32270 55350
rect 32090 54890 32270 55290
rect 32510 55110 32590 55366
rect 40970 55366 40976 55760
rect 41714 55798 41784 55808
rect 41046 55754 41632 55760
rect 41046 55702 41354 55754
rect 41406 55702 41632 55754
rect 41046 55690 41632 55702
rect 41046 55638 41354 55690
rect 41406 55638 41632 55690
rect 41046 55632 41632 55638
rect 41046 55366 41050 55632
rect 41128 55576 41714 55582
rect 41128 55524 41268 55576
rect 41320 55524 41440 55576
rect 41492 55524 41714 55576
rect 41128 55512 41714 55524
rect 41128 55460 41268 55512
rect 41320 55460 41440 55512
rect 41492 55460 41714 55512
rect 41128 55454 41714 55460
rect 40970 55110 41050 55366
rect 41710 55366 41714 55454
rect 50176 55798 50246 55808
rect 41784 55366 41790 55582
rect 32510 55090 32600 55110
rect 32510 55020 32520 55090
rect 32590 55020 32600 55090
rect 32510 55010 32600 55020
rect 40960 55090 41050 55110
rect 40960 55020 40970 55090
rect 41040 55020 41050 55090
rect 40960 55010 41050 55020
rect 41290 55350 41470 55360
rect 41290 55290 41293 55350
rect 41467 55290 41470 55350
rect 41290 54890 41470 55290
rect 41710 55110 41790 55366
rect 50170 55366 50176 55760
rect 50914 55798 50984 55808
rect 50246 55754 50832 55760
rect 50246 55702 50554 55754
rect 50606 55702 50832 55754
rect 50246 55690 50832 55702
rect 50246 55638 50554 55690
rect 50606 55638 50832 55690
rect 50246 55632 50832 55638
rect 50246 55366 50250 55632
rect 50328 55576 50914 55582
rect 50328 55524 50468 55576
rect 50520 55524 50640 55576
rect 50692 55524 50914 55576
rect 50328 55512 50914 55524
rect 50328 55460 50468 55512
rect 50520 55460 50640 55512
rect 50692 55460 50914 55512
rect 50328 55454 50914 55460
rect 50170 55110 50250 55366
rect 50910 55366 50914 55454
rect 59376 55798 59446 55808
rect 50984 55366 50990 55582
rect 41710 55090 41800 55110
rect 41710 55020 41720 55090
rect 41790 55020 41800 55090
rect 41710 55010 41800 55020
rect 50160 55090 50250 55110
rect 50160 55020 50170 55090
rect 50240 55020 50250 55090
rect 50160 55010 50250 55020
rect 50490 55350 50670 55360
rect 50490 55290 50493 55350
rect 50667 55290 50670 55350
rect 50490 54890 50670 55290
rect 50910 55110 50990 55366
rect 59370 55366 59376 55760
rect 60114 55798 60184 55808
rect 59446 55754 60032 55760
rect 59446 55702 59754 55754
rect 59806 55702 60032 55754
rect 59446 55690 60032 55702
rect 59446 55638 59754 55690
rect 59806 55638 60032 55690
rect 59446 55632 60032 55638
rect 59446 55366 59450 55632
rect 59528 55576 60114 55582
rect 59528 55524 59668 55576
rect 59720 55524 59840 55576
rect 59892 55524 60114 55576
rect 59528 55512 60114 55524
rect 59528 55460 59668 55512
rect 59720 55460 59840 55512
rect 59892 55460 60114 55512
rect 59528 55454 60114 55460
rect 59370 55110 59450 55366
rect 60110 55366 60114 55454
rect 68576 55798 68646 55808
rect 60184 55366 60190 55582
rect 50910 55090 51000 55110
rect 50910 55020 50920 55090
rect 50990 55020 51000 55090
rect 50910 55010 51000 55020
rect 59360 55090 59450 55110
rect 59360 55020 59370 55090
rect 59440 55020 59450 55090
rect 59360 55010 59450 55020
rect 59690 55350 59870 55360
rect 59690 55290 59693 55350
rect 59867 55290 59870 55350
rect 59690 54890 59870 55290
rect 60110 55110 60190 55366
rect 68570 55366 68576 55760
rect 69314 55798 69384 55808
rect 68646 55754 69232 55760
rect 68646 55702 68954 55754
rect 69006 55702 69232 55754
rect 68646 55690 69232 55702
rect 68646 55638 68954 55690
rect 69006 55638 69232 55690
rect 68646 55632 69232 55638
rect 68646 55366 68650 55632
rect 68728 55576 69314 55582
rect 68728 55524 68868 55576
rect 68920 55524 69040 55576
rect 69092 55524 69314 55576
rect 68728 55512 69314 55524
rect 68728 55460 68868 55512
rect 68920 55460 69040 55512
rect 69092 55460 69314 55512
rect 68728 55454 69314 55460
rect 68570 55110 68650 55366
rect 69310 55366 69314 55454
rect 69384 55366 69390 55582
rect 60110 55090 60200 55110
rect 60110 55020 60120 55090
rect 60190 55020 60200 55090
rect 60110 55010 60200 55020
rect 68560 55090 68650 55110
rect 68560 55020 68570 55090
rect 68640 55020 68650 55090
rect 68560 55010 68650 55020
rect 68890 55350 69070 55360
rect 68890 55290 68893 55350
rect 69067 55290 69070 55350
rect 68890 54890 69070 55290
rect 69310 55110 69390 55366
rect 69310 55090 69400 55110
rect 69310 55020 69320 55090
rect 69390 55020 69400 55090
rect 69310 55010 69400 55020
rect 0 52890 81600 54890
rect -6880 46140 -220 46160
rect -6880 46080 -490 46140
rect -240 46080 -220 46140
rect -6880 46060 -220 46080
rect -6880 6640 -4870 46060
rect 4176 45918 4246 45928
rect 4170 45486 4176 45880
rect 4914 45918 4984 45928
rect 4246 45874 4832 45880
rect 4246 45822 4554 45874
rect 4606 45822 4832 45874
rect 4246 45810 4832 45822
rect 4246 45758 4554 45810
rect 4606 45758 4832 45810
rect 4246 45752 4832 45758
rect 4246 45486 4250 45752
rect 4328 45696 4914 45702
rect 4328 45644 4468 45696
rect 4520 45644 4640 45696
rect 4692 45644 4914 45696
rect 4328 45632 4914 45644
rect 4328 45580 4468 45632
rect 4520 45580 4640 45632
rect 4692 45580 4914 45632
rect 4328 45574 4914 45580
rect -240 45350 0 45360
rect -240 45290 -230 45350
rect -170 45290 0 45350
rect -240 45280 0 45290
rect -160 45010 0 45280
rect 4170 45230 4250 45486
rect 4910 45486 4914 45574
rect 13376 45918 13446 45928
rect 4984 45486 4990 45702
rect 4160 45210 4250 45230
rect 4160 45140 4170 45210
rect 4240 45140 4250 45210
rect 4160 45130 4250 45140
rect 4490 45470 4670 45480
rect 4490 45410 4493 45470
rect 4667 45410 4670 45470
rect 4490 45010 4670 45410
rect 4910 45230 4990 45486
rect 13370 45486 13376 45880
rect 14114 45918 14184 45928
rect 13446 45874 14032 45880
rect 13446 45822 13754 45874
rect 13806 45822 14032 45874
rect 13446 45810 14032 45822
rect 13446 45758 13754 45810
rect 13806 45758 14032 45810
rect 13446 45752 14032 45758
rect 13446 45486 13450 45752
rect 13528 45696 14114 45702
rect 13528 45644 13668 45696
rect 13720 45644 13840 45696
rect 13892 45644 14114 45696
rect 13528 45632 14114 45644
rect 13528 45580 13668 45632
rect 13720 45580 13840 45632
rect 13892 45580 14114 45632
rect 13528 45574 14114 45580
rect 13370 45230 13450 45486
rect 14110 45486 14114 45574
rect 22576 45918 22646 45928
rect 14184 45486 14190 45702
rect 4910 45210 5000 45230
rect 4910 45140 4920 45210
rect 4990 45140 5000 45210
rect 4910 45130 5000 45140
rect 13360 45210 13450 45230
rect 13360 45140 13370 45210
rect 13440 45140 13450 45210
rect 13360 45130 13450 45140
rect 13690 45470 13870 45480
rect 13690 45410 13693 45470
rect 13867 45410 13870 45470
rect 13690 45010 13870 45410
rect 14110 45230 14190 45486
rect 22570 45486 22576 45880
rect 23314 45918 23384 45928
rect 22646 45874 23232 45880
rect 22646 45822 22954 45874
rect 23006 45822 23232 45874
rect 22646 45810 23232 45822
rect 22646 45758 22954 45810
rect 23006 45758 23232 45810
rect 22646 45752 23232 45758
rect 22646 45486 22650 45752
rect 22728 45696 23314 45702
rect 22728 45644 22868 45696
rect 22920 45644 23040 45696
rect 23092 45644 23314 45696
rect 22728 45632 23314 45644
rect 22728 45580 22868 45632
rect 22920 45580 23040 45632
rect 23092 45580 23314 45632
rect 22728 45574 23314 45580
rect 22570 45230 22650 45486
rect 23310 45486 23314 45574
rect 31776 45918 31846 45928
rect 23384 45486 23390 45702
rect 14110 45210 14200 45230
rect 14110 45140 14120 45210
rect 14190 45140 14200 45210
rect 14110 45130 14200 45140
rect 22560 45210 22650 45230
rect 22560 45140 22570 45210
rect 22640 45140 22650 45210
rect 22560 45130 22650 45140
rect 22890 45470 23070 45480
rect 22890 45410 22893 45470
rect 23067 45410 23070 45470
rect 22890 45010 23070 45410
rect 23310 45230 23390 45486
rect 31770 45486 31776 45880
rect 32514 45918 32584 45928
rect 31846 45874 32432 45880
rect 31846 45822 32154 45874
rect 32206 45822 32432 45874
rect 31846 45810 32432 45822
rect 31846 45758 32154 45810
rect 32206 45758 32432 45810
rect 31846 45752 32432 45758
rect 31846 45486 31850 45752
rect 31928 45696 32514 45702
rect 31928 45644 32068 45696
rect 32120 45644 32240 45696
rect 32292 45644 32514 45696
rect 31928 45632 32514 45644
rect 31928 45580 32068 45632
rect 32120 45580 32240 45632
rect 32292 45580 32514 45632
rect 31928 45574 32514 45580
rect 31770 45230 31850 45486
rect 32510 45486 32514 45574
rect 40976 45918 41046 45928
rect 32584 45486 32590 45702
rect 23310 45210 23400 45230
rect 23310 45140 23320 45210
rect 23390 45140 23400 45210
rect 23310 45130 23400 45140
rect 31760 45210 31850 45230
rect 31760 45140 31770 45210
rect 31840 45140 31850 45210
rect 31760 45130 31850 45140
rect 32090 45470 32270 45480
rect 32090 45410 32093 45470
rect 32267 45410 32270 45470
rect 32090 45010 32270 45410
rect 32510 45230 32590 45486
rect 40970 45486 40976 45880
rect 41714 45918 41784 45928
rect 41046 45874 41632 45880
rect 41046 45822 41354 45874
rect 41406 45822 41632 45874
rect 41046 45810 41632 45822
rect 41046 45758 41354 45810
rect 41406 45758 41632 45810
rect 41046 45752 41632 45758
rect 41046 45486 41050 45752
rect 41128 45696 41714 45702
rect 41128 45644 41268 45696
rect 41320 45644 41440 45696
rect 41492 45644 41714 45696
rect 41128 45632 41714 45644
rect 41128 45580 41268 45632
rect 41320 45580 41440 45632
rect 41492 45580 41714 45632
rect 41128 45574 41714 45580
rect 40970 45230 41050 45486
rect 41710 45486 41714 45574
rect 50176 45918 50246 45928
rect 41784 45486 41790 45702
rect 32510 45210 32600 45230
rect 32510 45140 32520 45210
rect 32590 45140 32600 45210
rect 32510 45130 32600 45140
rect 40960 45210 41050 45230
rect 40960 45140 40970 45210
rect 41040 45140 41050 45210
rect 40960 45130 41050 45140
rect 41290 45470 41470 45480
rect 41290 45410 41293 45470
rect 41467 45410 41470 45470
rect 41290 45010 41470 45410
rect 41710 45230 41790 45486
rect 50170 45486 50176 45880
rect 50914 45918 50984 45928
rect 50246 45874 50832 45880
rect 50246 45822 50554 45874
rect 50606 45822 50832 45874
rect 50246 45810 50832 45822
rect 50246 45758 50554 45810
rect 50606 45758 50832 45810
rect 50246 45752 50832 45758
rect 50246 45486 50250 45752
rect 50328 45696 50914 45702
rect 50328 45644 50468 45696
rect 50520 45644 50640 45696
rect 50692 45644 50914 45696
rect 50328 45632 50914 45644
rect 50328 45580 50468 45632
rect 50520 45580 50640 45632
rect 50692 45580 50914 45632
rect 50328 45574 50914 45580
rect 50170 45230 50250 45486
rect 50910 45486 50914 45574
rect 59376 45918 59446 45928
rect 50984 45486 50990 45702
rect 41710 45210 41800 45230
rect 41710 45140 41720 45210
rect 41790 45140 41800 45210
rect 41710 45130 41800 45140
rect 50160 45210 50250 45230
rect 50160 45140 50170 45210
rect 50240 45140 50250 45210
rect 50160 45130 50250 45140
rect 50490 45470 50670 45480
rect 50490 45410 50493 45470
rect 50667 45410 50670 45470
rect 50490 45010 50670 45410
rect 50910 45230 50990 45486
rect 59370 45486 59376 45880
rect 60114 45918 60184 45928
rect 59446 45874 60032 45880
rect 59446 45822 59754 45874
rect 59806 45822 60032 45874
rect 59446 45810 60032 45822
rect 59446 45758 59754 45810
rect 59806 45758 60032 45810
rect 59446 45752 60032 45758
rect 59446 45486 59450 45752
rect 59528 45696 60114 45702
rect 59528 45644 59668 45696
rect 59720 45644 59840 45696
rect 59892 45644 60114 45696
rect 59528 45632 60114 45644
rect 59528 45580 59668 45632
rect 59720 45580 59840 45632
rect 59892 45580 60114 45632
rect 59528 45574 60114 45580
rect 59370 45230 59450 45486
rect 60110 45486 60114 45574
rect 68576 45918 68646 45928
rect 60184 45486 60190 45702
rect 50910 45210 51000 45230
rect 50910 45140 50920 45210
rect 50990 45140 51000 45210
rect 50910 45130 51000 45140
rect 59360 45210 59450 45230
rect 59360 45140 59370 45210
rect 59440 45140 59450 45210
rect 59360 45130 59450 45140
rect 59690 45470 59870 45480
rect 59690 45410 59693 45470
rect 59867 45410 59870 45470
rect 59690 45010 59870 45410
rect 60110 45230 60190 45486
rect 68570 45486 68576 45880
rect 69314 45918 69384 45928
rect 68646 45874 69232 45880
rect 68646 45822 68954 45874
rect 69006 45822 69232 45874
rect 68646 45810 69232 45822
rect 68646 45758 68954 45810
rect 69006 45758 69232 45810
rect 68646 45752 69232 45758
rect 68646 45486 68650 45752
rect 68728 45696 69314 45702
rect 68728 45644 68868 45696
rect 68920 45644 69040 45696
rect 69092 45644 69314 45696
rect 68728 45632 69314 45644
rect 68728 45580 68868 45632
rect 68920 45580 69040 45632
rect 69092 45580 69314 45632
rect 68728 45574 69314 45580
rect 68570 45230 68650 45486
rect 69310 45486 69314 45574
rect 69384 45486 69390 45702
rect 60110 45210 60200 45230
rect 60110 45140 60120 45210
rect 60190 45140 60200 45210
rect 60110 45130 60200 45140
rect 68560 45210 68650 45230
rect 68560 45140 68570 45210
rect 68640 45140 68650 45210
rect 68560 45130 68650 45140
rect 68890 45470 69070 45480
rect 68890 45410 68893 45470
rect 69067 45410 69070 45470
rect 68890 45010 69070 45410
rect 69310 45230 69390 45486
rect 69310 45210 69400 45230
rect 69310 45140 69320 45210
rect 69390 45140 69400 45210
rect 69310 45130 69400 45140
rect 79600 45010 81600 52890
rect -160 43010 82600 45010
rect 4176 36038 4246 36048
rect 4170 35606 4176 36000
rect 4914 36038 4984 36048
rect 4246 35994 4832 36000
rect 4246 35942 4554 35994
rect 4606 35942 4832 35994
rect 4246 35930 4832 35942
rect 4246 35878 4554 35930
rect 4606 35878 4832 35930
rect 4246 35872 4832 35878
rect 4246 35606 4250 35872
rect 4328 35816 4914 35822
rect 4328 35764 4468 35816
rect 4520 35764 4640 35816
rect 4692 35764 4914 35816
rect 4328 35752 4914 35764
rect 4328 35700 4468 35752
rect 4520 35700 4640 35752
rect 4692 35700 4914 35752
rect 4328 35694 4914 35700
rect 4170 35350 4250 35606
rect 4910 35606 4914 35694
rect 13376 36038 13446 36048
rect 4984 35606 4990 35822
rect 4160 35330 4250 35350
rect 4160 35260 4170 35330
rect 4240 35260 4250 35330
rect 4160 35250 4250 35260
rect 4490 35590 4670 35600
rect 4490 35530 4493 35590
rect 4667 35530 4670 35590
rect 4490 35130 4670 35530
rect 4910 35350 4990 35606
rect 13370 35606 13376 36000
rect 14114 36038 14184 36048
rect 13446 35994 14032 36000
rect 13446 35942 13754 35994
rect 13806 35942 14032 35994
rect 13446 35930 14032 35942
rect 13446 35878 13754 35930
rect 13806 35878 14032 35930
rect 13446 35872 14032 35878
rect 13446 35606 13450 35872
rect 13528 35816 14114 35822
rect 13528 35764 13668 35816
rect 13720 35764 13840 35816
rect 13892 35764 14114 35816
rect 13528 35752 14114 35764
rect 13528 35700 13668 35752
rect 13720 35700 13840 35752
rect 13892 35700 14114 35752
rect 13528 35694 14114 35700
rect 13370 35350 13450 35606
rect 14110 35606 14114 35694
rect 22576 36038 22646 36048
rect 14184 35606 14190 35822
rect 4910 35330 5000 35350
rect 4910 35260 4920 35330
rect 4990 35260 5000 35330
rect 4910 35250 5000 35260
rect 13360 35330 13450 35350
rect 13360 35260 13370 35330
rect 13440 35260 13450 35330
rect 13360 35250 13450 35260
rect 13690 35590 13870 35600
rect 13690 35530 13693 35590
rect 13867 35530 13870 35590
rect 13690 35130 13870 35530
rect 14110 35350 14190 35606
rect 22570 35606 22576 36000
rect 23314 36038 23384 36048
rect 22646 35994 23232 36000
rect 22646 35942 22954 35994
rect 23006 35942 23232 35994
rect 22646 35930 23232 35942
rect 22646 35878 22954 35930
rect 23006 35878 23232 35930
rect 22646 35872 23232 35878
rect 22646 35606 22650 35872
rect 22728 35816 23314 35822
rect 22728 35764 22868 35816
rect 22920 35764 23040 35816
rect 23092 35764 23314 35816
rect 22728 35752 23314 35764
rect 22728 35700 22868 35752
rect 22920 35700 23040 35752
rect 23092 35700 23314 35752
rect 22728 35694 23314 35700
rect 22570 35350 22650 35606
rect 23310 35606 23314 35694
rect 31776 36038 31846 36048
rect 23384 35606 23390 35822
rect 14110 35330 14200 35350
rect 14110 35260 14120 35330
rect 14190 35260 14200 35330
rect 14110 35250 14200 35260
rect 22560 35330 22650 35350
rect 22560 35260 22570 35330
rect 22640 35260 22650 35330
rect 22560 35250 22650 35260
rect 22890 35590 23070 35600
rect 22890 35530 22893 35590
rect 23067 35530 23070 35590
rect 22890 35130 23070 35530
rect 23310 35350 23390 35606
rect 31770 35606 31776 36000
rect 32514 36038 32584 36048
rect 31846 35994 32432 36000
rect 31846 35942 32154 35994
rect 32206 35942 32432 35994
rect 31846 35930 32432 35942
rect 31846 35878 32154 35930
rect 32206 35878 32432 35930
rect 31846 35872 32432 35878
rect 31846 35606 31850 35872
rect 31928 35816 32514 35822
rect 31928 35764 32068 35816
rect 32120 35764 32240 35816
rect 32292 35764 32514 35816
rect 31928 35752 32514 35764
rect 31928 35700 32068 35752
rect 32120 35700 32240 35752
rect 32292 35700 32514 35752
rect 31928 35694 32514 35700
rect 31770 35350 31850 35606
rect 32510 35606 32514 35694
rect 40976 36038 41046 36048
rect 32584 35606 32590 35822
rect 23310 35330 23400 35350
rect 23310 35260 23320 35330
rect 23390 35260 23400 35330
rect 23310 35250 23400 35260
rect 31760 35330 31850 35350
rect 31760 35260 31770 35330
rect 31840 35260 31850 35330
rect 31760 35250 31850 35260
rect 32090 35590 32270 35600
rect 32090 35530 32093 35590
rect 32267 35530 32270 35590
rect 32090 35130 32270 35530
rect 32510 35350 32590 35606
rect 40970 35606 40976 36000
rect 41714 36038 41784 36048
rect 41046 35994 41632 36000
rect 41046 35942 41354 35994
rect 41406 35942 41632 35994
rect 41046 35930 41632 35942
rect 41046 35878 41354 35930
rect 41406 35878 41632 35930
rect 41046 35872 41632 35878
rect 41046 35606 41050 35872
rect 41128 35816 41714 35822
rect 41128 35764 41268 35816
rect 41320 35764 41440 35816
rect 41492 35764 41714 35816
rect 41128 35752 41714 35764
rect 41128 35700 41268 35752
rect 41320 35700 41440 35752
rect 41492 35700 41714 35752
rect 41128 35694 41714 35700
rect 40970 35350 41050 35606
rect 41710 35606 41714 35694
rect 50176 36038 50246 36048
rect 41784 35606 41790 35822
rect 32510 35330 32600 35350
rect 32510 35260 32520 35330
rect 32590 35260 32600 35330
rect 32510 35250 32600 35260
rect 40960 35330 41050 35350
rect 40960 35260 40970 35330
rect 41040 35260 41050 35330
rect 40960 35250 41050 35260
rect 41290 35590 41470 35600
rect 41290 35530 41293 35590
rect 41467 35530 41470 35590
rect 41290 35130 41470 35530
rect 41710 35350 41790 35606
rect 50170 35606 50176 36000
rect 50914 36038 50984 36048
rect 50246 35994 50832 36000
rect 50246 35942 50554 35994
rect 50606 35942 50832 35994
rect 50246 35930 50832 35942
rect 50246 35878 50554 35930
rect 50606 35878 50832 35930
rect 50246 35872 50832 35878
rect 50246 35606 50250 35872
rect 50328 35816 50914 35822
rect 50328 35764 50468 35816
rect 50520 35764 50640 35816
rect 50692 35764 50914 35816
rect 50328 35752 50914 35764
rect 50328 35700 50468 35752
rect 50520 35700 50640 35752
rect 50692 35700 50914 35752
rect 50328 35694 50914 35700
rect 50170 35350 50250 35606
rect 50910 35606 50914 35694
rect 59376 36038 59446 36048
rect 50984 35606 50990 35822
rect 41710 35330 41800 35350
rect 41710 35260 41720 35330
rect 41790 35260 41800 35330
rect 41710 35250 41800 35260
rect 50160 35330 50250 35350
rect 50160 35260 50170 35330
rect 50240 35260 50250 35330
rect 50160 35250 50250 35260
rect 50490 35590 50670 35600
rect 50490 35530 50493 35590
rect 50667 35530 50670 35590
rect 50490 35130 50670 35530
rect 50910 35350 50990 35606
rect 59370 35606 59376 36000
rect 60114 36038 60184 36048
rect 59446 35994 60032 36000
rect 59446 35942 59754 35994
rect 59806 35942 60032 35994
rect 59446 35930 60032 35942
rect 59446 35878 59754 35930
rect 59806 35878 60032 35930
rect 59446 35872 60032 35878
rect 59446 35606 59450 35872
rect 59528 35816 60114 35822
rect 59528 35764 59668 35816
rect 59720 35764 59840 35816
rect 59892 35764 60114 35816
rect 59528 35752 60114 35764
rect 59528 35700 59668 35752
rect 59720 35700 59840 35752
rect 59892 35700 60114 35752
rect 59528 35694 60114 35700
rect 59370 35350 59450 35606
rect 60110 35606 60114 35694
rect 68576 36038 68646 36048
rect 60184 35606 60190 35822
rect 50910 35330 51000 35350
rect 50910 35260 50920 35330
rect 50990 35260 51000 35330
rect 50910 35250 51000 35260
rect 59360 35330 59450 35350
rect 59360 35260 59370 35330
rect 59440 35260 59450 35330
rect 59360 35250 59450 35260
rect 59690 35590 59870 35600
rect 59690 35530 59693 35590
rect 59867 35530 59870 35590
rect 59690 35130 59870 35530
rect 60110 35350 60190 35606
rect 68570 35606 68576 36000
rect 69314 36038 69384 36048
rect 68646 35994 69232 36000
rect 68646 35942 68954 35994
rect 69006 35942 69232 35994
rect 68646 35930 69232 35942
rect 68646 35878 68954 35930
rect 69006 35878 69232 35930
rect 68646 35872 69232 35878
rect 68646 35606 68650 35872
rect 68728 35816 69314 35822
rect 68728 35764 68868 35816
rect 68920 35764 69040 35816
rect 69092 35764 69314 35816
rect 68728 35752 69314 35764
rect 68728 35700 68868 35752
rect 68920 35700 69040 35752
rect 69092 35700 69314 35752
rect 68728 35694 69314 35700
rect 68570 35350 68650 35606
rect 69310 35606 69314 35694
rect 69384 35606 69390 35822
rect 60110 35330 60200 35350
rect 60110 35260 60120 35330
rect 60190 35260 60200 35330
rect 60110 35250 60200 35260
rect 68560 35330 68650 35350
rect 68560 35260 68570 35330
rect 68640 35260 68650 35330
rect 68560 35250 68650 35260
rect 68890 35590 69070 35600
rect 68890 35530 68893 35590
rect 69067 35530 69070 35590
rect 68890 35130 69070 35530
rect 69310 35350 69390 35606
rect 69310 35330 69400 35350
rect 69310 35260 69320 35330
rect 69390 35260 69400 35330
rect 69310 35250 69400 35260
rect 0 33130 81600 35130
rect 4176 26158 4246 26168
rect 4170 25726 4176 26120
rect 4914 26158 4984 26168
rect 4246 26114 4832 26120
rect 4246 26062 4554 26114
rect 4606 26062 4832 26114
rect 4246 26050 4832 26062
rect 4246 25998 4554 26050
rect 4606 25998 4832 26050
rect 4246 25992 4832 25998
rect 4246 25726 4250 25992
rect 4328 25936 4914 25942
rect 4328 25884 4468 25936
rect 4520 25884 4640 25936
rect 4692 25884 4914 25936
rect 4328 25872 4914 25884
rect 4328 25820 4468 25872
rect 4520 25820 4640 25872
rect 4692 25820 4914 25872
rect 4328 25814 4914 25820
rect 4170 25470 4250 25726
rect 4910 25726 4914 25814
rect 13376 26158 13446 26168
rect 4984 25726 4990 25942
rect 4160 25450 4250 25470
rect 4160 25380 4170 25450
rect 4240 25380 4250 25450
rect 4160 25370 4250 25380
rect 4490 25710 4670 25720
rect 4490 25650 4493 25710
rect 4667 25650 4670 25710
rect 4490 25250 4670 25650
rect 4910 25470 4990 25726
rect 13370 25726 13376 26120
rect 14114 26158 14184 26168
rect 13446 26114 14032 26120
rect 13446 26062 13754 26114
rect 13806 26062 14032 26114
rect 13446 26050 14032 26062
rect 13446 25998 13754 26050
rect 13806 25998 14032 26050
rect 13446 25992 14032 25998
rect 13446 25726 13450 25992
rect 13528 25936 14114 25942
rect 13528 25884 13668 25936
rect 13720 25884 13840 25936
rect 13892 25884 14114 25936
rect 13528 25872 14114 25884
rect 13528 25820 13668 25872
rect 13720 25820 13840 25872
rect 13892 25820 14114 25872
rect 13528 25814 14114 25820
rect 13370 25470 13450 25726
rect 14110 25726 14114 25814
rect 22576 26158 22646 26168
rect 14184 25726 14190 25942
rect 4910 25450 5000 25470
rect 4910 25380 4920 25450
rect 4990 25380 5000 25450
rect 4910 25370 5000 25380
rect 13360 25450 13450 25470
rect 13360 25380 13370 25450
rect 13440 25380 13450 25450
rect 13360 25370 13450 25380
rect 13690 25710 13870 25720
rect 13690 25650 13693 25710
rect 13867 25650 13870 25710
rect 13690 25250 13870 25650
rect 14110 25470 14190 25726
rect 22570 25726 22576 26120
rect 23314 26158 23384 26168
rect 22646 26114 23232 26120
rect 22646 26062 22954 26114
rect 23006 26062 23232 26114
rect 22646 26050 23232 26062
rect 22646 25998 22954 26050
rect 23006 25998 23232 26050
rect 22646 25992 23232 25998
rect 22646 25726 22650 25992
rect 22728 25936 23314 25942
rect 22728 25884 22868 25936
rect 22920 25884 23040 25936
rect 23092 25884 23314 25936
rect 22728 25872 23314 25884
rect 22728 25820 22868 25872
rect 22920 25820 23040 25872
rect 23092 25820 23314 25872
rect 22728 25814 23314 25820
rect 22570 25470 22650 25726
rect 23310 25726 23314 25814
rect 31776 26158 31846 26168
rect 23384 25726 23390 25942
rect 14110 25450 14200 25470
rect 14110 25380 14120 25450
rect 14190 25380 14200 25450
rect 14110 25370 14200 25380
rect 22560 25450 22650 25470
rect 22560 25380 22570 25450
rect 22640 25380 22650 25450
rect 22560 25370 22650 25380
rect 22890 25710 23070 25720
rect 22890 25650 22893 25710
rect 23067 25650 23070 25710
rect 22890 25250 23070 25650
rect 23310 25470 23390 25726
rect 31770 25726 31776 26120
rect 32514 26158 32584 26168
rect 31846 26114 32432 26120
rect 31846 26062 32154 26114
rect 32206 26062 32432 26114
rect 31846 26050 32432 26062
rect 31846 25998 32154 26050
rect 32206 25998 32432 26050
rect 31846 25992 32432 25998
rect 31846 25726 31850 25992
rect 31928 25936 32514 25942
rect 31928 25884 32068 25936
rect 32120 25884 32240 25936
rect 32292 25884 32514 25936
rect 31928 25872 32514 25884
rect 31928 25820 32068 25872
rect 32120 25820 32240 25872
rect 32292 25820 32514 25872
rect 31928 25814 32514 25820
rect 31770 25470 31850 25726
rect 32510 25726 32514 25814
rect 40976 26158 41046 26168
rect 32584 25726 32590 25942
rect 23310 25450 23400 25470
rect 23310 25380 23320 25450
rect 23390 25380 23400 25450
rect 23310 25370 23400 25380
rect 31760 25450 31850 25470
rect 31760 25380 31770 25450
rect 31840 25380 31850 25450
rect 31760 25370 31850 25380
rect 32090 25710 32270 25720
rect 32090 25650 32093 25710
rect 32267 25650 32270 25710
rect 32090 25250 32270 25650
rect 32510 25470 32590 25726
rect 40970 25726 40976 26120
rect 41714 26158 41784 26168
rect 41046 26114 41632 26120
rect 41046 26062 41354 26114
rect 41406 26062 41632 26114
rect 41046 26050 41632 26062
rect 41046 25998 41354 26050
rect 41406 25998 41632 26050
rect 41046 25992 41632 25998
rect 41046 25726 41050 25992
rect 41128 25936 41714 25942
rect 41128 25884 41268 25936
rect 41320 25884 41440 25936
rect 41492 25884 41714 25936
rect 41128 25872 41714 25884
rect 41128 25820 41268 25872
rect 41320 25820 41440 25872
rect 41492 25820 41714 25872
rect 41128 25814 41714 25820
rect 40970 25470 41050 25726
rect 41710 25726 41714 25814
rect 50176 26158 50246 26168
rect 41784 25726 41790 25942
rect 32510 25450 32600 25470
rect 32510 25380 32520 25450
rect 32590 25380 32600 25450
rect 32510 25370 32600 25380
rect 40960 25450 41050 25470
rect 40960 25380 40970 25450
rect 41040 25380 41050 25450
rect 40960 25370 41050 25380
rect 41290 25710 41470 25720
rect 41290 25650 41293 25710
rect 41467 25650 41470 25710
rect 41290 25250 41470 25650
rect 41710 25470 41790 25726
rect 50170 25726 50176 26120
rect 50914 26158 50984 26168
rect 50246 26114 50832 26120
rect 50246 26062 50554 26114
rect 50606 26062 50832 26114
rect 50246 26050 50832 26062
rect 50246 25998 50554 26050
rect 50606 25998 50832 26050
rect 50246 25992 50832 25998
rect 50246 25726 50250 25992
rect 50328 25936 50914 25942
rect 50328 25884 50468 25936
rect 50520 25884 50640 25936
rect 50692 25884 50914 25936
rect 50328 25872 50914 25884
rect 50328 25820 50468 25872
rect 50520 25820 50640 25872
rect 50692 25820 50914 25872
rect 50328 25814 50914 25820
rect 50170 25470 50250 25726
rect 50910 25726 50914 25814
rect 59376 26158 59446 26168
rect 50984 25726 50990 25942
rect 41710 25450 41800 25470
rect 41710 25380 41720 25450
rect 41790 25380 41800 25450
rect 41710 25370 41800 25380
rect 50160 25450 50250 25470
rect 50160 25380 50170 25450
rect 50240 25380 50250 25450
rect 50160 25370 50250 25380
rect 50490 25710 50670 25720
rect 50490 25650 50493 25710
rect 50667 25650 50670 25710
rect 50490 25250 50670 25650
rect 50910 25470 50990 25726
rect 59370 25726 59376 26120
rect 60114 26158 60184 26168
rect 59446 26114 60032 26120
rect 59446 26062 59754 26114
rect 59806 26062 60032 26114
rect 59446 26050 60032 26062
rect 59446 25998 59754 26050
rect 59806 25998 60032 26050
rect 59446 25992 60032 25998
rect 59446 25726 59450 25992
rect 59528 25936 60114 25942
rect 59528 25884 59668 25936
rect 59720 25884 59840 25936
rect 59892 25884 60114 25936
rect 59528 25872 60114 25884
rect 59528 25820 59668 25872
rect 59720 25820 59840 25872
rect 59892 25820 60114 25872
rect 59528 25814 60114 25820
rect 59370 25470 59450 25726
rect 60110 25726 60114 25814
rect 68576 26158 68646 26168
rect 60184 25726 60190 25942
rect 50910 25450 51000 25470
rect 50910 25380 50920 25450
rect 50990 25380 51000 25450
rect 50910 25370 51000 25380
rect 59360 25450 59450 25470
rect 59360 25380 59370 25450
rect 59440 25380 59450 25450
rect 59360 25370 59450 25380
rect 59690 25710 59870 25720
rect 59690 25650 59693 25710
rect 59867 25650 59870 25710
rect 59690 25250 59870 25650
rect 60110 25470 60190 25726
rect 68570 25726 68576 26120
rect 69314 26158 69384 26168
rect 68646 26114 69232 26120
rect 68646 26062 68954 26114
rect 69006 26062 69232 26114
rect 68646 26050 69232 26062
rect 68646 25998 68954 26050
rect 69006 25998 69232 26050
rect 68646 25992 69232 25998
rect 68646 25726 68650 25992
rect 68728 25936 69314 25942
rect 68728 25884 68868 25936
rect 68920 25884 69040 25936
rect 69092 25884 69314 25936
rect 68728 25872 69314 25884
rect 68728 25820 68868 25872
rect 68920 25820 69040 25872
rect 69092 25820 69314 25872
rect 68728 25814 69314 25820
rect 68570 25470 68650 25726
rect 69310 25726 69314 25814
rect 69384 25726 69390 25942
rect 60110 25450 60200 25470
rect 60110 25380 60120 25450
rect 60190 25380 60200 25450
rect 60110 25370 60200 25380
rect 68560 25450 68650 25470
rect 68560 25380 68570 25450
rect 68640 25380 68650 25450
rect 68560 25370 68650 25380
rect 68890 25710 69070 25720
rect 68890 25650 68893 25710
rect 69067 25650 69070 25710
rect 68890 25250 69070 25650
rect 69310 25470 69390 25726
rect 69310 25450 69400 25470
rect 69310 25380 69320 25450
rect 69390 25380 69400 25450
rect 69310 25370 69400 25380
rect 79600 25250 81600 33130
rect 0 23250 81600 25250
rect 4176 16278 4246 16288
rect 4170 15846 4176 16240
rect 4914 16278 4984 16288
rect 4246 16234 4832 16240
rect 4246 16182 4554 16234
rect 4606 16182 4832 16234
rect 4246 16170 4832 16182
rect 4246 16118 4554 16170
rect 4606 16118 4832 16170
rect 4246 16112 4832 16118
rect 4246 15846 4250 16112
rect 4328 16056 4914 16062
rect 4328 16004 4468 16056
rect 4520 16004 4640 16056
rect 4692 16004 4914 16056
rect 4328 15992 4914 16004
rect 4328 15940 4468 15992
rect 4520 15940 4640 15992
rect 4692 15940 4914 15992
rect 4328 15934 4914 15940
rect 4170 15590 4250 15846
rect 4910 15846 4914 15934
rect 13376 16278 13446 16288
rect 4984 15846 4990 16062
rect 4160 15570 4250 15590
rect 4160 15500 4170 15570
rect 4240 15500 4250 15570
rect 4160 15490 4250 15500
rect 4490 15830 4670 15840
rect 4490 15770 4493 15830
rect 4667 15770 4670 15830
rect 4490 15370 4670 15770
rect 4910 15590 4990 15846
rect 13370 15846 13376 16240
rect 14114 16278 14184 16288
rect 13446 16234 14032 16240
rect 13446 16182 13754 16234
rect 13806 16182 14032 16234
rect 13446 16170 14032 16182
rect 13446 16118 13754 16170
rect 13806 16118 14032 16170
rect 13446 16112 14032 16118
rect 13446 15846 13450 16112
rect 13528 16056 14114 16062
rect 13528 16004 13668 16056
rect 13720 16004 13840 16056
rect 13892 16004 14114 16056
rect 13528 15992 14114 16004
rect 13528 15940 13668 15992
rect 13720 15940 13840 15992
rect 13892 15940 14114 15992
rect 13528 15934 14114 15940
rect 13370 15590 13450 15846
rect 14110 15846 14114 15934
rect 22576 16278 22646 16288
rect 14184 15846 14190 16062
rect 4910 15570 5000 15590
rect 4910 15500 4920 15570
rect 4990 15500 5000 15570
rect 4910 15490 5000 15500
rect 13360 15570 13450 15590
rect 13360 15500 13370 15570
rect 13440 15500 13450 15570
rect 13360 15490 13450 15500
rect 13690 15830 13870 15840
rect 13690 15770 13693 15830
rect 13867 15770 13870 15830
rect 13690 15370 13870 15770
rect 14110 15590 14190 15846
rect 22570 15846 22576 16240
rect 23314 16278 23384 16288
rect 22646 16234 23232 16240
rect 22646 16182 22954 16234
rect 23006 16182 23232 16234
rect 22646 16170 23232 16182
rect 22646 16118 22954 16170
rect 23006 16118 23232 16170
rect 22646 16112 23232 16118
rect 22646 15846 22650 16112
rect 22728 16056 23314 16062
rect 22728 16004 22868 16056
rect 22920 16004 23040 16056
rect 23092 16004 23314 16056
rect 22728 15992 23314 16004
rect 22728 15940 22868 15992
rect 22920 15940 23040 15992
rect 23092 15940 23314 15992
rect 22728 15934 23314 15940
rect 22570 15590 22650 15846
rect 23310 15846 23314 15934
rect 31776 16278 31846 16288
rect 23384 15846 23390 16062
rect 14110 15570 14200 15590
rect 14110 15500 14120 15570
rect 14190 15500 14200 15570
rect 14110 15490 14200 15500
rect 22560 15570 22650 15590
rect 22560 15500 22570 15570
rect 22640 15500 22650 15570
rect 22560 15490 22650 15500
rect 22890 15830 23070 15840
rect 22890 15770 22893 15830
rect 23067 15770 23070 15830
rect 22890 15370 23070 15770
rect 23310 15590 23390 15846
rect 31770 15846 31776 16240
rect 32514 16278 32584 16288
rect 31846 16234 32432 16240
rect 31846 16182 32154 16234
rect 32206 16182 32432 16234
rect 31846 16170 32432 16182
rect 31846 16118 32154 16170
rect 32206 16118 32432 16170
rect 31846 16112 32432 16118
rect 31846 15846 31850 16112
rect 31928 16056 32514 16062
rect 31928 16004 32068 16056
rect 32120 16004 32240 16056
rect 32292 16004 32514 16056
rect 31928 15992 32514 16004
rect 31928 15940 32068 15992
rect 32120 15940 32240 15992
rect 32292 15940 32514 15992
rect 31928 15934 32514 15940
rect 31770 15590 31850 15846
rect 32510 15846 32514 15934
rect 40976 16278 41046 16288
rect 32584 15846 32590 16062
rect 23310 15570 23400 15590
rect 23310 15500 23320 15570
rect 23390 15500 23400 15570
rect 23310 15490 23400 15500
rect 31760 15570 31850 15590
rect 31760 15500 31770 15570
rect 31840 15500 31850 15570
rect 31760 15490 31850 15500
rect 32090 15830 32270 15840
rect 32090 15770 32093 15830
rect 32267 15770 32270 15830
rect 32090 15370 32270 15770
rect 32510 15590 32590 15846
rect 40970 15846 40976 16240
rect 41714 16278 41784 16288
rect 41046 16234 41632 16240
rect 41046 16182 41354 16234
rect 41406 16182 41632 16234
rect 41046 16170 41632 16182
rect 41046 16118 41354 16170
rect 41406 16118 41632 16170
rect 41046 16112 41632 16118
rect 41046 15846 41050 16112
rect 41128 16056 41714 16062
rect 41128 16004 41268 16056
rect 41320 16004 41440 16056
rect 41492 16004 41714 16056
rect 41128 15992 41714 16004
rect 41128 15940 41268 15992
rect 41320 15940 41440 15992
rect 41492 15940 41714 15992
rect 41128 15934 41714 15940
rect 40970 15590 41050 15846
rect 41710 15846 41714 15934
rect 50176 16278 50246 16288
rect 41784 15846 41790 16062
rect 32510 15570 32600 15590
rect 32510 15500 32520 15570
rect 32590 15500 32600 15570
rect 32510 15490 32600 15500
rect 40960 15570 41050 15590
rect 40960 15500 40970 15570
rect 41040 15500 41050 15570
rect 40960 15490 41050 15500
rect 41290 15830 41470 15840
rect 41290 15770 41293 15830
rect 41467 15770 41470 15830
rect 41290 15370 41470 15770
rect 41710 15590 41790 15846
rect 50170 15846 50176 16240
rect 50914 16278 50984 16288
rect 50246 16234 50832 16240
rect 50246 16182 50554 16234
rect 50606 16182 50832 16234
rect 50246 16170 50832 16182
rect 50246 16118 50554 16170
rect 50606 16118 50832 16170
rect 50246 16112 50832 16118
rect 50246 15846 50250 16112
rect 50328 16056 50914 16062
rect 50328 16004 50468 16056
rect 50520 16004 50640 16056
rect 50692 16004 50914 16056
rect 50328 15992 50914 16004
rect 50328 15940 50468 15992
rect 50520 15940 50640 15992
rect 50692 15940 50914 15992
rect 50328 15934 50914 15940
rect 50170 15590 50250 15846
rect 50910 15846 50914 15934
rect 59376 16278 59446 16288
rect 50984 15846 50990 16062
rect 41710 15570 41800 15590
rect 41710 15500 41720 15570
rect 41790 15500 41800 15570
rect 41710 15490 41800 15500
rect 50160 15570 50250 15590
rect 50160 15500 50170 15570
rect 50240 15500 50250 15570
rect 50160 15490 50250 15500
rect 50490 15830 50670 15840
rect 50490 15770 50493 15830
rect 50667 15770 50670 15830
rect 50490 15370 50670 15770
rect 50910 15590 50990 15846
rect 59370 15846 59376 16240
rect 60114 16278 60184 16288
rect 59446 16234 60032 16240
rect 59446 16182 59754 16234
rect 59806 16182 60032 16234
rect 59446 16170 60032 16182
rect 59446 16118 59754 16170
rect 59806 16118 60032 16170
rect 59446 16112 60032 16118
rect 59446 15846 59450 16112
rect 59528 16056 60114 16062
rect 59528 16004 59668 16056
rect 59720 16004 59840 16056
rect 59892 16004 60114 16056
rect 59528 15992 60114 16004
rect 59528 15940 59668 15992
rect 59720 15940 59840 15992
rect 59892 15940 60114 15992
rect 59528 15934 60114 15940
rect 59370 15590 59450 15846
rect 60110 15846 60114 15934
rect 68576 16278 68646 16288
rect 60184 15846 60190 16062
rect 50910 15570 51000 15590
rect 50910 15500 50920 15570
rect 50990 15500 51000 15570
rect 50910 15490 51000 15500
rect 59360 15570 59450 15590
rect 59360 15500 59370 15570
rect 59440 15500 59450 15570
rect 59360 15490 59450 15500
rect 59690 15830 59870 15840
rect 59690 15770 59693 15830
rect 59867 15770 59870 15830
rect 59690 15370 59870 15770
rect 60110 15590 60190 15846
rect 68570 15846 68576 16240
rect 69314 16278 69384 16288
rect 68646 16234 69232 16240
rect 68646 16182 68954 16234
rect 69006 16182 69232 16234
rect 68646 16170 69232 16182
rect 68646 16118 68954 16170
rect 69006 16118 69232 16170
rect 68646 16112 69232 16118
rect 68646 15846 68650 16112
rect 68728 16056 69314 16062
rect 68728 16004 68868 16056
rect 68920 16004 69040 16056
rect 69092 16004 69314 16056
rect 68728 15992 69314 16004
rect 68728 15940 68868 15992
rect 68920 15940 69040 15992
rect 69092 15940 69314 15992
rect 68728 15934 69314 15940
rect 68570 15590 68650 15846
rect 69310 15846 69314 15934
rect 69384 15846 69390 16062
rect 60110 15570 60200 15590
rect 60110 15500 60120 15570
rect 60190 15500 60200 15570
rect 60110 15490 60200 15500
rect 68560 15570 68650 15590
rect 68560 15500 68570 15570
rect 68640 15500 68650 15570
rect 68560 15490 68650 15500
rect 68890 15830 69070 15840
rect 68890 15770 68893 15830
rect 69067 15770 69070 15830
rect 68890 15370 69070 15770
rect 69310 15590 69390 15846
rect 69310 15570 69400 15590
rect 69310 15500 69320 15570
rect 69390 15500 69400 15570
rect 69310 15490 69400 15500
rect 79600 15370 81600 23250
rect 0 13370 81600 15370
rect -6880 6620 -220 6640
rect -6880 6560 -490 6620
rect -240 6560 -220 6620
rect -6880 6540 -220 6560
rect -6880 -10 -4870 6540
rect 4176 6398 4246 6408
rect 4170 5966 4176 6360
rect 4914 6398 4984 6408
rect 4246 6354 4832 6360
rect 4246 6302 4554 6354
rect 4606 6302 4832 6354
rect 4246 6290 4832 6302
rect 4246 6238 4554 6290
rect 4606 6238 4832 6290
rect 4246 6232 4832 6238
rect 4246 5966 4250 6232
rect 4328 6176 4914 6182
rect 4328 6124 4468 6176
rect 4520 6124 4640 6176
rect 4692 6124 4914 6176
rect 4328 6112 4914 6124
rect 4328 6060 4468 6112
rect 4520 6060 4640 6112
rect 4692 6060 4914 6112
rect 4328 6054 4914 6060
rect -240 5830 0 5840
rect -240 5770 -230 5830
rect -170 5770 0 5830
rect -240 5760 0 5770
rect -160 5490 0 5760
rect 4170 5710 4250 5966
rect 4910 5966 4914 6054
rect 13376 6398 13446 6408
rect 4984 5966 4990 6182
rect 4160 5690 4250 5710
rect 4160 5620 4170 5690
rect 4240 5620 4250 5690
rect 4160 5610 4250 5620
rect 4490 5950 4670 5960
rect 4490 5890 4493 5950
rect 4667 5890 4670 5950
rect 4490 5490 4670 5890
rect 4910 5710 4990 5966
rect 13370 5966 13376 6360
rect 14114 6398 14184 6408
rect 13446 6354 14032 6360
rect 13446 6302 13754 6354
rect 13806 6302 14032 6354
rect 13446 6290 14032 6302
rect 13446 6238 13754 6290
rect 13806 6238 14032 6290
rect 13446 6232 14032 6238
rect 13446 5966 13450 6232
rect 13528 6176 14114 6182
rect 13528 6124 13668 6176
rect 13720 6124 13840 6176
rect 13892 6124 14114 6176
rect 13528 6112 14114 6124
rect 13528 6060 13668 6112
rect 13720 6060 13840 6112
rect 13892 6060 14114 6112
rect 13528 6054 14114 6060
rect 13370 5710 13450 5966
rect 14110 5966 14114 6054
rect 22576 6398 22646 6408
rect 14184 5966 14190 6182
rect 4910 5690 5000 5710
rect 4910 5620 4920 5690
rect 4990 5620 5000 5690
rect 4910 5610 5000 5620
rect 13360 5690 13450 5710
rect 13360 5620 13370 5690
rect 13440 5620 13450 5690
rect 13360 5610 13450 5620
rect 13690 5950 13870 5960
rect 13690 5890 13693 5950
rect 13867 5890 13870 5950
rect 13690 5490 13870 5890
rect 14110 5710 14190 5966
rect 22570 5966 22576 6360
rect 23314 6398 23384 6408
rect 22646 6354 23232 6360
rect 22646 6302 22954 6354
rect 23006 6302 23232 6354
rect 22646 6290 23232 6302
rect 22646 6238 22954 6290
rect 23006 6238 23232 6290
rect 22646 6232 23232 6238
rect 22646 5966 22650 6232
rect 22728 6176 23314 6182
rect 22728 6124 22868 6176
rect 22920 6124 23040 6176
rect 23092 6124 23314 6176
rect 22728 6112 23314 6124
rect 22728 6060 22868 6112
rect 22920 6060 23040 6112
rect 23092 6060 23314 6112
rect 22728 6054 23314 6060
rect 22570 5710 22650 5966
rect 23310 5966 23314 6054
rect 31776 6398 31846 6408
rect 23384 5966 23390 6182
rect 14110 5690 14200 5710
rect 14110 5620 14120 5690
rect 14190 5620 14200 5690
rect 14110 5610 14200 5620
rect 22560 5690 22650 5710
rect 22560 5620 22570 5690
rect 22640 5620 22650 5690
rect 22560 5610 22650 5620
rect 22890 5950 23070 5960
rect 22890 5890 22893 5950
rect 23067 5890 23070 5950
rect 22890 5490 23070 5890
rect 23310 5710 23390 5966
rect 31770 5966 31776 6360
rect 32514 6398 32584 6408
rect 31846 6354 32432 6360
rect 31846 6302 32154 6354
rect 32206 6302 32432 6354
rect 31846 6290 32432 6302
rect 31846 6238 32154 6290
rect 32206 6238 32432 6290
rect 31846 6232 32432 6238
rect 31846 5966 31850 6232
rect 31928 6176 32514 6182
rect 31928 6124 32068 6176
rect 32120 6124 32240 6176
rect 32292 6124 32514 6176
rect 31928 6112 32514 6124
rect 31928 6060 32068 6112
rect 32120 6060 32240 6112
rect 32292 6060 32514 6112
rect 31928 6054 32514 6060
rect 31770 5710 31850 5966
rect 32510 5966 32514 6054
rect 40976 6398 41046 6408
rect 32584 5966 32590 6182
rect 23310 5690 23400 5710
rect 23310 5620 23320 5690
rect 23390 5620 23400 5690
rect 23310 5610 23400 5620
rect 31760 5690 31850 5710
rect 31760 5620 31770 5690
rect 31840 5620 31850 5690
rect 31760 5610 31850 5620
rect 32090 5950 32270 5960
rect 32090 5890 32093 5950
rect 32267 5890 32270 5950
rect 32090 5490 32270 5890
rect 32510 5710 32590 5966
rect 40970 5966 40976 6360
rect 41714 6398 41784 6408
rect 41046 6354 41632 6360
rect 41046 6302 41354 6354
rect 41406 6302 41632 6354
rect 41046 6290 41632 6302
rect 41046 6238 41354 6290
rect 41406 6238 41632 6290
rect 41046 6232 41632 6238
rect 41046 5966 41050 6232
rect 41128 6176 41714 6182
rect 41128 6124 41268 6176
rect 41320 6124 41440 6176
rect 41492 6124 41714 6176
rect 41128 6112 41714 6124
rect 41128 6060 41268 6112
rect 41320 6060 41440 6112
rect 41492 6060 41714 6112
rect 41128 6054 41714 6060
rect 40970 5710 41050 5966
rect 41710 5966 41714 6054
rect 50176 6398 50246 6408
rect 41784 5966 41790 6182
rect 32510 5690 32600 5710
rect 32510 5620 32520 5690
rect 32590 5620 32600 5690
rect 32510 5610 32600 5620
rect 40960 5690 41050 5710
rect 40960 5620 40970 5690
rect 41040 5620 41050 5690
rect 40960 5610 41050 5620
rect 41290 5950 41470 5960
rect 41290 5890 41293 5950
rect 41467 5890 41470 5950
rect 41290 5490 41470 5890
rect 41710 5710 41790 5966
rect 50170 5966 50176 6360
rect 50914 6398 50984 6408
rect 50246 6354 50832 6360
rect 50246 6302 50554 6354
rect 50606 6302 50832 6354
rect 50246 6290 50832 6302
rect 50246 6238 50554 6290
rect 50606 6238 50832 6290
rect 50246 6232 50832 6238
rect 50246 5966 50250 6232
rect 50328 6176 50914 6182
rect 50328 6124 50468 6176
rect 50520 6124 50640 6176
rect 50692 6124 50914 6176
rect 50328 6112 50914 6124
rect 50328 6060 50468 6112
rect 50520 6060 50640 6112
rect 50692 6060 50914 6112
rect 50328 6054 50914 6060
rect 50170 5710 50250 5966
rect 50910 5966 50914 6054
rect 59376 6398 59446 6408
rect 50984 5966 50990 6182
rect 41710 5690 41800 5710
rect 41710 5620 41720 5690
rect 41790 5620 41800 5690
rect 41710 5610 41800 5620
rect 50160 5690 50250 5710
rect 50160 5620 50170 5690
rect 50240 5620 50250 5690
rect 50160 5610 50250 5620
rect 50490 5950 50670 5960
rect 50490 5890 50493 5950
rect 50667 5890 50670 5950
rect 50490 5490 50670 5890
rect 50910 5710 50990 5966
rect 59370 5966 59376 6360
rect 60114 6398 60184 6408
rect 59446 6354 60032 6360
rect 59446 6302 59754 6354
rect 59806 6302 60032 6354
rect 59446 6290 60032 6302
rect 59446 6238 59754 6290
rect 59806 6238 60032 6290
rect 59446 6232 60032 6238
rect 59446 5966 59450 6232
rect 59528 6176 60114 6182
rect 59528 6124 59668 6176
rect 59720 6124 59840 6176
rect 59892 6124 60114 6176
rect 59528 6112 60114 6124
rect 59528 6060 59668 6112
rect 59720 6060 59840 6112
rect 59892 6060 60114 6112
rect 59528 6054 60114 6060
rect 59370 5710 59450 5966
rect 60110 5966 60114 6054
rect 68576 6398 68646 6408
rect 60184 5966 60190 6182
rect 50910 5690 51000 5710
rect 50910 5620 50920 5690
rect 50990 5620 51000 5690
rect 50910 5610 51000 5620
rect 59360 5690 59450 5710
rect 59360 5620 59370 5690
rect 59440 5620 59450 5690
rect 59360 5610 59450 5620
rect 59690 5950 59870 5960
rect 59690 5890 59693 5950
rect 59867 5890 59870 5950
rect 59690 5490 59870 5890
rect 60110 5710 60190 5966
rect 68570 5966 68576 6360
rect 69314 6398 69384 6408
rect 68646 6354 69232 6360
rect 68646 6302 68954 6354
rect 69006 6302 69232 6354
rect 68646 6290 69232 6302
rect 68646 6238 68954 6290
rect 69006 6238 69232 6290
rect 68646 6232 69232 6238
rect 68646 5966 68650 6232
rect 68728 6176 69314 6182
rect 68728 6124 68868 6176
rect 68920 6124 69040 6176
rect 69092 6124 69314 6176
rect 68728 6112 69314 6124
rect 68728 6060 68868 6112
rect 68920 6060 69040 6112
rect 69092 6060 69314 6112
rect 68728 6054 69314 6060
rect 68570 5710 68650 5966
rect 69310 5966 69314 6054
rect 69384 5966 69390 6182
rect 60110 5690 60200 5710
rect 60110 5620 60120 5690
rect 60190 5620 60200 5690
rect 60110 5610 60200 5620
rect 68560 5690 68650 5710
rect 68560 5620 68570 5690
rect 68640 5620 68650 5690
rect 68560 5610 68650 5620
rect 68890 5950 69070 5960
rect 68890 5890 68893 5950
rect 69067 5890 69070 5950
rect 68890 5490 69070 5890
rect 69310 5710 69390 5966
rect 69310 5690 69400 5710
rect 69310 5620 69320 5690
rect 69390 5620 69400 5690
rect 69310 5610 69400 5620
rect 79600 5490 81600 13370
rect -160 3490 82600 5490
<< via2 >>
rect 4170 94540 4240 94610
rect 4920 94540 4990 94610
rect 4170 84660 4240 84730
rect 4920 84660 4990 84730
rect 13370 84660 13440 84730
rect 14120 84660 14190 84730
rect 4170 74780 4240 74850
rect 4920 74780 4990 74850
rect 13370 74780 13440 74850
rect 14120 74780 14190 74850
rect 22570 74780 22640 74850
rect 23320 74780 23390 74850
rect 31770 74780 31840 74850
rect 32520 74780 32590 74850
rect 4170 64900 4240 64970
rect 4920 64900 4990 64970
rect 13370 64900 13440 64970
rect 14120 64900 14190 64970
rect 22570 64900 22640 64970
rect 23320 64900 23390 64970
rect 31770 64900 31840 64970
rect 32520 64900 32590 64970
rect 40970 64900 41040 64970
rect 41720 64900 41790 64970
rect 50170 64900 50240 64970
rect 50920 64900 50990 64970
rect 59370 64900 59440 64970
rect 60120 64900 60190 64970
rect 68570 64900 68640 64970
rect 69320 64900 69390 64970
rect 4170 55020 4240 55090
rect 4920 55020 4990 55090
rect 13370 55020 13440 55090
rect 14120 55020 14190 55090
rect 22570 55020 22640 55090
rect 23320 55020 23390 55090
rect 31770 55020 31840 55090
rect 32520 55020 32590 55090
rect 40970 55020 41040 55090
rect 41720 55020 41790 55090
rect 50170 55020 50240 55090
rect 50920 55020 50990 55090
rect 59370 55020 59440 55090
rect 60120 55020 60190 55090
rect 68570 55020 68640 55090
rect 69320 55020 69390 55090
rect 4170 45140 4240 45210
rect 4920 45140 4990 45210
rect 13370 45140 13440 45210
rect 14120 45140 14190 45210
rect 22570 45140 22640 45210
rect 23320 45140 23390 45210
rect 31770 45140 31840 45210
rect 32520 45140 32590 45210
rect 40970 45140 41040 45210
rect 41720 45140 41790 45210
rect 50170 45140 50240 45210
rect 50920 45140 50990 45210
rect 59370 45140 59440 45210
rect 60120 45140 60190 45210
rect 68570 45140 68640 45210
rect 69320 45140 69390 45210
rect 4170 35260 4240 35330
rect 4920 35260 4990 35330
rect 13370 35260 13440 35330
rect 14120 35260 14190 35330
rect 22570 35260 22640 35330
rect 23320 35260 23390 35330
rect 31770 35260 31840 35330
rect 32520 35260 32590 35330
rect 40970 35260 41040 35330
rect 41720 35260 41790 35330
rect 50170 35260 50240 35330
rect 50920 35260 50990 35330
rect 59370 35260 59440 35330
rect 60120 35260 60190 35330
rect 68570 35260 68640 35330
rect 69320 35260 69390 35330
rect 4170 25380 4240 25450
rect 4920 25380 4990 25450
rect 13370 25380 13440 25450
rect 14120 25380 14190 25450
rect 22570 25380 22640 25450
rect 23320 25380 23390 25450
rect 31770 25380 31840 25450
rect 32520 25380 32590 25450
rect 40970 25380 41040 25450
rect 41720 25380 41790 25450
rect 50170 25380 50240 25450
rect 50920 25380 50990 25450
rect 59370 25380 59440 25450
rect 60120 25380 60190 25450
rect 68570 25380 68640 25450
rect 69320 25380 69390 25450
rect 4170 15500 4240 15570
rect 4920 15500 4990 15570
rect 13370 15500 13440 15570
rect 14120 15500 14190 15570
rect 22570 15500 22640 15570
rect 23320 15500 23390 15570
rect 31770 15500 31840 15570
rect 32520 15500 32590 15570
rect 40970 15500 41040 15570
rect 41720 15500 41790 15570
rect 50170 15500 50240 15570
rect 50920 15500 50990 15570
rect 59370 15500 59440 15570
rect 60120 15500 60190 15570
rect 68570 15500 68640 15570
rect 69320 15500 69390 15570
rect 4170 5620 4240 5690
rect 4920 5620 4990 5690
rect 13370 5620 13440 5690
rect 14120 5620 14190 5690
rect 22570 5620 22640 5690
rect 23320 5620 23390 5690
rect 31770 5620 31840 5690
rect 32520 5620 32590 5690
rect 40970 5620 41040 5690
rect 41720 5620 41790 5690
rect 50170 5620 50240 5690
rect 50920 5620 50990 5690
rect 59370 5620 59440 5690
rect 60120 5620 60190 5690
rect 68570 5620 68640 5690
rect 69320 5620 69390 5690
<< metal3 >>
rect -6874 109790 70726 109796
rect -9760 107810 6220 109790
rect 8200 107810 15420 109790
rect 17400 107810 24620 109790
rect 26600 107810 33820 109790
rect 35800 107810 43020 109790
rect 45000 107810 52220 109790
rect 54200 109780 70726 109790
rect 72610 109780 82600 109800
rect 54200 107810 61420 109780
rect -9760 107800 61420 107810
rect 63400 107800 70620 109780
rect 72600 107800 82600 109780
rect -9760 107790 72610 107800
rect -9760 103780 70720 103790
rect 72610 103780 82600 103790
rect -9760 101800 1010 103780
rect 2990 101800 10210 103780
rect 12190 101800 19410 103780
rect 21390 101800 28610 103780
rect 30590 101800 37810 103780
rect 39790 101800 47010 103780
rect 48990 101800 56210 103780
rect 58190 101800 65410 103780
rect 67390 101800 82600 103780
rect -9760 101790 82600 101800
rect 3085 95702 4044 95730
rect 3085 94898 3960 95702
rect 4024 94898 4044 95702
rect 3085 94870 4044 94898
rect 5164 95702 6123 95730
rect 5164 94898 5184 95702
rect 5248 94898 6123 95702
rect 5164 94870 6123 94898
rect 3940 94620 4260 94630
rect 3940 94530 3950 94620
rect 4030 94610 4260 94620
rect 4030 94540 4170 94610
rect 4240 94540 4260 94610
rect 4030 94530 4260 94540
rect 3940 94520 4260 94530
rect 4900 94620 5270 94630
rect 4900 94610 5180 94620
rect 4900 94540 4920 94610
rect 4990 94540 5180 94610
rect 4900 94530 5180 94540
rect 5260 94530 5270 94620
rect 4900 94520 5270 94530
rect 3085 85822 4044 85850
rect 3085 85018 3960 85822
rect 4024 85018 4044 85822
rect 3085 84990 4044 85018
rect 5164 85822 6123 85850
rect 5164 85018 5184 85822
rect 5248 85018 6123 85822
rect 5164 84990 6123 85018
rect 12285 85822 13244 85850
rect 12285 85018 13160 85822
rect 13224 85018 13244 85822
rect 12285 84990 13244 85018
rect 14364 85822 15323 85850
rect 14364 85018 14384 85822
rect 14448 85018 15323 85822
rect 14364 84990 15323 85018
rect 3940 84740 4260 84750
rect 3940 84650 3950 84740
rect 4030 84730 4260 84740
rect 4030 84660 4170 84730
rect 4240 84660 4260 84730
rect 4030 84650 4260 84660
rect 3940 84640 4260 84650
rect 4900 84740 5270 84750
rect 4900 84730 5180 84740
rect 4900 84660 4920 84730
rect 4990 84660 5180 84730
rect 4900 84650 5180 84660
rect 5260 84650 5270 84740
rect 4900 84640 5270 84650
rect 13140 84740 13460 84750
rect 13140 84650 13150 84740
rect 13230 84730 13460 84740
rect 13230 84660 13370 84730
rect 13440 84660 13460 84730
rect 13230 84650 13460 84660
rect 13140 84640 13460 84650
rect 14100 84740 14470 84750
rect 14100 84730 14380 84740
rect 14100 84660 14120 84730
rect 14190 84660 14380 84730
rect 14100 84650 14380 84660
rect 14460 84650 14470 84740
rect 14100 84640 14470 84650
rect 3085 75942 4044 75970
rect 3085 75138 3960 75942
rect 4024 75138 4044 75942
rect 3085 75110 4044 75138
rect 5164 75942 6123 75970
rect 5164 75138 5184 75942
rect 5248 75138 6123 75942
rect 5164 75110 6123 75138
rect 12285 75942 13244 75970
rect 12285 75138 13160 75942
rect 13224 75138 13244 75942
rect 12285 75110 13244 75138
rect 14364 75942 15323 75970
rect 14364 75138 14384 75942
rect 14448 75138 15323 75942
rect 14364 75110 15323 75138
rect 21485 75942 22444 75970
rect 21485 75138 22360 75942
rect 22424 75138 22444 75942
rect 21485 75110 22444 75138
rect 23564 75942 24523 75970
rect 23564 75138 23584 75942
rect 23648 75138 24523 75942
rect 23564 75110 24523 75138
rect 30685 75942 31644 75970
rect 30685 75138 31560 75942
rect 31624 75138 31644 75942
rect 30685 75110 31644 75138
rect 32764 75942 33723 75970
rect 32764 75138 32784 75942
rect 32848 75138 33723 75942
rect 32764 75110 33723 75138
rect 3940 74860 4260 74870
rect 3940 74770 3950 74860
rect 4030 74850 4260 74860
rect 4030 74780 4170 74850
rect 4240 74780 4260 74850
rect 4030 74770 4260 74780
rect 3940 74760 4260 74770
rect 4900 74860 5270 74870
rect 4900 74850 5180 74860
rect 4900 74780 4920 74850
rect 4990 74780 5180 74850
rect 4900 74770 5180 74780
rect 5260 74770 5270 74860
rect 4900 74760 5270 74770
rect 13140 74860 13460 74870
rect 13140 74770 13150 74860
rect 13230 74850 13460 74860
rect 13230 74780 13370 74850
rect 13440 74780 13460 74850
rect 13230 74770 13460 74780
rect 13140 74760 13460 74770
rect 14100 74860 14470 74870
rect 14100 74850 14380 74860
rect 14100 74780 14120 74850
rect 14190 74780 14380 74850
rect 14100 74770 14380 74780
rect 14460 74770 14470 74860
rect 14100 74760 14470 74770
rect 22340 74860 22660 74870
rect 22340 74770 22350 74860
rect 22430 74850 22660 74860
rect 22430 74780 22570 74850
rect 22640 74780 22660 74850
rect 22430 74770 22660 74780
rect 22340 74760 22660 74770
rect 23300 74860 23670 74870
rect 23300 74850 23580 74860
rect 23300 74780 23320 74850
rect 23390 74780 23580 74850
rect 23300 74770 23580 74780
rect 23660 74770 23670 74860
rect 23300 74760 23670 74770
rect 31540 74860 31860 74870
rect 31540 74770 31550 74860
rect 31630 74850 31860 74860
rect 31630 74780 31770 74850
rect 31840 74780 31860 74850
rect 31630 74770 31860 74780
rect 31540 74760 31860 74770
rect 32500 74860 32870 74870
rect 32500 74850 32780 74860
rect 32500 74780 32520 74850
rect 32590 74780 32780 74850
rect 32500 74770 32780 74780
rect 32860 74770 32870 74860
rect 32500 74760 32870 74770
rect 3085 66062 4044 66090
rect 3085 65258 3960 66062
rect 4024 65258 4044 66062
rect 3085 65230 4044 65258
rect 5164 66062 6123 66090
rect 5164 65258 5184 66062
rect 5248 65258 6123 66062
rect 5164 65230 6123 65258
rect 12285 66062 13244 66090
rect 12285 65258 13160 66062
rect 13224 65258 13244 66062
rect 12285 65230 13244 65258
rect 14364 66062 15323 66090
rect 14364 65258 14384 66062
rect 14448 65258 15323 66062
rect 14364 65230 15323 65258
rect 21485 66062 22444 66090
rect 21485 65258 22360 66062
rect 22424 65258 22444 66062
rect 21485 65230 22444 65258
rect 23564 66062 24523 66090
rect 23564 65258 23584 66062
rect 23648 65258 24523 66062
rect 23564 65230 24523 65258
rect 30685 66062 31644 66090
rect 30685 65258 31560 66062
rect 31624 65258 31644 66062
rect 30685 65230 31644 65258
rect 32764 66062 33723 66090
rect 32764 65258 32784 66062
rect 32848 65258 33723 66062
rect 32764 65230 33723 65258
rect 39885 66062 40844 66090
rect 39885 65258 40760 66062
rect 40824 65258 40844 66062
rect 39885 65230 40844 65258
rect 41964 66062 42923 66090
rect 41964 65258 41984 66062
rect 42048 65258 42923 66062
rect 41964 65230 42923 65258
rect 49085 66062 50044 66090
rect 49085 65258 49960 66062
rect 50024 65258 50044 66062
rect 49085 65230 50044 65258
rect 51164 66062 52123 66090
rect 51164 65258 51184 66062
rect 51248 65258 52123 66062
rect 51164 65230 52123 65258
rect 58285 66062 59244 66090
rect 58285 65258 59160 66062
rect 59224 65258 59244 66062
rect 58285 65230 59244 65258
rect 60364 66062 61323 66090
rect 60364 65258 60384 66062
rect 60448 65258 61323 66062
rect 60364 65230 61323 65258
rect 67485 66062 68444 66090
rect 67485 65258 68360 66062
rect 68424 65258 68444 66062
rect 67485 65230 68444 65258
rect 69564 66062 70523 66090
rect 69564 65258 69584 66062
rect 69648 65258 70523 66062
rect 69564 65230 70523 65258
rect 3940 64980 4260 64990
rect 3940 64890 3950 64980
rect 4030 64970 4260 64980
rect 4030 64900 4170 64970
rect 4240 64900 4260 64970
rect 4030 64890 4260 64900
rect 3940 64880 4260 64890
rect 4900 64980 5270 64990
rect 4900 64970 5180 64980
rect 4900 64900 4920 64970
rect 4990 64900 5180 64970
rect 4900 64890 5180 64900
rect 5260 64890 5270 64980
rect 4900 64880 5270 64890
rect 13140 64980 13460 64990
rect 13140 64890 13150 64980
rect 13230 64970 13460 64980
rect 13230 64900 13370 64970
rect 13440 64900 13460 64970
rect 13230 64890 13460 64900
rect 13140 64880 13460 64890
rect 14100 64980 14470 64990
rect 14100 64970 14380 64980
rect 14100 64900 14120 64970
rect 14190 64900 14380 64970
rect 14100 64890 14380 64900
rect 14460 64890 14470 64980
rect 14100 64880 14470 64890
rect 22340 64980 22660 64990
rect 22340 64890 22350 64980
rect 22430 64970 22660 64980
rect 22430 64900 22570 64970
rect 22640 64900 22660 64970
rect 22430 64890 22660 64900
rect 22340 64880 22660 64890
rect 23300 64980 23670 64990
rect 23300 64970 23580 64980
rect 23300 64900 23320 64970
rect 23390 64900 23580 64970
rect 23300 64890 23580 64900
rect 23660 64890 23670 64980
rect 23300 64880 23670 64890
rect 31540 64980 31860 64990
rect 31540 64890 31550 64980
rect 31630 64970 31860 64980
rect 31630 64900 31770 64970
rect 31840 64900 31860 64970
rect 31630 64890 31860 64900
rect 31540 64880 31860 64890
rect 32500 64980 32870 64990
rect 32500 64970 32780 64980
rect 32500 64900 32520 64970
rect 32590 64900 32780 64970
rect 32500 64890 32780 64900
rect 32860 64890 32870 64980
rect 32500 64880 32870 64890
rect 40740 64980 41060 64990
rect 40740 64890 40750 64980
rect 40830 64970 41060 64980
rect 40830 64900 40970 64970
rect 41040 64900 41060 64970
rect 40830 64890 41060 64900
rect 40740 64880 41060 64890
rect 41700 64980 42070 64990
rect 41700 64970 41980 64980
rect 41700 64900 41720 64970
rect 41790 64900 41980 64970
rect 41700 64890 41980 64900
rect 42060 64890 42070 64980
rect 41700 64880 42070 64890
rect 49940 64980 50260 64990
rect 49940 64890 49950 64980
rect 50030 64970 50260 64980
rect 50030 64900 50170 64970
rect 50240 64900 50260 64970
rect 50030 64890 50260 64900
rect 49940 64880 50260 64890
rect 50900 64980 51270 64990
rect 50900 64970 51180 64980
rect 50900 64900 50920 64970
rect 50990 64900 51180 64970
rect 50900 64890 51180 64900
rect 51260 64890 51270 64980
rect 50900 64880 51270 64890
rect 59140 64980 59460 64990
rect 59140 64890 59150 64980
rect 59230 64970 59460 64980
rect 59230 64900 59370 64970
rect 59440 64900 59460 64970
rect 59230 64890 59460 64900
rect 59140 64880 59460 64890
rect 60100 64980 60470 64990
rect 60100 64970 60380 64980
rect 60100 64900 60120 64970
rect 60190 64900 60380 64970
rect 60100 64890 60380 64900
rect 60460 64890 60470 64980
rect 60100 64880 60470 64890
rect 68340 64980 68660 64990
rect 68340 64890 68350 64980
rect 68430 64970 68660 64980
rect 68430 64900 68570 64970
rect 68640 64900 68660 64970
rect 68430 64890 68660 64900
rect 68340 64880 68660 64890
rect 69300 64980 69670 64990
rect 69300 64970 69580 64980
rect 69300 64900 69320 64970
rect 69390 64900 69580 64970
rect 69300 64890 69580 64900
rect 69660 64890 69670 64980
rect 69300 64880 69670 64890
rect 3085 56182 4044 56210
rect 3085 55378 3960 56182
rect 4024 55378 4044 56182
rect 3085 55350 4044 55378
rect 5164 56182 6123 56210
rect 5164 55378 5184 56182
rect 5248 55378 6123 56182
rect 5164 55350 6123 55378
rect 12285 56182 13244 56210
rect 12285 55378 13160 56182
rect 13224 55378 13244 56182
rect 12285 55350 13244 55378
rect 14364 56182 15323 56210
rect 14364 55378 14384 56182
rect 14448 55378 15323 56182
rect 14364 55350 15323 55378
rect 21485 56182 22444 56210
rect 21485 55378 22360 56182
rect 22424 55378 22444 56182
rect 21485 55350 22444 55378
rect 23564 56182 24523 56210
rect 23564 55378 23584 56182
rect 23648 55378 24523 56182
rect 23564 55350 24523 55378
rect 30685 56182 31644 56210
rect 30685 55378 31560 56182
rect 31624 55378 31644 56182
rect 30685 55350 31644 55378
rect 32764 56182 33723 56210
rect 32764 55378 32784 56182
rect 32848 55378 33723 56182
rect 32764 55350 33723 55378
rect 39885 56182 40844 56210
rect 39885 55378 40760 56182
rect 40824 55378 40844 56182
rect 39885 55350 40844 55378
rect 41964 56182 42923 56210
rect 41964 55378 41984 56182
rect 42048 55378 42923 56182
rect 41964 55350 42923 55378
rect 49085 56182 50044 56210
rect 49085 55378 49960 56182
rect 50024 55378 50044 56182
rect 49085 55350 50044 55378
rect 51164 56182 52123 56210
rect 51164 55378 51184 56182
rect 51248 55378 52123 56182
rect 51164 55350 52123 55378
rect 58285 56182 59244 56210
rect 58285 55378 59160 56182
rect 59224 55378 59244 56182
rect 58285 55350 59244 55378
rect 60364 56182 61323 56210
rect 60364 55378 60384 56182
rect 60448 55378 61323 56182
rect 60364 55350 61323 55378
rect 67485 56182 68444 56210
rect 67485 55378 68360 56182
rect 68424 55378 68444 56182
rect 67485 55350 68444 55378
rect 69564 56182 70523 56210
rect 69564 55378 69584 56182
rect 69648 55378 70523 56182
rect 69564 55350 70523 55378
rect 3940 55100 4260 55110
rect 3940 55010 3950 55100
rect 4030 55090 4260 55100
rect 4030 55020 4170 55090
rect 4240 55020 4260 55090
rect 4030 55010 4260 55020
rect 3940 55000 4260 55010
rect 4900 55100 5270 55110
rect 4900 55090 5180 55100
rect 4900 55020 4920 55090
rect 4990 55020 5180 55090
rect 4900 55010 5180 55020
rect 5260 55010 5270 55100
rect 4900 55000 5270 55010
rect 13140 55100 13460 55110
rect 13140 55010 13150 55100
rect 13230 55090 13460 55100
rect 13230 55020 13370 55090
rect 13440 55020 13460 55090
rect 13230 55010 13460 55020
rect 13140 55000 13460 55010
rect 14100 55100 14470 55110
rect 14100 55090 14380 55100
rect 14100 55020 14120 55090
rect 14190 55020 14380 55090
rect 14100 55010 14380 55020
rect 14460 55010 14470 55100
rect 14100 55000 14470 55010
rect 22340 55100 22660 55110
rect 22340 55010 22350 55100
rect 22430 55090 22660 55100
rect 22430 55020 22570 55090
rect 22640 55020 22660 55090
rect 22430 55010 22660 55020
rect 22340 55000 22660 55010
rect 23300 55100 23670 55110
rect 23300 55090 23580 55100
rect 23300 55020 23320 55090
rect 23390 55020 23580 55090
rect 23300 55010 23580 55020
rect 23660 55010 23670 55100
rect 23300 55000 23670 55010
rect 31540 55100 31860 55110
rect 31540 55010 31550 55100
rect 31630 55090 31860 55100
rect 31630 55020 31770 55090
rect 31840 55020 31860 55090
rect 31630 55010 31860 55020
rect 31540 55000 31860 55010
rect 32500 55100 32870 55110
rect 32500 55090 32780 55100
rect 32500 55020 32520 55090
rect 32590 55020 32780 55090
rect 32500 55010 32780 55020
rect 32860 55010 32870 55100
rect 32500 55000 32870 55010
rect 40740 55100 41060 55110
rect 40740 55010 40750 55100
rect 40830 55090 41060 55100
rect 40830 55020 40970 55090
rect 41040 55020 41060 55090
rect 40830 55010 41060 55020
rect 40740 55000 41060 55010
rect 41700 55100 42070 55110
rect 41700 55090 41980 55100
rect 41700 55020 41720 55090
rect 41790 55020 41980 55090
rect 41700 55010 41980 55020
rect 42060 55010 42070 55100
rect 41700 55000 42070 55010
rect 49940 55100 50260 55110
rect 49940 55010 49950 55100
rect 50030 55090 50260 55100
rect 50030 55020 50170 55090
rect 50240 55020 50260 55090
rect 50030 55010 50260 55020
rect 49940 55000 50260 55010
rect 50900 55100 51270 55110
rect 50900 55090 51180 55100
rect 50900 55020 50920 55090
rect 50990 55020 51180 55090
rect 50900 55010 51180 55020
rect 51260 55010 51270 55100
rect 50900 55000 51270 55010
rect 59140 55100 59460 55110
rect 59140 55010 59150 55100
rect 59230 55090 59460 55100
rect 59230 55020 59370 55090
rect 59440 55020 59460 55090
rect 59230 55010 59460 55020
rect 59140 55000 59460 55010
rect 60100 55100 60470 55110
rect 60100 55090 60380 55100
rect 60100 55020 60120 55090
rect 60190 55020 60380 55090
rect 60100 55010 60380 55020
rect 60460 55010 60470 55100
rect 60100 55000 60470 55010
rect 68340 55100 68660 55110
rect 68340 55010 68350 55100
rect 68430 55090 68660 55100
rect 68430 55020 68570 55090
rect 68640 55020 68660 55090
rect 68430 55010 68660 55020
rect 68340 55000 68660 55010
rect 69300 55100 69670 55110
rect 69300 55090 69580 55100
rect 69300 55020 69320 55090
rect 69390 55020 69580 55090
rect 69300 55010 69580 55020
rect 69660 55010 69670 55100
rect 69300 55000 69670 55010
rect 3085 46302 4044 46330
rect 3085 45498 3960 46302
rect 4024 45498 4044 46302
rect 3085 45470 4044 45498
rect 5164 46302 6123 46330
rect 5164 45498 5184 46302
rect 5248 45498 6123 46302
rect 5164 45470 6123 45498
rect 12285 46302 13244 46330
rect 12285 45498 13160 46302
rect 13224 45498 13244 46302
rect 12285 45470 13244 45498
rect 14364 46302 15323 46330
rect 14364 45498 14384 46302
rect 14448 45498 15323 46302
rect 14364 45470 15323 45498
rect 21485 46302 22444 46330
rect 21485 45498 22360 46302
rect 22424 45498 22444 46302
rect 21485 45470 22444 45498
rect 23564 46302 24523 46330
rect 23564 45498 23584 46302
rect 23648 45498 24523 46302
rect 23564 45470 24523 45498
rect 30685 46302 31644 46330
rect 30685 45498 31560 46302
rect 31624 45498 31644 46302
rect 30685 45470 31644 45498
rect 32764 46302 33723 46330
rect 32764 45498 32784 46302
rect 32848 45498 33723 46302
rect 32764 45470 33723 45498
rect 39885 46302 40844 46330
rect 39885 45498 40760 46302
rect 40824 45498 40844 46302
rect 39885 45470 40844 45498
rect 41964 46302 42923 46330
rect 41964 45498 41984 46302
rect 42048 45498 42923 46302
rect 41964 45470 42923 45498
rect 49085 46302 50044 46330
rect 49085 45498 49960 46302
rect 50024 45498 50044 46302
rect 49085 45470 50044 45498
rect 51164 46302 52123 46330
rect 51164 45498 51184 46302
rect 51248 45498 52123 46302
rect 51164 45470 52123 45498
rect 58285 46302 59244 46330
rect 58285 45498 59160 46302
rect 59224 45498 59244 46302
rect 58285 45470 59244 45498
rect 60364 46302 61323 46330
rect 60364 45498 60384 46302
rect 60448 45498 61323 46302
rect 60364 45470 61323 45498
rect 67485 46302 68444 46330
rect 67485 45498 68360 46302
rect 68424 45498 68444 46302
rect 67485 45470 68444 45498
rect 69564 46302 70523 46330
rect 69564 45498 69584 46302
rect 69648 45498 70523 46302
rect 69564 45470 70523 45498
rect 3940 45220 4260 45230
rect 3940 45130 3950 45220
rect 4030 45210 4260 45220
rect 4030 45140 4170 45210
rect 4240 45140 4260 45210
rect 4030 45130 4260 45140
rect 3940 45120 4260 45130
rect 4900 45220 5270 45230
rect 4900 45210 5180 45220
rect 4900 45140 4920 45210
rect 4990 45140 5180 45210
rect 4900 45130 5180 45140
rect 5260 45130 5270 45220
rect 4900 45120 5270 45130
rect 13140 45220 13460 45230
rect 13140 45130 13150 45220
rect 13230 45210 13460 45220
rect 13230 45140 13370 45210
rect 13440 45140 13460 45210
rect 13230 45130 13460 45140
rect 13140 45120 13460 45130
rect 14100 45220 14470 45230
rect 14100 45210 14380 45220
rect 14100 45140 14120 45210
rect 14190 45140 14380 45210
rect 14100 45130 14380 45140
rect 14460 45130 14470 45220
rect 14100 45120 14470 45130
rect 22340 45220 22660 45230
rect 22340 45130 22350 45220
rect 22430 45210 22660 45220
rect 22430 45140 22570 45210
rect 22640 45140 22660 45210
rect 22430 45130 22660 45140
rect 22340 45120 22660 45130
rect 23300 45220 23670 45230
rect 23300 45210 23580 45220
rect 23300 45140 23320 45210
rect 23390 45140 23580 45210
rect 23300 45130 23580 45140
rect 23660 45130 23670 45220
rect 23300 45120 23670 45130
rect 31540 45220 31860 45230
rect 31540 45130 31550 45220
rect 31630 45210 31860 45220
rect 31630 45140 31770 45210
rect 31840 45140 31860 45210
rect 31630 45130 31860 45140
rect 31540 45120 31860 45130
rect 32500 45220 32870 45230
rect 32500 45210 32780 45220
rect 32500 45140 32520 45210
rect 32590 45140 32780 45210
rect 32500 45130 32780 45140
rect 32860 45130 32870 45220
rect 32500 45120 32870 45130
rect 40740 45220 41060 45230
rect 40740 45130 40750 45220
rect 40830 45210 41060 45220
rect 40830 45140 40970 45210
rect 41040 45140 41060 45210
rect 40830 45130 41060 45140
rect 40740 45120 41060 45130
rect 41700 45220 42070 45230
rect 41700 45210 41980 45220
rect 41700 45140 41720 45210
rect 41790 45140 41980 45210
rect 41700 45130 41980 45140
rect 42060 45130 42070 45220
rect 41700 45120 42070 45130
rect 49940 45220 50260 45230
rect 49940 45130 49950 45220
rect 50030 45210 50260 45220
rect 50030 45140 50170 45210
rect 50240 45140 50260 45210
rect 50030 45130 50260 45140
rect 49940 45120 50260 45130
rect 50900 45220 51270 45230
rect 50900 45210 51180 45220
rect 50900 45140 50920 45210
rect 50990 45140 51180 45210
rect 50900 45130 51180 45140
rect 51260 45130 51270 45220
rect 50900 45120 51270 45130
rect 59140 45220 59460 45230
rect 59140 45130 59150 45220
rect 59230 45210 59460 45220
rect 59230 45140 59370 45210
rect 59440 45140 59460 45210
rect 59230 45130 59460 45140
rect 59140 45120 59460 45130
rect 60100 45220 60470 45230
rect 60100 45210 60380 45220
rect 60100 45140 60120 45210
rect 60190 45140 60380 45210
rect 60100 45130 60380 45140
rect 60460 45130 60470 45220
rect 60100 45120 60470 45130
rect 68340 45220 68660 45230
rect 68340 45130 68350 45220
rect 68430 45210 68660 45220
rect 68430 45140 68570 45210
rect 68640 45140 68660 45210
rect 68430 45130 68660 45140
rect 68340 45120 68660 45130
rect 69300 45220 69670 45230
rect 69300 45210 69580 45220
rect 69300 45140 69320 45210
rect 69390 45140 69580 45210
rect 69300 45130 69580 45140
rect 69660 45130 69670 45220
rect 69300 45120 69670 45130
rect 3085 36422 4044 36450
rect 3085 35618 3960 36422
rect 4024 35618 4044 36422
rect 3085 35590 4044 35618
rect 5164 36422 6123 36450
rect 5164 35618 5184 36422
rect 5248 35618 6123 36422
rect 5164 35590 6123 35618
rect 12285 36422 13244 36450
rect 12285 35618 13160 36422
rect 13224 35618 13244 36422
rect 12285 35590 13244 35618
rect 14364 36422 15323 36450
rect 14364 35618 14384 36422
rect 14448 35618 15323 36422
rect 14364 35590 15323 35618
rect 21485 36422 22444 36450
rect 21485 35618 22360 36422
rect 22424 35618 22444 36422
rect 21485 35590 22444 35618
rect 23564 36422 24523 36450
rect 23564 35618 23584 36422
rect 23648 35618 24523 36422
rect 23564 35590 24523 35618
rect 30685 36422 31644 36450
rect 30685 35618 31560 36422
rect 31624 35618 31644 36422
rect 30685 35590 31644 35618
rect 32764 36422 33723 36450
rect 32764 35618 32784 36422
rect 32848 35618 33723 36422
rect 32764 35590 33723 35618
rect 39885 36422 40844 36450
rect 39885 35618 40760 36422
rect 40824 35618 40844 36422
rect 39885 35590 40844 35618
rect 41964 36422 42923 36450
rect 41964 35618 41984 36422
rect 42048 35618 42923 36422
rect 41964 35590 42923 35618
rect 49085 36422 50044 36450
rect 49085 35618 49960 36422
rect 50024 35618 50044 36422
rect 49085 35590 50044 35618
rect 51164 36422 52123 36450
rect 51164 35618 51184 36422
rect 51248 35618 52123 36422
rect 51164 35590 52123 35618
rect 58285 36422 59244 36450
rect 58285 35618 59160 36422
rect 59224 35618 59244 36422
rect 58285 35590 59244 35618
rect 60364 36422 61323 36450
rect 60364 35618 60384 36422
rect 60448 35618 61323 36422
rect 60364 35590 61323 35618
rect 67485 36422 68444 36450
rect 67485 35618 68360 36422
rect 68424 35618 68444 36422
rect 67485 35590 68444 35618
rect 69564 36422 70523 36450
rect 69564 35618 69584 36422
rect 69648 35618 70523 36422
rect 69564 35590 70523 35618
rect 3940 35340 4260 35350
rect 3940 35250 3950 35340
rect 4030 35330 4260 35340
rect 4030 35260 4170 35330
rect 4240 35260 4260 35330
rect 4030 35250 4260 35260
rect 3940 35240 4260 35250
rect 4900 35340 5270 35350
rect 4900 35330 5180 35340
rect 4900 35260 4920 35330
rect 4990 35260 5180 35330
rect 4900 35250 5180 35260
rect 5260 35250 5270 35340
rect 4900 35240 5270 35250
rect 13140 35340 13460 35350
rect 13140 35250 13150 35340
rect 13230 35330 13460 35340
rect 13230 35260 13370 35330
rect 13440 35260 13460 35330
rect 13230 35250 13460 35260
rect 13140 35240 13460 35250
rect 14100 35340 14470 35350
rect 14100 35330 14380 35340
rect 14100 35260 14120 35330
rect 14190 35260 14380 35330
rect 14100 35250 14380 35260
rect 14460 35250 14470 35340
rect 14100 35240 14470 35250
rect 22340 35340 22660 35350
rect 22340 35250 22350 35340
rect 22430 35330 22660 35340
rect 22430 35260 22570 35330
rect 22640 35260 22660 35330
rect 22430 35250 22660 35260
rect 22340 35240 22660 35250
rect 23300 35340 23670 35350
rect 23300 35330 23580 35340
rect 23300 35260 23320 35330
rect 23390 35260 23580 35330
rect 23300 35250 23580 35260
rect 23660 35250 23670 35340
rect 23300 35240 23670 35250
rect 31540 35340 31860 35350
rect 31540 35250 31550 35340
rect 31630 35330 31860 35340
rect 31630 35260 31770 35330
rect 31840 35260 31860 35330
rect 31630 35250 31860 35260
rect 31540 35240 31860 35250
rect 32500 35340 32870 35350
rect 32500 35330 32780 35340
rect 32500 35260 32520 35330
rect 32590 35260 32780 35330
rect 32500 35250 32780 35260
rect 32860 35250 32870 35340
rect 32500 35240 32870 35250
rect 40740 35340 41060 35350
rect 40740 35250 40750 35340
rect 40830 35330 41060 35340
rect 40830 35260 40970 35330
rect 41040 35260 41060 35330
rect 40830 35250 41060 35260
rect 40740 35240 41060 35250
rect 41700 35340 42070 35350
rect 41700 35330 41980 35340
rect 41700 35260 41720 35330
rect 41790 35260 41980 35330
rect 41700 35250 41980 35260
rect 42060 35250 42070 35340
rect 41700 35240 42070 35250
rect 49940 35340 50260 35350
rect 49940 35250 49950 35340
rect 50030 35330 50260 35340
rect 50030 35260 50170 35330
rect 50240 35260 50260 35330
rect 50030 35250 50260 35260
rect 49940 35240 50260 35250
rect 50900 35340 51270 35350
rect 50900 35330 51180 35340
rect 50900 35260 50920 35330
rect 50990 35260 51180 35330
rect 50900 35250 51180 35260
rect 51260 35250 51270 35340
rect 50900 35240 51270 35250
rect 59140 35340 59460 35350
rect 59140 35250 59150 35340
rect 59230 35330 59460 35340
rect 59230 35260 59370 35330
rect 59440 35260 59460 35330
rect 59230 35250 59460 35260
rect 59140 35240 59460 35250
rect 60100 35340 60470 35350
rect 60100 35330 60380 35340
rect 60100 35260 60120 35330
rect 60190 35260 60380 35330
rect 60100 35250 60380 35260
rect 60460 35250 60470 35340
rect 60100 35240 60470 35250
rect 68340 35340 68660 35350
rect 68340 35250 68350 35340
rect 68430 35330 68660 35340
rect 68430 35260 68570 35330
rect 68640 35260 68660 35330
rect 68430 35250 68660 35260
rect 68340 35240 68660 35250
rect 69300 35340 69670 35350
rect 69300 35330 69580 35340
rect 69300 35260 69320 35330
rect 69390 35260 69580 35330
rect 69300 35250 69580 35260
rect 69660 35250 69670 35340
rect 69300 35240 69670 35250
rect 3085 26542 4044 26570
rect 3085 25738 3960 26542
rect 4024 25738 4044 26542
rect 3085 25710 4044 25738
rect 5164 26542 6123 26570
rect 5164 25738 5184 26542
rect 5248 25738 6123 26542
rect 5164 25710 6123 25738
rect 12285 26542 13244 26570
rect 12285 25738 13160 26542
rect 13224 25738 13244 26542
rect 12285 25710 13244 25738
rect 14364 26542 15323 26570
rect 14364 25738 14384 26542
rect 14448 25738 15323 26542
rect 14364 25710 15323 25738
rect 21485 26542 22444 26570
rect 21485 25738 22360 26542
rect 22424 25738 22444 26542
rect 21485 25710 22444 25738
rect 23564 26542 24523 26570
rect 23564 25738 23584 26542
rect 23648 25738 24523 26542
rect 23564 25710 24523 25738
rect 30685 26542 31644 26570
rect 30685 25738 31560 26542
rect 31624 25738 31644 26542
rect 30685 25710 31644 25738
rect 32764 26542 33723 26570
rect 32764 25738 32784 26542
rect 32848 25738 33723 26542
rect 32764 25710 33723 25738
rect 39885 26542 40844 26570
rect 39885 25738 40760 26542
rect 40824 25738 40844 26542
rect 39885 25710 40844 25738
rect 41964 26542 42923 26570
rect 41964 25738 41984 26542
rect 42048 25738 42923 26542
rect 41964 25710 42923 25738
rect 49085 26542 50044 26570
rect 49085 25738 49960 26542
rect 50024 25738 50044 26542
rect 49085 25710 50044 25738
rect 51164 26542 52123 26570
rect 51164 25738 51184 26542
rect 51248 25738 52123 26542
rect 51164 25710 52123 25738
rect 58285 26542 59244 26570
rect 58285 25738 59160 26542
rect 59224 25738 59244 26542
rect 58285 25710 59244 25738
rect 60364 26542 61323 26570
rect 60364 25738 60384 26542
rect 60448 25738 61323 26542
rect 60364 25710 61323 25738
rect 67485 26542 68444 26570
rect 67485 25738 68360 26542
rect 68424 25738 68444 26542
rect 67485 25710 68444 25738
rect 69564 26542 70523 26570
rect 69564 25738 69584 26542
rect 69648 25738 70523 26542
rect 69564 25710 70523 25738
rect 3940 25460 4260 25470
rect 3940 25370 3950 25460
rect 4030 25450 4260 25460
rect 4030 25380 4170 25450
rect 4240 25380 4260 25450
rect 4030 25370 4260 25380
rect 3940 25360 4260 25370
rect 4900 25460 5270 25470
rect 4900 25450 5180 25460
rect 4900 25380 4920 25450
rect 4990 25380 5180 25450
rect 4900 25370 5180 25380
rect 5260 25370 5270 25460
rect 4900 25360 5270 25370
rect 13140 25460 13460 25470
rect 13140 25370 13150 25460
rect 13230 25450 13460 25460
rect 13230 25380 13370 25450
rect 13440 25380 13460 25450
rect 13230 25370 13460 25380
rect 13140 25360 13460 25370
rect 14100 25460 14470 25470
rect 14100 25450 14380 25460
rect 14100 25380 14120 25450
rect 14190 25380 14380 25450
rect 14100 25370 14380 25380
rect 14460 25370 14470 25460
rect 14100 25360 14470 25370
rect 22340 25460 22660 25470
rect 22340 25370 22350 25460
rect 22430 25450 22660 25460
rect 22430 25380 22570 25450
rect 22640 25380 22660 25450
rect 22430 25370 22660 25380
rect 22340 25360 22660 25370
rect 23300 25460 23670 25470
rect 23300 25450 23580 25460
rect 23300 25380 23320 25450
rect 23390 25380 23580 25450
rect 23300 25370 23580 25380
rect 23660 25370 23670 25460
rect 23300 25360 23670 25370
rect 31540 25460 31860 25470
rect 31540 25370 31550 25460
rect 31630 25450 31860 25460
rect 31630 25380 31770 25450
rect 31840 25380 31860 25450
rect 31630 25370 31860 25380
rect 31540 25360 31860 25370
rect 32500 25460 32870 25470
rect 32500 25450 32780 25460
rect 32500 25380 32520 25450
rect 32590 25380 32780 25450
rect 32500 25370 32780 25380
rect 32860 25370 32870 25460
rect 32500 25360 32870 25370
rect 40740 25460 41060 25470
rect 40740 25370 40750 25460
rect 40830 25450 41060 25460
rect 40830 25380 40970 25450
rect 41040 25380 41060 25450
rect 40830 25370 41060 25380
rect 40740 25360 41060 25370
rect 41700 25460 42070 25470
rect 41700 25450 41980 25460
rect 41700 25380 41720 25450
rect 41790 25380 41980 25450
rect 41700 25370 41980 25380
rect 42060 25370 42070 25460
rect 41700 25360 42070 25370
rect 49940 25460 50260 25470
rect 49940 25370 49950 25460
rect 50030 25450 50260 25460
rect 50030 25380 50170 25450
rect 50240 25380 50260 25450
rect 50030 25370 50260 25380
rect 49940 25360 50260 25370
rect 50900 25460 51270 25470
rect 50900 25450 51180 25460
rect 50900 25380 50920 25450
rect 50990 25380 51180 25450
rect 50900 25370 51180 25380
rect 51260 25370 51270 25460
rect 50900 25360 51270 25370
rect 59140 25460 59460 25470
rect 59140 25370 59150 25460
rect 59230 25450 59460 25460
rect 59230 25380 59370 25450
rect 59440 25380 59460 25450
rect 59230 25370 59460 25380
rect 59140 25360 59460 25370
rect 60100 25460 60470 25470
rect 60100 25450 60380 25460
rect 60100 25380 60120 25450
rect 60190 25380 60380 25450
rect 60100 25370 60380 25380
rect 60460 25370 60470 25460
rect 60100 25360 60470 25370
rect 68340 25460 68660 25470
rect 68340 25370 68350 25460
rect 68430 25450 68660 25460
rect 68430 25380 68570 25450
rect 68640 25380 68660 25450
rect 68430 25370 68660 25380
rect 68340 25360 68660 25370
rect 69300 25460 69670 25470
rect 69300 25450 69580 25460
rect 69300 25380 69320 25450
rect 69390 25380 69580 25450
rect 69300 25370 69580 25380
rect 69660 25370 69670 25460
rect 69300 25360 69670 25370
rect 3085 16662 4044 16690
rect 3085 15858 3960 16662
rect 4024 15858 4044 16662
rect 3085 15830 4044 15858
rect 5164 16662 6123 16690
rect 5164 15858 5184 16662
rect 5248 15858 6123 16662
rect 5164 15830 6123 15858
rect 12285 16662 13244 16690
rect 12285 15858 13160 16662
rect 13224 15858 13244 16662
rect 12285 15830 13244 15858
rect 14364 16662 15323 16690
rect 14364 15858 14384 16662
rect 14448 15858 15323 16662
rect 14364 15830 15323 15858
rect 21485 16662 22444 16690
rect 21485 15858 22360 16662
rect 22424 15858 22444 16662
rect 21485 15830 22444 15858
rect 23564 16662 24523 16690
rect 23564 15858 23584 16662
rect 23648 15858 24523 16662
rect 23564 15830 24523 15858
rect 30685 16662 31644 16690
rect 30685 15858 31560 16662
rect 31624 15858 31644 16662
rect 30685 15830 31644 15858
rect 32764 16662 33723 16690
rect 32764 15858 32784 16662
rect 32848 15858 33723 16662
rect 32764 15830 33723 15858
rect 39885 16662 40844 16690
rect 39885 15858 40760 16662
rect 40824 15858 40844 16662
rect 39885 15830 40844 15858
rect 41964 16662 42923 16690
rect 41964 15858 41984 16662
rect 42048 15858 42923 16662
rect 41964 15830 42923 15858
rect 49085 16662 50044 16690
rect 49085 15858 49960 16662
rect 50024 15858 50044 16662
rect 49085 15830 50044 15858
rect 51164 16662 52123 16690
rect 51164 15858 51184 16662
rect 51248 15858 52123 16662
rect 51164 15830 52123 15858
rect 58285 16662 59244 16690
rect 58285 15858 59160 16662
rect 59224 15858 59244 16662
rect 58285 15830 59244 15858
rect 60364 16662 61323 16690
rect 60364 15858 60384 16662
rect 60448 15858 61323 16662
rect 60364 15830 61323 15858
rect 67485 16662 68444 16690
rect 67485 15858 68360 16662
rect 68424 15858 68444 16662
rect 67485 15830 68444 15858
rect 69564 16662 70523 16690
rect 69564 15858 69584 16662
rect 69648 15858 70523 16662
rect 69564 15830 70523 15858
rect 3940 15580 4260 15590
rect 3940 15490 3950 15580
rect 4030 15570 4260 15580
rect 4030 15500 4170 15570
rect 4240 15500 4260 15570
rect 4030 15490 4260 15500
rect 3940 15480 4260 15490
rect 4900 15580 5270 15590
rect 4900 15570 5180 15580
rect 4900 15500 4920 15570
rect 4990 15500 5180 15570
rect 4900 15490 5180 15500
rect 5260 15490 5270 15580
rect 4900 15480 5270 15490
rect 13140 15580 13460 15590
rect 13140 15490 13150 15580
rect 13230 15570 13460 15580
rect 13230 15500 13370 15570
rect 13440 15500 13460 15570
rect 13230 15490 13460 15500
rect 13140 15480 13460 15490
rect 14100 15580 14470 15590
rect 14100 15570 14380 15580
rect 14100 15500 14120 15570
rect 14190 15500 14380 15570
rect 14100 15490 14380 15500
rect 14460 15490 14470 15580
rect 14100 15480 14470 15490
rect 22340 15580 22660 15590
rect 22340 15490 22350 15580
rect 22430 15570 22660 15580
rect 22430 15500 22570 15570
rect 22640 15500 22660 15570
rect 22430 15490 22660 15500
rect 22340 15480 22660 15490
rect 23300 15580 23670 15590
rect 23300 15570 23580 15580
rect 23300 15500 23320 15570
rect 23390 15500 23580 15570
rect 23300 15490 23580 15500
rect 23660 15490 23670 15580
rect 23300 15480 23670 15490
rect 31540 15580 31860 15590
rect 31540 15490 31550 15580
rect 31630 15570 31860 15580
rect 31630 15500 31770 15570
rect 31840 15500 31860 15570
rect 31630 15490 31860 15500
rect 31540 15480 31860 15490
rect 32500 15580 32870 15590
rect 32500 15570 32780 15580
rect 32500 15500 32520 15570
rect 32590 15500 32780 15570
rect 32500 15490 32780 15500
rect 32860 15490 32870 15580
rect 32500 15480 32870 15490
rect 40740 15580 41060 15590
rect 40740 15490 40750 15580
rect 40830 15570 41060 15580
rect 40830 15500 40970 15570
rect 41040 15500 41060 15570
rect 40830 15490 41060 15500
rect 40740 15480 41060 15490
rect 41700 15580 42070 15590
rect 41700 15570 41980 15580
rect 41700 15500 41720 15570
rect 41790 15500 41980 15570
rect 41700 15490 41980 15500
rect 42060 15490 42070 15580
rect 41700 15480 42070 15490
rect 49940 15580 50260 15590
rect 49940 15490 49950 15580
rect 50030 15570 50260 15580
rect 50030 15500 50170 15570
rect 50240 15500 50260 15570
rect 50030 15490 50260 15500
rect 49940 15480 50260 15490
rect 50900 15580 51270 15590
rect 50900 15570 51180 15580
rect 50900 15500 50920 15570
rect 50990 15500 51180 15570
rect 50900 15490 51180 15500
rect 51260 15490 51270 15580
rect 50900 15480 51270 15490
rect 59140 15580 59460 15590
rect 59140 15490 59150 15580
rect 59230 15570 59460 15580
rect 59230 15500 59370 15570
rect 59440 15500 59460 15570
rect 59230 15490 59460 15500
rect 59140 15480 59460 15490
rect 60100 15580 60470 15590
rect 60100 15570 60380 15580
rect 60100 15500 60120 15570
rect 60190 15500 60380 15570
rect 60100 15490 60380 15500
rect 60460 15490 60470 15580
rect 60100 15480 60470 15490
rect 68340 15580 68660 15590
rect 68340 15490 68350 15580
rect 68430 15570 68660 15580
rect 68430 15500 68570 15570
rect 68640 15500 68660 15570
rect 68430 15490 68660 15500
rect 68340 15480 68660 15490
rect 69300 15580 69670 15590
rect 69300 15570 69580 15580
rect 69300 15500 69320 15570
rect 69390 15500 69580 15570
rect 69300 15490 69580 15500
rect 69660 15490 69670 15580
rect 69300 15480 69670 15490
rect 3085 6782 4044 6810
rect 3085 5978 3960 6782
rect 4024 5978 4044 6782
rect 3085 5950 4044 5978
rect 5164 6782 6123 6810
rect 5164 5978 5184 6782
rect 5248 5978 6123 6782
rect 5164 5950 6123 5978
rect 12285 6782 13244 6810
rect 12285 5978 13160 6782
rect 13224 5978 13244 6782
rect 12285 5950 13244 5978
rect 14364 6782 15323 6810
rect 14364 5978 14384 6782
rect 14448 5978 15323 6782
rect 14364 5950 15323 5978
rect 21485 6782 22444 6810
rect 21485 5978 22360 6782
rect 22424 5978 22444 6782
rect 21485 5950 22444 5978
rect 23564 6782 24523 6810
rect 23564 5978 23584 6782
rect 23648 5978 24523 6782
rect 23564 5950 24523 5978
rect 30685 6782 31644 6810
rect 30685 5978 31560 6782
rect 31624 5978 31644 6782
rect 30685 5950 31644 5978
rect 32764 6782 33723 6810
rect 32764 5978 32784 6782
rect 32848 5978 33723 6782
rect 32764 5950 33723 5978
rect 39885 6782 40844 6810
rect 39885 5978 40760 6782
rect 40824 5978 40844 6782
rect 39885 5950 40844 5978
rect 41964 6782 42923 6810
rect 41964 5978 41984 6782
rect 42048 5978 42923 6782
rect 41964 5950 42923 5978
rect 49085 6782 50044 6810
rect 49085 5978 49960 6782
rect 50024 5978 50044 6782
rect 49085 5950 50044 5978
rect 51164 6782 52123 6810
rect 51164 5978 51184 6782
rect 51248 5978 52123 6782
rect 51164 5950 52123 5978
rect 58285 6782 59244 6810
rect 58285 5978 59160 6782
rect 59224 5978 59244 6782
rect 58285 5950 59244 5978
rect 60364 6782 61323 6810
rect 60364 5978 60384 6782
rect 60448 5978 61323 6782
rect 60364 5950 61323 5978
rect 67485 6782 68444 6810
rect 67485 5978 68360 6782
rect 68424 5978 68444 6782
rect 67485 5950 68444 5978
rect 69564 6782 70523 6810
rect 69564 5978 69584 6782
rect 69648 5978 70523 6782
rect 69564 5950 70523 5978
rect 3940 5700 4260 5710
rect 3940 5610 3950 5700
rect 4030 5690 4260 5700
rect 4030 5620 4170 5690
rect 4240 5620 4260 5690
rect 4030 5610 4260 5620
rect 3940 5600 4260 5610
rect 4900 5700 5270 5710
rect 4900 5690 5180 5700
rect 4900 5620 4920 5690
rect 4990 5620 5180 5690
rect 4900 5610 5180 5620
rect 5260 5610 5270 5700
rect 4900 5600 5270 5610
rect 13140 5700 13460 5710
rect 13140 5610 13150 5700
rect 13230 5690 13460 5700
rect 13230 5620 13370 5690
rect 13440 5620 13460 5690
rect 13230 5610 13460 5620
rect 13140 5600 13460 5610
rect 14100 5700 14470 5710
rect 14100 5690 14380 5700
rect 14100 5620 14120 5690
rect 14190 5620 14380 5690
rect 14100 5610 14380 5620
rect 14460 5610 14470 5700
rect 14100 5600 14470 5610
rect 22340 5700 22660 5710
rect 22340 5610 22350 5700
rect 22430 5690 22660 5700
rect 22430 5620 22570 5690
rect 22640 5620 22660 5690
rect 22430 5610 22660 5620
rect 22340 5600 22660 5610
rect 23300 5700 23670 5710
rect 23300 5690 23580 5700
rect 23300 5620 23320 5690
rect 23390 5620 23580 5690
rect 23300 5610 23580 5620
rect 23660 5610 23670 5700
rect 23300 5600 23670 5610
rect 31540 5700 31860 5710
rect 31540 5610 31550 5700
rect 31630 5690 31860 5700
rect 31630 5620 31770 5690
rect 31840 5620 31860 5690
rect 31630 5610 31860 5620
rect 31540 5600 31860 5610
rect 32500 5700 32870 5710
rect 32500 5690 32780 5700
rect 32500 5620 32520 5690
rect 32590 5620 32780 5690
rect 32500 5610 32780 5620
rect 32860 5610 32870 5700
rect 32500 5600 32870 5610
rect 40740 5700 41060 5710
rect 40740 5610 40750 5700
rect 40830 5690 41060 5700
rect 40830 5620 40970 5690
rect 41040 5620 41060 5690
rect 40830 5610 41060 5620
rect 40740 5600 41060 5610
rect 41700 5700 42070 5710
rect 41700 5690 41980 5700
rect 41700 5620 41720 5690
rect 41790 5620 41980 5690
rect 41700 5610 41980 5620
rect 42060 5610 42070 5700
rect 41700 5600 42070 5610
rect 49940 5700 50260 5710
rect 49940 5610 49950 5700
rect 50030 5690 50260 5700
rect 50030 5620 50170 5690
rect 50240 5620 50260 5690
rect 50030 5610 50260 5620
rect 49940 5600 50260 5610
rect 50900 5700 51270 5710
rect 50900 5690 51180 5700
rect 50900 5620 50920 5690
rect 50990 5620 51180 5690
rect 50900 5610 51180 5620
rect 51260 5610 51270 5700
rect 50900 5600 51270 5610
rect 59140 5700 59460 5710
rect 59140 5610 59150 5700
rect 59230 5690 59460 5700
rect 59230 5620 59370 5690
rect 59440 5620 59460 5690
rect 59230 5610 59460 5620
rect 59140 5600 59460 5610
rect 60100 5700 60470 5710
rect 60100 5690 60380 5700
rect 60100 5620 60120 5690
rect 60190 5620 60380 5690
rect 60100 5610 60380 5620
rect 60460 5610 60470 5700
rect 60100 5600 60470 5610
rect 68340 5700 68660 5710
rect 68340 5610 68350 5700
rect 68430 5690 68660 5700
rect 68430 5620 68570 5690
rect 68640 5620 68660 5690
rect 68430 5610 68660 5620
rect 68340 5600 68660 5610
rect 69300 5700 69670 5710
rect 69300 5690 69580 5700
rect 69300 5620 69320 5690
rect 69390 5620 69580 5690
rect 69300 5610 69580 5620
rect 69660 5610 69670 5700
rect 69300 5600 69670 5610
<< via3 >>
rect 6220 107810 8200 109790
rect 15420 107810 17400 109790
rect 24620 107810 26600 109790
rect 33820 107810 35800 109790
rect 43020 107810 45000 109790
rect 52220 107810 54200 109790
rect 61420 107800 63400 109780
rect 70620 107800 72600 109780
rect 1010 101800 2990 103780
rect 10210 101800 12190 103780
rect 19410 101800 21390 103780
rect 28610 101800 30590 103780
rect 37810 101800 39790 103780
rect 47010 101800 48990 103780
rect 56210 101800 58190 103780
rect 65410 101800 67390 103780
rect 3960 94898 4024 95702
rect 5184 94898 5248 95702
rect 3950 94530 4030 94620
rect 5180 94530 5260 94620
rect 3960 85018 4024 85822
rect 5184 85018 5248 85822
rect 13160 85018 13224 85822
rect 14384 85018 14448 85822
rect 3950 84650 4030 84740
rect 5180 84650 5260 84740
rect 13150 84650 13230 84740
rect 14380 84650 14460 84740
rect 3960 75138 4024 75942
rect 5184 75138 5248 75942
rect 13160 75138 13224 75942
rect 14384 75138 14448 75942
rect 22360 75138 22424 75942
rect 23584 75138 23648 75942
rect 31560 75138 31624 75942
rect 32784 75138 32848 75942
rect 3950 74770 4030 74860
rect 5180 74770 5260 74860
rect 13150 74770 13230 74860
rect 14380 74770 14460 74860
rect 22350 74770 22430 74860
rect 23580 74770 23660 74860
rect 31550 74770 31630 74860
rect 32780 74770 32860 74860
rect 3960 65258 4024 66062
rect 5184 65258 5248 66062
rect 13160 65258 13224 66062
rect 14384 65258 14448 66062
rect 22360 65258 22424 66062
rect 23584 65258 23648 66062
rect 31560 65258 31624 66062
rect 32784 65258 32848 66062
rect 40760 65258 40824 66062
rect 41984 65258 42048 66062
rect 49960 65258 50024 66062
rect 51184 65258 51248 66062
rect 59160 65258 59224 66062
rect 60384 65258 60448 66062
rect 68360 65258 68424 66062
rect 69584 65258 69648 66062
rect 3950 64890 4030 64980
rect 5180 64890 5260 64980
rect 13150 64890 13230 64980
rect 14380 64890 14460 64980
rect 22350 64890 22430 64980
rect 23580 64890 23660 64980
rect 31550 64890 31630 64980
rect 32780 64890 32860 64980
rect 40750 64890 40830 64980
rect 41980 64890 42060 64980
rect 49950 64890 50030 64980
rect 51180 64890 51260 64980
rect 59150 64890 59230 64980
rect 60380 64890 60460 64980
rect 68350 64890 68430 64980
rect 69580 64890 69660 64980
rect 3960 55378 4024 56182
rect 5184 55378 5248 56182
rect 13160 55378 13224 56182
rect 14384 55378 14448 56182
rect 22360 55378 22424 56182
rect 23584 55378 23648 56182
rect 31560 55378 31624 56182
rect 32784 55378 32848 56182
rect 40760 55378 40824 56182
rect 41984 55378 42048 56182
rect 49960 55378 50024 56182
rect 51184 55378 51248 56182
rect 59160 55378 59224 56182
rect 60384 55378 60448 56182
rect 68360 55378 68424 56182
rect 69584 55378 69648 56182
rect 3950 55010 4030 55100
rect 5180 55010 5260 55100
rect 13150 55010 13230 55100
rect 14380 55010 14460 55100
rect 22350 55010 22430 55100
rect 23580 55010 23660 55100
rect 31550 55010 31630 55100
rect 32780 55010 32860 55100
rect 40750 55010 40830 55100
rect 41980 55010 42060 55100
rect 49950 55010 50030 55100
rect 51180 55010 51260 55100
rect 59150 55010 59230 55100
rect 60380 55010 60460 55100
rect 68350 55010 68430 55100
rect 69580 55010 69660 55100
rect 3960 45498 4024 46302
rect 5184 45498 5248 46302
rect 13160 45498 13224 46302
rect 14384 45498 14448 46302
rect 22360 45498 22424 46302
rect 23584 45498 23648 46302
rect 31560 45498 31624 46302
rect 32784 45498 32848 46302
rect 40760 45498 40824 46302
rect 41984 45498 42048 46302
rect 49960 45498 50024 46302
rect 51184 45498 51248 46302
rect 59160 45498 59224 46302
rect 60384 45498 60448 46302
rect 68360 45498 68424 46302
rect 69584 45498 69648 46302
rect 3950 45130 4030 45220
rect 5180 45130 5260 45220
rect 13150 45130 13230 45220
rect 14380 45130 14460 45220
rect 22350 45130 22430 45220
rect 23580 45130 23660 45220
rect 31550 45130 31630 45220
rect 32780 45130 32860 45220
rect 40750 45130 40830 45220
rect 41980 45130 42060 45220
rect 49950 45130 50030 45220
rect 51180 45130 51260 45220
rect 59150 45130 59230 45220
rect 60380 45130 60460 45220
rect 68350 45130 68430 45220
rect 69580 45130 69660 45220
rect 3960 35618 4024 36422
rect 5184 35618 5248 36422
rect 13160 35618 13224 36422
rect 14384 35618 14448 36422
rect 22360 35618 22424 36422
rect 23584 35618 23648 36422
rect 31560 35618 31624 36422
rect 32784 35618 32848 36422
rect 40760 35618 40824 36422
rect 41984 35618 42048 36422
rect 49960 35618 50024 36422
rect 51184 35618 51248 36422
rect 59160 35618 59224 36422
rect 60384 35618 60448 36422
rect 68360 35618 68424 36422
rect 69584 35618 69648 36422
rect 3950 35250 4030 35340
rect 5180 35250 5260 35340
rect 13150 35250 13230 35340
rect 14380 35250 14460 35340
rect 22350 35250 22430 35340
rect 23580 35250 23660 35340
rect 31550 35250 31630 35340
rect 32780 35250 32860 35340
rect 40750 35250 40830 35340
rect 41980 35250 42060 35340
rect 49950 35250 50030 35340
rect 51180 35250 51260 35340
rect 59150 35250 59230 35340
rect 60380 35250 60460 35340
rect 68350 35250 68430 35340
rect 69580 35250 69660 35340
rect 3960 25738 4024 26542
rect 5184 25738 5248 26542
rect 13160 25738 13224 26542
rect 14384 25738 14448 26542
rect 22360 25738 22424 26542
rect 23584 25738 23648 26542
rect 31560 25738 31624 26542
rect 32784 25738 32848 26542
rect 40760 25738 40824 26542
rect 41984 25738 42048 26542
rect 49960 25738 50024 26542
rect 51184 25738 51248 26542
rect 59160 25738 59224 26542
rect 60384 25738 60448 26542
rect 68360 25738 68424 26542
rect 69584 25738 69648 26542
rect 3950 25370 4030 25460
rect 5180 25370 5260 25460
rect 13150 25370 13230 25460
rect 14380 25370 14460 25460
rect 22350 25370 22430 25460
rect 23580 25370 23660 25460
rect 31550 25370 31630 25460
rect 32780 25370 32860 25460
rect 40750 25370 40830 25460
rect 41980 25370 42060 25460
rect 49950 25370 50030 25460
rect 51180 25370 51260 25460
rect 59150 25370 59230 25460
rect 60380 25370 60460 25460
rect 68350 25370 68430 25460
rect 69580 25370 69660 25460
rect 3960 15858 4024 16662
rect 5184 15858 5248 16662
rect 13160 15858 13224 16662
rect 14384 15858 14448 16662
rect 22360 15858 22424 16662
rect 23584 15858 23648 16662
rect 31560 15858 31624 16662
rect 32784 15858 32848 16662
rect 40760 15858 40824 16662
rect 41984 15858 42048 16662
rect 49960 15858 50024 16662
rect 51184 15858 51248 16662
rect 59160 15858 59224 16662
rect 60384 15858 60448 16662
rect 68360 15858 68424 16662
rect 69584 15858 69648 16662
rect 3950 15490 4030 15580
rect 5180 15490 5260 15580
rect 13150 15490 13230 15580
rect 14380 15490 14460 15580
rect 22350 15490 22430 15580
rect 23580 15490 23660 15580
rect 31550 15490 31630 15580
rect 32780 15490 32860 15580
rect 40750 15490 40830 15580
rect 41980 15490 42060 15580
rect 49950 15490 50030 15580
rect 51180 15490 51260 15580
rect 59150 15490 59230 15580
rect 60380 15490 60460 15580
rect 68350 15490 68430 15580
rect 69580 15490 69660 15580
rect 3960 5978 4024 6782
rect 5184 5978 5248 6782
rect 13160 5978 13224 6782
rect 14384 5978 14448 6782
rect 22360 5978 22424 6782
rect 23584 5978 23648 6782
rect 31560 5978 31624 6782
rect 32784 5978 32848 6782
rect 40760 5978 40824 6782
rect 41984 5978 42048 6782
rect 49960 5978 50024 6782
rect 51184 5978 51248 6782
rect 59160 5978 59224 6782
rect 60384 5978 60448 6782
rect 68360 5978 68424 6782
rect 69584 5978 69648 6782
rect 3950 5610 4030 5700
rect 5180 5610 5260 5700
rect 13150 5610 13230 5700
rect 14380 5610 14460 5700
rect 22350 5610 22430 5700
rect 23580 5610 23660 5700
rect 31550 5610 31630 5700
rect 32780 5610 32860 5700
rect 40750 5610 40830 5700
rect 41980 5610 42060 5700
rect 49950 5610 50030 5700
rect 51180 5610 51260 5700
rect 59150 5610 59230 5700
rect 60380 5610 60460 5700
rect 68350 5610 68430 5700
rect 69580 5610 69660 5700
<< mimcap >>
rect 3185 95590 3845 95630
rect 3185 95010 3225 95590
rect 3805 95010 3845 95590
rect 3185 94970 3845 95010
rect 5363 95590 6023 95630
rect 5363 95010 5403 95590
rect 5983 95010 6023 95590
rect 5363 94970 6023 95010
rect 3185 85710 3845 85750
rect 3185 85130 3225 85710
rect 3805 85130 3845 85710
rect 3185 85090 3845 85130
rect 5363 85710 6023 85750
rect 5363 85130 5403 85710
rect 5983 85130 6023 85710
rect 5363 85090 6023 85130
rect 12385 85710 13045 85750
rect 12385 85130 12425 85710
rect 13005 85130 13045 85710
rect 12385 85090 13045 85130
rect 14563 85710 15223 85750
rect 14563 85130 14603 85710
rect 15183 85130 15223 85710
rect 14563 85090 15223 85130
rect 3185 75830 3845 75870
rect 3185 75250 3225 75830
rect 3805 75250 3845 75830
rect 3185 75210 3845 75250
rect 5363 75830 6023 75870
rect 5363 75250 5403 75830
rect 5983 75250 6023 75830
rect 5363 75210 6023 75250
rect 12385 75830 13045 75870
rect 12385 75250 12425 75830
rect 13005 75250 13045 75830
rect 12385 75210 13045 75250
rect 14563 75830 15223 75870
rect 14563 75250 14603 75830
rect 15183 75250 15223 75830
rect 14563 75210 15223 75250
rect 21585 75830 22245 75870
rect 21585 75250 21625 75830
rect 22205 75250 22245 75830
rect 21585 75210 22245 75250
rect 23763 75830 24423 75870
rect 23763 75250 23803 75830
rect 24383 75250 24423 75830
rect 23763 75210 24423 75250
rect 30785 75830 31445 75870
rect 30785 75250 30825 75830
rect 31405 75250 31445 75830
rect 30785 75210 31445 75250
rect 32963 75830 33623 75870
rect 32963 75250 33003 75830
rect 33583 75250 33623 75830
rect 32963 75210 33623 75250
rect 3185 65950 3845 65990
rect 3185 65370 3225 65950
rect 3805 65370 3845 65950
rect 3185 65330 3845 65370
rect 5363 65950 6023 65990
rect 5363 65370 5403 65950
rect 5983 65370 6023 65950
rect 5363 65330 6023 65370
rect 12385 65950 13045 65990
rect 12385 65370 12425 65950
rect 13005 65370 13045 65950
rect 12385 65330 13045 65370
rect 14563 65950 15223 65990
rect 14563 65370 14603 65950
rect 15183 65370 15223 65950
rect 14563 65330 15223 65370
rect 21585 65950 22245 65990
rect 21585 65370 21625 65950
rect 22205 65370 22245 65950
rect 21585 65330 22245 65370
rect 23763 65950 24423 65990
rect 23763 65370 23803 65950
rect 24383 65370 24423 65950
rect 23763 65330 24423 65370
rect 30785 65950 31445 65990
rect 30785 65370 30825 65950
rect 31405 65370 31445 65950
rect 30785 65330 31445 65370
rect 32963 65950 33623 65990
rect 32963 65370 33003 65950
rect 33583 65370 33623 65950
rect 32963 65330 33623 65370
rect 39985 65950 40645 65990
rect 39985 65370 40025 65950
rect 40605 65370 40645 65950
rect 39985 65330 40645 65370
rect 42163 65950 42823 65990
rect 42163 65370 42203 65950
rect 42783 65370 42823 65950
rect 42163 65330 42823 65370
rect 49185 65950 49845 65990
rect 49185 65370 49225 65950
rect 49805 65370 49845 65950
rect 49185 65330 49845 65370
rect 51363 65950 52023 65990
rect 51363 65370 51403 65950
rect 51983 65370 52023 65950
rect 51363 65330 52023 65370
rect 58385 65950 59045 65990
rect 58385 65370 58425 65950
rect 59005 65370 59045 65950
rect 58385 65330 59045 65370
rect 60563 65950 61223 65990
rect 60563 65370 60603 65950
rect 61183 65370 61223 65950
rect 60563 65330 61223 65370
rect 67585 65950 68245 65990
rect 67585 65370 67625 65950
rect 68205 65370 68245 65950
rect 67585 65330 68245 65370
rect 69763 65950 70423 65990
rect 69763 65370 69803 65950
rect 70383 65370 70423 65950
rect 69763 65330 70423 65370
rect 3185 56070 3845 56110
rect 3185 55490 3225 56070
rect 3805 55490 3845 56070
rect 3185 55450 3845 55490
rect 5363 56070 6023 56110
rect 5363 55490 5403 56070
rect 5983 55490 6023 56070
rect 5363 55450 6023 55490
rect 12385 56070 13045 56110
rect 12385 55490 12425 56070
rect 13005 55490 13045 56070
rect 12385 55450 13045 55490
rect 14563 56070 15223 56110
rect 14563 55490 14603 56070
rect 15183 55490 15223 56070
rect 14563 55450 15223 55490
rect 21585 56070 22245 56110
rect 21585 55490 21625 56070
rect 22205 55490 22245 56070
rect 21585 55450 22245 55490
rect 23763 56070 24423 56110
rect 23763 55490 23803 56070
rect 24383 55490 24423 56070
rect 23763 55450 24423 55490
rect 30785 56070 31445 56110
rect 30785 55490 30825 56070
rect 31405 55490 31445 56070
rect 30785 55450 31445 55490
rect 32963 56070 33623 56110
rect 32963 55490 33003 56070
rect 33583 55490 33623 56070
rect 32963 55450 33623 55490
rect 39985 56070 40645 56110
rect 39985 55490 40025 56070
rect 40605 55490 40645 56070
rect 39985 55450 40645 55490
rect 42163 56070 42823 56110
rect 42163 55490 42203 56070
rect 42783 55490 42823 56070
rect 42163 55450 42823 55490
rect 49185 56070 49845 56110
rect 49185 55490 49225 56070
rect 49805 55490 49845 56070
rect 49185 55450 49845 55490
rect 51363 56070 52023 56110
rect 51363 55490 51403 56070
rect 51983 55490 52023 56070
rect 51363 55450 52023 55490
rect 58385 56070 59045 56110
rect 58385 55490 58425 56070
rect 59005 55490 59045 56070
rect 58385 55450 59045 55490
rect 60563 56070 61223 56110
rect 60563 55490 60603 56070
rect 61183 55490 61223 56070
rect 60563 55450 61223 55490
rect 67585 56070 68245 56110
rect 67585 55490 67625 56070
rect 68205 55490 68245 56070
rect 67585 55450 68245 55490
rect 69763 56070 70423 56110
rect 69763 55490 69803 56070
rect 70383 55490 70423 56070
rect 69763 55450 70423 55490
rect 3185 46190 3845 46230
rect 3185 45610 3225 46190
rect 3805 45610 3845 46190
rect 3185 45570 3845 45610
rect 5363 46190 6023 46230
rect 5363 45610 5403 46190
rect 5983 45610 6023 46190
rect 5363 45570 6023 45610
rect 12385 46190 13045 46230
rect 12385 45610 12425 46190
rect 13005 45610 13045 46190
rect 12385 45570 13045 45610
rect 14563 46190 15223 46230
rect 14563 45610 14603 46190
rect 15183 45610 15223 46190
rect 14563 45570 15223 45610
rect 21585 46190 22245 46230
rect 21585 45610 21625 46190
rect 22205 45610 22245 46190
rect 21585 45570 22245 45610
rect 23763 46190 24423 46230
rect 23763 45610 23803 46190
rect 24383 45610 24423 46190
rect 23763 45570 24423 45610
rect 30785 46190 31445 46230
rect 30785 45610 30825 46190
rect 31405 45610 31445 46190
rect 30785 45570 31445 45610
rect 32963 46190 33623 46230
rect 32963 45610 33003 46190
rect 33583 45610 33623 46190
rect 32963 45570 33623 45610
rect 39985 46190 40645 46230
rect 39985 45610 40025 46190
rect 40605 45610 40645 46190
rect 39985 45570 40645 45610
rect 42163 46190 42823 46230
rect 42163 45610 42203 46190
rect 42783 45610 42823 46190
rect 42163 45570 42823 45610
rect 49185 46190 49845 46230
rect 49185 45610 49225 46190
rect 49805 45610 49845 46190
rect 49185 45570 49845 45610
rect 51363 46190 52023 46230
rect 51363 45610 51403 46190
rect 51983 45610 52023 46190
rect 51363 45570 52023 45610
rect 58385 46190 59045 46230
rect 58385 45610 58425 46190
rect 59005 45610 59045 46190
rect 58385 45570 59045 45610
rect 60563 46190 61223 46230
rect 60563 45610 60603 46190
rect 61183 45610 61223 46190
rect 60563 45570 61223 45610
rect 67585 46190 68245 46230
rect 67585 45610 67625 46190
rect 68205 45610 68245 46190
rect 67585 45570 68245 45610
rect 69763 46190 70423 46230
rect 69763 45610 69803 46190
rect 70383 45610 70423 46190
rect 69763 45570 70423 45610
rect 3185 36310 3845 36350
rect 3185 35730 3225 36310
rect 3805 35730 3845 36310
rect 3185 35690 3845 35730
rect 5363 36310 6023 36350
rect 5363 35730 5403 36310
rect 5983 35730 6023 36310
rect 5363 35690 6023 35730
rect 12385 36310 13045 36350
rect 12385 35730 12425 36310
rect 13005 35730 13045 36310
rect 12385 35690 13045 35730
rect 14563 36310 15223 36350
rect 14563 35730 14603 36310
rect 15183 35730 15223 36310
rect 14563 35690 15223 35730
rect 21585 36310 22245 36350
rect 21585 35730 21625 36310
rect 22205 35730 22245 36310
rect 21585 35690 22245 35730
rect 23763 36310 24423 36350
rect 23763 35730 23803 36310
rect 24383 35730 24423 36310
rect 23763 35690 24423 35730
rect 30785 36310 31445 36350
rect 30785 35730 30825 36310
rect 31405 35730 31445 36310
rect 30785 35690 31445 35730
rect 32963 36310 33623 36350
rect 32963 35730 33003 36310
rect 33583 35730 33623 36310
rect 32963 35690 33623 35730
rect 39985 36310 40645 36350
rect 39985 35730 40025 36310
rect 40605 35730 40645 36310
rect 39985 35690 40645 35730
rect 42163 36310 42823 36350
rect 42163 35730 42203 36310
rect 42783 35730 42823 36310
rect 42163 35690 42823 35730
rect 49185 36310 49845 36350
rect 49185 35730 49225 36310
rect 49805 35730 49845 36310
rect 49185 35690 49845 35730
rect 51363 36310 52023 36350
rect 51363 35730 51403 36310
rect 51983 35730 52023 36310
rect 51363 35690 52023 35730
rect 58385 36310 59045 36350
rect 58385 35730 58425 36310
rect 59005 35730 59045 36310
rect 58385 35690 59045 35730
rect 60563 36310 61223 36350
rect 60563 35730 60603 36310
rect 61183 35730 61223 36310
rect 60563 35690 61223 35730
rect 67585 36310 68245 36350
rect 67585 35730 67625 36310
rect 68205 35730 68245 36310
rect 67585 35690 68245 35730
rect 69763 36310 70423 36350
rect 69763 35730 69803 36310
rect 70383 35730 70423 36310
rect 69763 35690 70423 35730
rect 3185 26430 3845 26470
rect 3185 25850 3225 26430
rect 3805 25850 3845 26430
rect 3185 25810 3845 25850
rect 5363 26430 6023 26470
rect 5363 25850 5403 26430
rect 5983 25850 6023 26430
rect 5363 25810 6023 25850
rect 12385 26430 13045 26470
rect 12385 25850 12425 26430
rect 13005 25850 13045 26430
rect 12385 25810 13045 25850
rect 14563 26430 15223 26470
rect 14563 25850 14603 26430
rect 15183 25850 15223 26430
rect 14563 25810 15223 25850
rect 21585 26430 22245 26470
rect 21585 25850 21625 26430
rect 22205 25850 22245 26430
rect 21585 25810 22245 25850
rect 23763 26430 24423 26470
rect 23763 25850 23803 26430
rect 24383 25850 24423 26430
rect 23763 25810 24423 25850
rect 30785 26430 31445 26470
rect 30785 25850 30825 26430
rect 31405 25850 31445 26430
rect 30785 25810 31445 25850
rect 32963 26430 33623 26470
rect 32963 25850 33003 26430
rect 33583 25850 33623 26430
rect 32963 25810 33623 25850
rect 39985 26430 40645 26470
rect 39985 25850 40025 26430
rect 40605 25850 40645 26430
rect 39985 25810 40645 25850
rect 42163 26430 42823 26470
rect 42163 25850 42203 26430
rect 42783 25850 42823 26430
rect 42163 25810 42823 25850
rect 49185 26430 49845 26470
rect 49185 25850 49225 26430
rect 49805 25850 49845 26430
rect 49185 25810 49845 25850
rect 51363 26430 52023 26470
rect 51363 25850 51403 26430
rect 51983 25850 52023 26430
rect 51363 25810 52023 25850
rect 58385 26430 59045 26470
rect 58385 25850 58425 26430
rect 59005 25850 59045 26430
rect 58385 25810 59045 25850
rect 60563 26430 61223 26470
rect 60563 25850 60603 26430
rect 61183 25850 61223 26430
rect 60563 25810 61223 25850
rect 67585 26430 68245 26470
rect 67585 25850 67625 26430
rect 68205 25850 68245 26430
rect 67585 25810 68245 25850
rect 69763 26430 70423 26470
rect 69763 25850 69803 26430
rect 70383 25850 70423 26430
rect 69763 25810 70423 25850
rect 3185 16550 3845 16590
rect 3185 15970 3225 16550
rect 3805 15970 3845 16550
rect 3185 15930 3845 15970
rect 5363 16550 6023 16590
rect 5363 15970 5403 16550
rect 5983 15970 6023 16550
rect 5363 15930 6023 15970
rect 12385 16550 13045 16590
rect 12385 15970 12425 16550
rect 13005 15970 13045 16550
rect 12385 15930 13045 15970
rect 14563 16550 15223 16590
rect 14563 15970 14603 16550
rect 15183 15970 15223 16550
rect 14563 15930 15223 15970
rect 21585 16550 22245 16590
rect 21585 15970 21625 16550
rect 22205 15970 22245 16550
rect 21585 15930 22245 15970
rect 23763 16550 24423 16590
rect 23763 15970 23803 16550
rect 24383 15970 24423 16550
rect 23763 15930 24423 15970
rect 30785 16550 31445 16590
rect 30785 15970 30825 16550
rect 31405 15970 31445 16550
rect 30785 15930 31445 15970
rect 32963 16550 33623 16590
rect 32963 15970 33003 16550
rect 33583 15970 33623 16550
rect 32963 15930 33623 15970
rect 39985 16550 40645 16590
rect 39985 15970 40025 16550
rect 40605 15970 40645 16550
rect 39985 15930 40645 15970
rect 42163 16550 42823 16590
rect 42163 15970 42203 16550
rect 42783 15970 42823 16550
rect 42163 15930 42823 15970
rect 49185 16550 49845 16590
rect 49185 15970 49225 16550
rect 49805 15970 49845 16550
rect 49185 15930 49845 15970
rect 51363 16550 52023 16590
rect 51363 15970 51403 16550
rect 51983 15970 52023 16550
rect 51363 15930 52023 15970
rect 58385 16550 59045 16590
rect 58385 15970 58425 16550
rect 59005 15970 59045 16550
rect 58385 15930 59045 15970
rect 60563 16550 61223 16590
rect 60563 15970 60603 16550
rect 61183 15970 61223 16550
rect 60563 15930 61223 15970
rect 67585 16550 68245 16590
rect 67585 15970 67625 16550
rect 68205 15970 68245 16550
rect 67585 15930 68245 15970
rect 69763 16550 70423 16590
rect 69763 15970 69803 16550
rect 70383 15970 70423 16550
rect 69763 15930 70423 15970
rect 3185 6670 3845 6710
rect 3185 6090 3225 6670
rect 3805 6090 3845 6670
rect 3185 6050 3845 6090
rect 5363 6670 6023 6710
rect 5363 6090 5403 6670
rect 5983 6090 6023 6670
rect 5363 6050 6023 6090
rect 12385 6670 13045 6710
rect 12385 6090 12425 6670
rect 13005 6090 13045 6670
rect 12385 6050 13045 6090
rect 14563 6670 15223 6710
rect 14563 6090 14603 6670
rect 15183 6090 15223 6670
rect 14563 6050 15223 6090
rect 21585 6670 22245 6710
rect 21585 6090 21625 6670
rect 22205 6090 22245 6670
rect 21585 6050 22245 6090
rect 23763 6670 24423 6710
rect 23763 6090 23803 6670
rect 24383 6090 24423 6670
rect 23763 6050 24423 6090
rect 30785 6670 31445 6710
rect 30785 6090 30825 6670
rect 31405 6090 31445 6670
rect 30785 6050 31445 6090
rect 32963 6670 33623 6710
rect 32963 6090 33003 6670
rect 33583 6090 33623 6670
rect 32963 6050 33623 6090
rect 39985 6670 40645 6710
rect 39985 6090 40025 6670
rect 40605 6090 40645 6670
rect 39985 6050 40645 6090
rect 42163 6670 42823 6710
rect 42163 6090 42203 6670
rect 42783 6090 42823 6670
rect 42163 6050 42823 6090
rect 49185 6670 49845 6710
rect 49185 6090 49225 6670
rect 49805 6090 49845 6670
rect 49185 6050 49845 6090
rect 51363 6670 52023 6710
rect 51363 6090 51403 6670
rect 51983 6090 52023 6670
rect 51363 6050 52023 6090
rect 58385 6670 59045 6710
rect 58385 6090 58425 6670
rect 59005 6090 59045 6670
rect 58385 6050 59045 6090
rect 60563 6670 61223 6710
rect 60563 6090 60603 6670
rect 61183 6090 61223 6670
rect 60563 6050 61223 6090
rect 67585 6670 68245 6710
rect 67585 6090 67625 6670
rect 68205 6090 68245 6670
rect 67585 6050 68245 6090
rect 69763 6670 70423 6710
rect 69763 6090 69803 6670
rect 70383 6090 70423 6670
rect 69763 6050 70423 6090
<< mimcapcontact >>
rect 3225 95010 3805 95590
rect 5403 95010 5983 95590
rect 3225 85130 3805 85710
rect 5403 85130 5983 85710
rect 12425 85130 13005 85710
rect 14603 85130 15183 85710
rect 3225 75250 3805 75830
rect 5403 75250 5983 75830
rect 12425 75250 13005 75830
rect 14603 75250 15183 75830
rect 21625 75250 22205 75830
rect 23803 75250 24383 75830
rect 30825 75250 31405 75830
rect 33003 75250 33583 75830
rect 3225 65370 3805 65950
rect 5403 65370 5983 65950
rect 12425 65370 13005 65950
rect 14603 65370 15183 65950
rect 21625 65370 22205 65950
rect 23803 65370 24383 65950
rect 30825 65370 31405 65950
rect 33003 65370 33583 65950
rect 40025 65370 40605 65950
rect 42203 65370 42783 65950
rect 49225 65370 49805 65950
rect 51403 65370 51983 65950
rect 58425 65370 59005 65950
rect 60603 65370 61183 65950
rect 67625 65370 68205 65950
rect 69803 65370 70383 65950
rect 3225 55490 3805 56070
rect 5403 55490 5983 56070
rect 12425 55490 13005 56070
rect 14603 55490 15183 56070
rect 21625 55490 22205 56070
rect 23803 55490 24383 56070
rect 30825 55490 31405 56070
rect 33003 55490 33583 56070
rect 40025 55490 40605 56070
rect 42203 55490 42783 56070
rect 49225 55490 49805 56070
rect 51403 55490 51983 56070
rect 58425 55490 59005 56070
rect 60603 55490 61183 56070
rect 67625 55490 68205 56070
rect 69803 55490 70383 56070
rect 3225 45610 3805 46190
rect 5403 45610 5983 46190
rect 12425 45610 13005 46190
rect 14603 45610 15183 46190
rect 21625 45610 22205 46190
rect 23803 45610 24383 46190
rect 30825 45610 31405 46190
rect 33003 45610 33583 46190
rect 40025 45610 40605 46190
rect 42203 45610 42783 46190
rect 49225 45610 49805 46190
rect 51403 45610 51983 46190
rect 58425 45610 59005 46190
rect 60603 45610 61183 46190
rect 67625 45610 68205 46190
rect 69803 45610 70383 46190
rect 3225 35730 3805 36310
rect 5403 35730 5983 36310
rect 12425 35730 13005 36310
rect 14603 35730 15183 36310
rect 21625 35730 22205 36310
rect 23803 35730 24383 36310
rect 30825 35730 31405 36310
rect 33003 35730 33583 36310
rect 40025 35730 40605 36310
rect 42203 35730 42783 36310
rect 49225 35730 49805 36310
rect 51403 35730 51983 36310
rect 58425 35730 59005 36310
rect 60603 35730 61183 36310
rect 67625 35730 68205 36310
rect 69803 35730 70383 36310
rect 3225 25850 3805 26430
rect 5403 25850 5983 26430
rect 12425 25850 13005 26430
rect 14603 25850 15183 26430
rect 21625 25850 22205 26430
rect 23803 25850 24383 26430
rect 30825 25850 31405 26430
rect 33003 25850 33583 26430
rect 40025 25850 40605 26430
rect 42203 25850 42783 26430
rect 49225 25850 49805 26430
rect 51403 25850 51983 26430
rect 58425 25850 59005 26430
rect 60603 25850 61183 26430
rect 67625 25850 68205 26430
rect 69803 25850 70383 26430
rect 3225 15970 3805 16550
rect 5403 15970 5983 16550
rect 12425 15970 13005 16550
rect 14603 15970 15183 16550
rect 21625 15970 22205 16550
rect 23803 15970 24383 16550
rect 30825 15970 31405 16550
rect 33003 15970 33583 16550
rect 40025 15970 40605 16550
rect 42203 15970 42783 16550
rect 49225 15970 49805 16550
rect 51403 15970 51983 16550
rect 58425 15970 59005 16550
rect 60603 15970 61183 16550
rect 67625 15970 68205 16550
rect 69803 15970 70383 16550
rect 3225 6090 3805 6670
rect 5403 6090 5983 6670
rect 12425 6090 13005 6670
rect 14603 6090 15183 6670
rect 21625 6090 22205 6670
rect 23803 6090 24383 6670
rect 30825 6090 31405 6670
rect 33003 6090 33583 6670
rect 40025 6090 40605 6670
rect 42203 6090 42783 6670
rect 49225 6090 49805 6670
rect 51403 6090 51983 6670
rect 58425 6090 59005 6670
rect 60603 6090 61183 6670
rect 67625 6090 68205 6670
rect 69803 6090 70383 6670
<< metal4 >>
rect 1000 103780 3000 110790
rect 1000 101800 1010 103780
rect 2990 101800 3000 103780
rect 1000 95350 3000 101800
rect 6210 109790 8210 110790
rect 6210 107810 6220 109790
rect 8200 107810 8210 109790
rect 3940 95702 4040 95720
rect 5170 95718 5270 95720
rect 3224 95590 3806 95591
rect 3224 95350 3225 95590
rect 1000 95250 3225 95350
rect 1000 85470 3000 95250
rect 3224 95010 3225 95250
rect 3805 95010 3806 95590
rect 3224 95009 3806 95010
rect 3940 94898 3960 95702
rect 4024 94898 4040 95702
rect 3940 94620 4040 94898
rect 5168 95702 5270 95718
rect 5168 94898 5184 95702
rect 5248 94898 5270 95702
rect 5402 95590 5984 95591
rect 5402 95010 5403 95590
rect 5983 95350 5984 95590
rect 6210 95350 8210 107810
rect 5983 95250 8210 95350
rect 5983 95010 5984 95250
rect 5402 95009 5984 95010
rect 5168 94882 5270 94898
rect 3940 94530 3950 94620
rect 4030 94530 4040 94620
rect 3940 94520 4040 94530
rect 5170 94620 5270 94882
rect 5170 94530 5180 94620
rect 5260 94530 5270 94620
rect 5170 94520 5270 94530
rect 6210 92410 8210 95250
rect 6200 88910 8210 92410
rect 3940 85822 4040 85840
rect 5170 85838 5270 85840
rect 3224 85710 3806 85711
rect 3224 85470 3225 85710
rect 1000 85370 3225 85470
rect 1000 75590 3000 85370
rect 3224 85130 3225 85370
rect 3805 85130 3806 85710
rect 3224 85129 3806 85130
rect 3940 85018 3960 85822
rect 4024 85018 4040 85822
rect 3940 84740 4040 85018
rect 5168 85822 5270 85838
rect 5168 85018 5184 85822
rect 5248 85018 5270 85822
rect 5402 85710 5984 85711
rect 5402 85130 5403 85710
rect 5983 85470 5984 85710
rect 6210 85470 8210 88910
rect 5983 85370 8210 85470
rect 5983 85130 5984 85370
rect 5402 85129 5984 85130
rect 5168 85002 5270 85018
rect 3940 84650 3950 84740
rect 4030 84650 4040 84740
rect 3940 84640 4040 84650
rect 5170 84740 5270 85002
rect 5170 84650 5180 84740
rect 5260 84650 5270 84740
rect 5170 84640 5270 84650
rect 6210 82530 8210 85370
rect 6200 79030 8210 82530
rect 3940 75942 4040 75960
rect 5170 75958 5270 75960
rect 3224 75830 3806 75831
rect 3224 75590 3225 75830
rect 1000 75490 3225 75590
rect 1000 65710 3000 75490
rect 3224 75250 3225 75490
rect 3805 75250 3806 75830
rect 3224 75249 3806 75250
rect 3940 75138 3960 75942
rect 4024 75138 4040 75942
rect 3940 74860 4040 75138
rect 5168 75942 5270 75958
rect 5168 75138 5184 75942
rect 5248 75138 5270 75942
rect 5402 75830 5984 75831
rect 5402 75250 5403 75830
rect 5983 75590 5984 75830
rect 6210 75590 8210 79030
rect 5983 75490 8210 75590
rect 5983 75250 5984 75490
rect 5402 75249 5984 75250
rect 5168 75122 5270 75138
rect 3940 74770 3950 74860
rect 4030 74770 4040 74860
rect 3940 74760 4040 74770
rect 5170 74860 5270 75122
rect 5170 74770 5180 74860
rect 5260 74770 5270 74860
rect 5170 74760 5270 74770
rect 6210 72650 8210 75490
rect 6200 69150 8210 72650
rect 3940 66062 4040 66080
rect 5170 66078 5270 66080
rect 3224 65950 3806 65951
rect 3224 65710 3225 65950
rect 1000 65610 3225 65710
rect 1000 55830 3000 65610
rect 3224 65370 3225 65610
rect 3805 65370 3806 65950
rect 3224 65369 3806 65370
rect 3940 65258 3960 66062
rect 4024 65258 4040 66062
rect 3940 64980 4040 65258
rect 5168 66062 5270 66078
rect 5168 65258 5184 66062
rect 5248 65258 5270 66062
rect 5402 65950 5984 65951
rect 5402 65370 5403 65950
rect 5983 65710 5984 65950
rect 6210 65710 8210 69150
rect 5983 65610 8210 65710
rect 5983 65370 5984 65610
rect 5402 65369 5984 65370
rect 5168 65242 5270 65258
rect 3940 64890 3950 64980
rect 4030 64890 4040 64980
rect 3940 64880 4040 64890
rect 5170 64980 5270 65242
rect 5170 64890 5180 64980
rect 5260 64890 5270 64980
rect 5170 64880 5270 64890
rect 6210 62770 8210 65610
rect 6200 59270 8210 62770
rect 3940 56182 4040 56200
rect 5170 56198 5270 56200
rect 3224 56070 3806 56071
rect 3224 55830 3225 56070
rect 1000 55730 3225 55830
rect 1000 45950 3000 55730
rect 3224 55490 3225 55730
rect 3805 55490 3806 56070
rect 3224 55489 3806 55490
rect 3940 55378 3960 56182
rect 4024 55378 4040 56182
rect 3940 55100 4040 55378
rect 5168 56182 5270 56198
rect 5168 55378 5184 56182
rect 5248 55378 5270 56182
rect 5402 56070 5984 56071
rect 5402 55490 5403 56070
rect 5983 55830 5984 56070
rect 6210 55830 8210 59270
rect 5983 55730 8210 55830
rect 5983 55490 5984 55730
rect 5402 55489 5984 55490
rect 5168 55362 5270 55378
rect 3940 55010 3950 55100
rect 4030 55010 4040 55100
rect 3940 55000 4040 55010
rect 5170 55100 5270 55362
rect 5170 55010 5180 55100
rect 5260 55010 5270 55100
rect 5170 55000 5270 55010
rect 6210 52890 8210 55730
rect 6200 49390 8210 52890
rect 3940 46302 4040 46320
rect 5170 46318 5270 46320
rect 3224 46190 3806 46191
rect 3224 45950 3225 46190
rect 1000 45850 3225 45950
rect 1000 36070 3000 45850
rect 3224 45610 3225 45850
rect 3805 45610 3806 46190
rect 3224 45609 3806 45610
rect 3940 45498 3960 46302
rect 4024 45498 4040 46302
rect 3940 45220 4040 45498
rect 5168 46302 5270 46318
rect 5168 45498 5184 46302
rect 5248 45498 5270 46302
rect 5402 46190 5984 46191
rect 5402 45610 5403 46190
rect 5983 45950 5984 46190
rect 6210 45950 8210 49390
rect 5983 45850 8210 45950
rect 5983 45610 5984 45850
rect 5402 45609 5984 45610
rect 5168 45482 5270 45498
rect 3940 45130 3950 45220
rect 4030 45130 4040 45220
rect 3940 45120 4040 45130
rect 5170 45220 5270 45482
rect 5170 45130 5180 45220
rect 5260 45130 5270 45220
rect 5170 45120 5270 45130
rect 6210 43010 8210 45850
rect 6200 39510 8210 43010
rect 3940 36422 4040 36440
rect 5170 36438 5270 36440
rect 3224 36310 3806 36311
rect 3224 36070 3225 36310
rect 1000 35970 3225 36070
rect 1000 26190 3000 35970
rect 3224 35730 3225 35970
rect 3805 35730 3806 36310
rect 3224 35729 3806 35730
rect 3940 35618 3960 36422
rect 4024 35618 4040 36422
rect 3940 35340 4040 35618
rect 5168 36422 5270 36438
rect 5168 35618 5184 36422
rect 5248 35618 5270 36422
rect 5402 36310 5984 36311
rect 5402 35730 5403 36310
rect 5983 36070 5984 36310
rect 6210 36070 8210 39510
rect 5983 35970 8210 36070
rect 5983 35730 5984 35970
rect 5402 35729 5984 35730
rect 5168 35602 5270 35618
rect 3940 35250 3950 35340
rect 4030 35250 4040 35340
rect 3940 35240 4040 35250
rect 5170 35340 5270 35602
rect 5170 35250 5180 35340
rect 5260 35250 5270 35340
rect 5170 35240 5270 35250
rect 6210 33130 8210 35970
rect 6200 29630 8210 33130
rect 3940 26542 4040 26560
rect 5170 26558 5270 26560
rect 3224 26430 3806 26431
rect 3224 26190 3225 26430
rect 1000 26090 3225 26190
rect 1000 16310 3000 26090
rect 3224 25850 3225 26090
rect 3805 25850 3806 26430
rect 3224 25849 3806 25850
rect 3940 25738 3960 26542
rect 4024 25738 4040 26542
rect 3940 25460 4040 25738
rect 5168 26542 5270 26558
rect 5168 25738 5184 26542
rect 5248 25738 5270 26542
rect 5402 26430 5984 26431
rect 5402 25850 5403 26430
rect 5983 26190 5984 26430
rect 6210 26190 8210 29630
rect 5983 26090 8210 26190
rect 5983 25850 5984 26090
rect 5402 25849 5984 25850
rect 5168 25722 5270 25738
rect 3940 25370 3950 25460
rect 4030 25370 4040 25460
rect 3940 25360 4040 25370
rect 5170 25460 5270 25722
rect 5170 25370 5180 25460
rect 5260 25370 5270 25460
rect 5170 25360 5270 25370
rect 6210 23250 8210 26090
rect 6200 19750 8210 23250
rect 3940 16662 4040 16680
rect 5170 16678 5270 16680
rect 3224 16550 3806 16551
rect 3224 16310 3225 16550
rect 1000 16210 3225 16310
rect 1000 6430 3000 16210
rect 3224 15970 3225 16210
rect 3805 15970 3806 16550
rect 3224 15969 3806 15970
rect 3940 15858 3960 16662
rect 4024 15858 4040 16662
rect 3940 15580 4040 15858
rect 5168 16662 5270 16678
rect 5168 15858 5184 16662
rect 5248 15858 5270 16662
rect 5402 16550 5984 16551
rect 5402 15970 5403 16550
rect 5983 16310 5984 16550
rect 6210 16310 8210 19750
rect 5983 16210 8210 16310
rect 5983 15970 5984 16210
rect 5402 15969 5984 15970
rect 5168 15842 5270 15858
rect 3940 15490 3950 15580
rect 4030 15490 4040 15580
rect 3940 15480 4040 15490
rect 5170 15580 5270 15842
rect 5170 15490 5180 15580
rect 5260 15490 5270 15580
rect 5170 15480 5270 15490
rect 6210 13370 8210 16210
rect 6200 9870 8210 13370
rect 3940 6782 4040 6800
rect 5170 6798 5270 6800
rect 3224 6670 3806 6671
rect 3224 6430 3225 6670
rect 1000 6330 3225 6430
rect 1000 -10 3000 6330
rect 3224 6090 3225 6330
rect 3805 6090 3806 6670
rect 3224 6089 3806 6090
rect 3940 5978 3960 6782
rect 4024 5978 4040 6782
rect 3940 5700 4040 5978
rect 5168 6782 5270 6798
rect 5168 5978 5184 6782
rect 5248 5978 5270 6782
rect 5402 6670 5984 6671
rect 5402 6090 5403 6670
rect 5983 6430 5984 6670
rect 6210 6430 8210 9870
rect 5983 6330 8210 6430
rect 5983 6090 5984 6330
rect 5402 6089 5984 6090
rect 5168 5962 5270 5978
rect 3940 5610 3950 5700
rect 4030 5610 4040 5700
rect 3940 5600 4040 5610
rect 5170 5700 5270 5962
rect 5170 5610 5180 5700
rect 5260 5610 5270 5700
rect 5170 5600 5270 5610
rect 6210 3490 8210 6330
rect 6200 -10 8210 3490
rect 10200 103780 12200 110790
rect 10200 101800 10210 103780
rect 12190 101800 12200 103780
rect 10200 85470 12200 101800
rect 15410 109790 17410 110790
rect 15410 107810 15420 109790
rect 17400 107810 17410 109790
rect 13140 85822 13240 85840
rect 14370 85838 14470 85840
rect 12424 85710 13006 85711
rect 12424 85470 12425 85710
rect 10200 85370 12425 85470
rect 10200 75590 12200 85370
rect 12424 85130 12425 85370
rect 13005 85130 13006 85710
rect 12424 85129 13006 85130
rect 13140 85018 13160 85822
rect 13224 85018 13240 85822
rect 13140 84740 13240 85018
rect 14368 85822 14470 85838
rect 14368 85018 14384 85822
rect 14448 85018 14470 85822
rect 14602 85710 15184 85711
rect 14602 85130 14603 85710
rect 15183 85470 15184 85710
rect 15410 85470 17410 107810
rect 15183 85370 17410 85470
rect 15183 85130 15184 85370
rect 14602 85129 15184 85130
rect 14368 85002 14470 85018
rect 13140 84650 13150 84740
rect 13230 84650 13240 84740
rect 13140 84640 13240 84650
rect 14370 84740 14470 85002
rect 14370 84650 14380 84740
rect 14460 84650 14470 84740
rect 14370 84640 14470 84650
rect 15410 82530 17410 85370
rect 15400 79030 17410 82530
rect 13140 75942 13240 75960
rect 14370 75958 14470 75960
rect 12424 75830 13006 75831
rect 12424 75590 12425 75830
rect 10200 75490 12425 75590
rect 10200 65710 12200 75490
rect 12424 75250 12425 75490
rect 13005 75250 13006 75830
rect 12424 75249 13006 75250
rect 13140 75138 13160 75942
rect 13224 75138 13240 75942
rect 13140 74860 13240 75138
rect 14368 75942 14470 75958
rect 14368 75138 14384 75942
rect 14448 75138 14470 75942
rect 14602 75830 15184 75831
rect 14602 75250 14603 75830
rect 15183 75590 15184 75830
rect 15410 75590 17410 79030
rect 15183 75490 17410 75590
rect 15183 75250 15184 75490
rect 14602 75249 15184 75250
rect 14368 75122 14470 75138
rect 13140 74770 13150 74860
rect 13230 74770 13240 74860
rect 13140 74760 13240 74770
rect 14370 74860 14470 75122
rect 14370 74770 14380 74860
rect 14460 74770 14470 74860
rect 14370 74760 14470 74770
rect 15410 72650 17410 75490
rect 15400 69150 17410 72650
rect 13140 66062 13240 66080
rect 14370 66078 14470 66080
rect 12424 65950 13006 65951
rect 12424 65710 12425 65950
rect 10200 65610 12425 65710
rect 10200 55830 12200 65610
rect 12424 65370 12425 65610
rect 13005 65370 13006 65950
rect 12424 65369 13006 65370
rect 13140 65258 13160 66062
rect 13224 65258 13240 66062
rect 13140 64980 13240 65258
rect 14368 66062 14470 66078
rect 14368 65258 14384 66062
rect 14448 65258 14470 66062
rect 14602 65950 15184 65951
rect 14602 65370 14603 65950
rect 15183 65710 15184 65950
rect 15410 65710 17410 69150
rect 15183 65610 17410 65710
rect 15183 65370 15184 65610
rect 14602 65369 15184 65370
rect 14368 65242 14470 65258
rect 13140 64890 13150 64980
rect 13230 64890 13240 64980
rect 13140 64880 13240 64890
rect 14370 64980 14470 65242
rect 14370 64890 14380 64980
rect 14460 64890 14470 64980
rect 14370 64880 14470 64890
rect 15410 62770 17410 65610
rect 15400 59270 17410 62770
rect 13140 56182 13240 56200
rect 14370 56198 14470 56200
rect 12424 56070 13006 56071
rect 12424 55830 12425 56070
rect 10200 55730 12425 55830
rect 10200 45950 12200 55730
rect 12424 55490 12425 55730
rect 13005 55490 13006 56070
rect 12424 55489 13006 55490
rect 13140 55378 13160 56182
rect 13224 55378 13240 56182
rect 13140 55100 13240 55378
rect 14368 56182 14470 56198
rect 14368 55378 14384 56182
rect 14448 55378 14470 56182
rect 14602 56070 15184 56071
rect 14602 55490 14603 56070
rect 15183 55830 15184 56070
rect 15410 55830 17410 59270
rect 15183 55730 17410 55830
rect 15183 55490 15184 55730
rect 14602 55489 15184 55490
rect 14368 55362 14470 55378
rect 13140 55010 13150 55100
rect 13230 55010 13240 55100
rect 13140 55000 13240 55010
rect 14370 55100 14470 55362
rect 14370 55010 14380 55100
rect 14460 55010 14470 55100
rect 14370 55000 14470 55010
rect 15410 52890 17410 55730
rect 15400 49390 17410 52890
rect 13140 46302 13240 46320
rect 14370 46318 14470 46320
rect 12424 46190 13006 46191
rect 12424 45950 12425 46190
rect 10200 45850 12425 45950
rect 10200 36070 12200 45850
rect 12424 45610 12425 45850
rect 13005 45610 13006 46190
rect 12424 45609 13006 45610
rect 13140 45498 13160 46302
rect 13224 45498 13240 46302
rect 13140 45220 13240 45498
rect 14368 46302 14470 46318
rect 14368 45498 14384 46302
rect 14448 45498 14470 46302
rect 14602 46190 15184 46191
rect 14602 45610 14603 46190
rect 15183 45950 15184 46190
rect 15410 45950 17410 49390
rect 15183 45850 17410 45950
rect 15183 45610 15184 45850
rect 14602 45609 15184 45610
rect 14368 45482 14470 45498
rect 13140 45130 13150 45220
rect 13230 45130 13240 45220
rect 13140 45120 13240 45130
rect 14370 45220 14470 45482
rect 14370 45130 14380 45220
rect 14460 45130 14470 45220
rect 14370 45120 14470 45130
rect 15410 43010 17410 45850
rect 15400 39510 17410 43010
rect 13140 36422 13240 36440
rect 14370 36438 14470 36440
rect 12424 36310 13006 36311
rect 12424 36070 12425 36310
rect 10200 35970 12425 36070
rect 10200 26190 12200 35970
rect 12424 35730 12425 35970
rect 13005 35730 13006 36310
rect 12424 35729 13006 35730
rect 13140 35618 13160 36422
rect 13224 35618 13240 36422
rect 13140 35340 13240 35618
rect 14368 36422 14470 36438
rect 14368 35618 14384 36422
rect 14448 35618 14470 36422
rect 14602 36310 15184 36311
rect 14602 35730 14603 36310
rect 15183 36070 15184 36310
rect 15410 36070 17410 39510
rect 15183 35970 17410 36070
rect 15183 35730 15184 35970
rect 14602 35729 15184 35730
rect 14368 35602 14470 35618
rect 13140 35250 13150 35340
rect 13230 35250 13240 35340
rect 13140 35240 13240 35250
rect 14370 35340 14470 35602
rect 14370 35250 14380 35340
rect 14460 35250 14470 35340
rect 14370 35240 14470 35250
rect 15410 33130 17410 35970
rect 15400 29630 17410 33130
rect 13140 26542 13240 26560
rect 14370 26558 14470 26560
rect 12424 26430 13006 26431
rect 12424 26190 12425 26430
rect 10200 26090 12425 26190
rect 10200 16310 12200 26090
rect 12424 25850 12425 26090
rect 13005 25850 13006 26430
rect 12424 25849 13006 25850
rect 13140 25738 13160 26542
rect 13224 25738 13240 26542
rect 13140 25460 13240 25738
rect 14368 26542 14470 26558
rect 14368 25738 14384 26542
rect 14448 25738 14470 26542
rect 14602 26430 15184 26431
rect 14602 25850 14603 26430
rect 15183 26190 15184 26430
rect 15410 26190 17410 29630
rect 15183 26090 17410 26190
rect 15183 25850 15184 26090
rect 14602 25849 15184 25850
rect 14368 25722 14470 25738
rect 13140 25370 13150 25460
rect 13230 25370 13240 25460
rect 13140 25360 13240 25370
rect 14370 25460 14470 25722
rect 14370 25370 14380 25460
rect 14460 25370 14470 25460
rect 14370 25360 14470 25370
rect 15410 23250 17410 26090
rect 15400 19750 17410 23250
rect 13140 16662 13240 16680
rect 14370 16678 14470 16680
rect 12424 16550 13006 16551
rect 12424 16310 12425 16550
rect 10200 16210 12425 16310
rect 10200 6430 12200 16210
rect 12424 15970 12425 16210
rect 13005 15970 13006 16550
rect 12424 15969 13006 15970
rect 13140 15858 13160 16662
rect 13224 15858 13240 16662
rect 13140 15580 13240 15858
rect 14368 16662 14470 16678
rect 14368 15858 14384 16662
rect 14448 15858 14470 16662
rect 14602 16550 15184 16551
rect 14602 15970 14603 16550
rect 15183 16310 15184 16550
rect 15410 16310 17410 19750
rect 15183 16210 17410 16310
rect 15183 15970 15184 16210
rect 14602 15969 15184 15970
rect 14368 15842 14470 15858
rect 13140 15490 13150 15580
rect 13230 15490 13240 15580
rect 13140 15480 13240 15490
rect 14370 15580 14470 15842
rect 14370 15490 14380 15580
rect 14460 15490 14470 15580
rect 14370 15480 14470 15490
rect 15410 13370 17410 16210
rect 15400 9870 17410 13370
rect 13140 6782 13240 6800
rect 14370 6798 14470 6800
rect 12424 6670 13006 6671
rect 12424 6430 12425 6670
rect 10200 6330 12425 6430
rect 10200 -10 12200 6330
rect 12424 6090 12425 6330
rect 13005 6090 13006 6670
rect 12424 6089 13006 6090
rect 13140 5978 13160 6782
rect 13224 5978 13240 6782
rect 13140 5700 13240 5978
rect 14368 6782 14470 6798
rect 14368 5978 14384 6782
rect 14448 5978 14470 6782
rect 14602 6670 15184 6671
rect 14602 6090 14603 6670
rect 15183 6430 15184 6670
rect 15410 6430 17410 9870
rect 15183 6330 17410 6430
rect 15183 6090 15184 6330
rect 14602 6089 15184 6090
rect 14368 5962 14470 5978
rect 13140 5610 13150 5700
rect 13230 5610 13240 5700
rect 13140 5600 13240 5610
rect 14370 5700 14470 5962
rect 14370 5610 14380 5700
rect 14460 5610 14470 5700
rect 14370 5600 14470 5610
rect 15410 3490 17410 6330
rect 15400 -10 17410 3490
rect 19400 103780 21400 110790
rect 19400 101800 19410 103780
rect 21390 101800 21400 103780
rect 19400 75590 21400 101800
rect 24610 109790 26610 110790
rect 24610 107810 24620 109790
rect 26600 107810 26610 109790
rect 22340 75942 22440 75960
rect 23570 75958 23670 75960
rect 21624 75830 22206 75831
rect 21624 75590 21625 75830
rect 19400 75490 21625 75590
rect 19400 65710 21400 75490
rect 21624 75250 21625 75490
rect 22205 75250 22206 75830
rect 21624 75249 22206 75250
rect 22340 75138 22360 75942
rect 22424 75138 22440 75942
rect 22340 74860 22440 75138
rect 23568 75942 23670 75958
rect 23568 75138 23584 75942
rect 23648 75138 23670 75942
rect 23802 75830 24384 75831
rect 23802 75250 23803 75830
rect 24383 75590 24384 75830
rect 24610 75590 26610 107810
rect 24383 75490 26610 75590
rect 24383 75250 24384 75490
rect 23802 75249 24384 75250
rect 23568 75122 23670 75138
rect 22340 74770 22350 74860
rect 22430 74770 22440 74860
rect 22340 74760 22440 74770
rect 23570 74860 23670 75122
rect 23570 74770 23580 74860
rect 23660 74770 23670 74860
rect 23570 74760 23670 74770
rect 24610 72650 26610 75490
rect 24600 69150 26610 72650
rect 22340 66062 22440 66080
rect 23570 66078 23670 66080
rect 21624 65950 22206 65951
rect 21624 65710 21625 65950
rect 19400 65610 21625 65710
rect 19400 55830 21400 65610
rect 21624 65370 21625 65610
rect 22205 65370 22206 65950
rect 21624 65369 22206 65370
rect 22340 65258 22360 66062
rect 22424 65258 22440 66062
rect 22340 64980 22440 65258
rect 23568 66062 23670 66078
rect 23568 65258 23584 66062
rect 23648 65258 23670 66062
rect 23802 65950 24384 65951
rect 23802 65370 23803 65950
rect 24383 65710 24384 65950
rect 24610 65710 26610 69150
rect 24383 65610 26610 65710
rect 24383 65370 24384 65610
rect 23802 65369 24384 65370
rect 23568 65242 23670 65258
rect 22340 64890 22350 64980
rect 22430 64890 22440 64980
rect 22340 64880 22440 64890
rect 23570 64980 23670 65242
rect 23570 64890 23580 64980
rect 23660 64890 23670 64980
rect 23570 64880 23670 64890
rect 24610 62770 26610 65610
rect 24600 59270 26610 62770
rect 22340 56182 22440 56200
rect 23570 56198 23670 56200
rect 21624 56070 22206 56071
rect 21624 55830 21625 56070
rect 19400 55730 21625 55830
rect 19400 45950 21400 55730
rect 21624 55490 21625 55730
rect 22205 55490 22206 56070
rect 21624 55489 22206 55490
rect 22340 55378 22360 56182
rect 22424 55378 22440 56182
rect 22340 55100 22440 55378
rect 23568 56182 23670 56198
rect 23568 55378 23584 56182
rect 23648 55378 23670 56182
rect 23802 56070 24384 56071
rect 23802 55490 23803 56070
rect 24383 55830 24384 56070
rect 24610 55830 26610 59270
rect 24383 55730 26610 55830
rect 24383 55490 24384 55730
rect 23802 55489 24384 55490
rect 23568 55362 23670 55378
rect 22340 55010 22350 55100
rect 22430 55010 22440 55100
rect 22340 55000 22440 55010
rect 23570 55100 23670 55362
rect 23570 55010 23580 55100
rect 23660 55010 23670 55100
rect 23570 55000 23670 55010
rect 24610 52890 26610 55730
rect 24600 49390 26610 52890
rect 22340 46302 22440 46320
rect 23570 46318 23670 46320
rect 21624 46190 22206 46191
rect 21624 45950 21625 46190
rect 19400 45850 21625 45950
rect 19400 36070 21400 45850
rect 21624 45610 21625 45850
rect 22205 45610 22206 46190
rect 21624 45609 22206 45610
rect 22340 45498 22360 46302
rect 22424 45498 22440 46302
rect 22340 45220 22440 45498
rect 23568 46302 23670 46318
rect 23568 45498 23584 46302
rect 23648 45498 23670 46302
rect 23802 46190 24384 46191
rect 23802 45610 23803 46190
rect 24383 45950 24384 46190
rect 24610 45950 26610 49390
rect 24383 45850 26610 45950
rect 24383 45610 24384 45850
rect 23802 45609 24384 45610
rect 23568 45482 23670 45498
rect 22340 45130 22350 45220
rect 22430 45130 22440 45220
rect 22340 45120 22440 45130
rect 23570 45220 23670 45482
rect 23570 45130 23580 45220
rect 23660 45130 23670 45220
rect 23570 45120 23670 45130
rect 24610 43010 26610 45850
rect 24600 39510 26610 43010
rect 22340 36422 22440 36440
rect 23570 36438 23670 36440
rect 21624 36310 22206 36311
rect 21624 36070 21625 36310
rect 19400 35970 21625 36070
rect 19400 26190 21400 35970
rect 21624 35730 21625 35970
rect 22205 35730 22206 36310
rect 21624 35729 22206 35730
rect 22340 35618 22360 36422
rect 22424 35618 22440 36422
rect 22340 35340 22440 35618
rect 23568 36422 23670 36438
rect 23568 35618 23584 36422
rect 23648 35618 23670 36422
rect 23802 36310 24384 36311
rect 23802 35730 23803 36310
rect 24383 36070 24384 36310
rect 24610 36070 26610 39510
rect 24383 35970 26610 36070
rect 24383 35730 24384 35970
rect 23802 35729 24384 35730
rect 23568 35602 23670 35618
rect 22340 35250 22350 35340
rect 22430 35250 22440 35340
rect 22340 35240 22440 35250
rect 23570 35340 23670 35602
rect 23570 35250 23580 35340
rect 23660 35250 23670 35340
rect 23570 35240 23670 35250
rect 24610 33130 26610 35970
rect 24600 29630 26610 33130
rect 22340 26542 22440 26560
rect 23570 26558 23670 26560
rect 21624 26430 22206 26431
rect 21624 26190 21625 26430
rect 19400 26090 21625 26190
rect 19400 16310 21400 26090
rect 21624 25850 21625 26090
rect 22205 25850 22206 26430
rect 21624 25849 22206 25850
rect 22340 25738 22360 26542
rect 22424 25738 22440 26542
rect 22340 25460 22440 25738
rect 23568 26542 23670 26558
rect 23568 25738 23584 26542
rect 23648 25738 23670 26542
rect 23802 26430 24384 26431
rect 23802 25850 23803 26430
rect 24383 26190 24384 26430
rect 24610 26190 26610 29630
rect 24383 26090 26610 26190
rect 24383 25850 24384 26090
rect 23802 25849 24384 25850
rect 23568 25722 23670 25738
rect 22340 25370 22350 25460
rect 22430 25370 22440 25460
rect 22340 25360 22440 25370
rect 23570 25460 23670 25722
rect 23570 25370 23580 25460
rect 23660 25370 23670 25460
rect 23570 25360 23670 25370
rect 24610 23250 26610 26090
rect 24600 19750 26610 23250
rect 22340 16662 22440 16680
rect 23570 16678 23670 16680
rect 21624 16550 22206 16551
rect 21624 16310 21625 16550
rect 19400 16210 21625 16310
rect 19400 6430 21400 16210
rect 21624 15970 21625 16210
rect 22205 15970 22206 16550
rect 21624 15969 22206 15970
rect 22340 15858 22360 16662
rect 22424 15858 22440 16662
rect 22340 15580 22440 15858
rect 23568 16662 23670 16678
rect 23568 15858 23584 16662
rect 23648 15858 23670 16662
rect 23802 16550 24384 16551
rect 23802 15970 23803 16550
rect 24383 16310 24384 16550
rect 24610 16310 26610 19750
rect 24383 16210 26610 16310
rect 24383 15970 24384 16210
rect 23802 15969 24384 15970
rect 23568 15842 23670 15858
rect 22340 15490 22350 15580
rect 22430 15490 22440 15580
rect 22340 15480 22440 15490
rect 23570 15580 23670 15842
rect 23570 15490 23580 15580
rect 23660 15490 23670 15580
rect 23570 15480 23670 15490
rect 24610 13370 26610 16210
rect 24600 9870 26610 13370
rect 22340 6782 22440 6800
rect 23570 6798 23670 6800
rect 21624 6670 22206 6671
rect 21624 6430 21625 6670
rect 19400 6330 21625 6430
rect 19400 -10 21400 6330
rect 21624 6090 21625 6330
rect 22205 6090 22206 6670
rect 21624 6089 22206 6090
rect 22340 5978 22360 6782
rect 22424 5978 22440 6782
rect 22340 5700 22440 5978
rect 23568 6782 23670 6798
rect 23568 5978 23584 6782
rect 23648 5978 23670 6782
rect 23802 6670 24384 6671
rect 23802 6090 23803 6670
rect 24383 6430 24384 6670
rect 24610 6430 26610 9870
rect 24383 6330 26610 6430
rect 24383 6090 24384 6330
rect 23802 6089 24384 6090
rect 23568 5962 23670 5978
rect 22340 5610 22350 5700
rect 22430 5610 22440 5700
rect 22340 5600 22440 5610
rect 23570 5700 23670 5962
rect 23570 5610 23580 5700
rect 23660 5610 23670 5700
rect 23570 5600 23670 5610
rect 24610 3490 26610 6330
rect 24600 -10 26610 3490
rect 28600 103780 30600 110790
rect 28600 101800 28610 103780
rect 30590 101800 30600 103780
rect 28600 75590 30600 101800
rect 33810 109790 35810 110790
rect 33810 107810 33820 109790
rect 35800 107810 35810 109790
rect 31540 75942 31640 75960
rect 32770 75958 32870 75960
rect 30824 75830 31406 75831
rect 30824 75590 30825 75830
rect 28600 75490 30825 75590
rect 28600 65710 30600 75490
rect 30824 75250 30825 75490
rect 31405 75250 31406 75830
rect 30824 75249 31406 75250
rect 31540 75138 31560 75942
rect 31624 75138 31640 75942
rect 31540 74860 31640 75138
rect 32768 75942 32870 75958
rect 32768 75138 32784 75942
rect 32848 75138 32870 75942
rect 33002 75830 33584 75831
rect 33002 75250 33003 75830
rect 33583 75590 33584 75830
rect 33810 75590 35810 107810
rect 33583 75490 35810 75590
rect 33583 75250 33584 75490
rect 33002 75249 33584 75250
rect 32768 75122 32870 75138
rect 31540 74770 31550 74860
rect 31630 74770 31640 74860
rect 31540 74760 31640 74770
rect 32770 74860 32870 75122
rect 32770 74770 32780 74860
rect 32860 74770 32870 74860
rect 32770 74760 32870 74770
rect 33810 72650 35810 75490
rect 33800 69150 35810 72650
rect 31540 66062 31640 66080
rect 32770 66078 32870 66080
rect 30824 65950 31406 65951
rect 30824 65710 30825 65950
rect 28600 65610 30825 65710
rect 28600 55830 30600 65610
rect 30824 65370 30825 65610
rect 31405 65370 31406 65950
rect 30824 65369 31406 65370
rect 31540 65258 31560 66062
rect 31624 65258 31640 66062
rect 31540 64980 31640 65258
rect 32768 66062 32870 66078
rect 32768 65258 32784 66062
rect 32848 65258 32870 66062
rect 33002 65950 33584 65951
rect 33002 65370 33003 65950
rect 33583 65710 33584 65950
rect 33810 65710 35810 69150
rect 33583 65610 35810 65710
rect 33583 65370 33584 65610
rect 33002 65369 33584 65370
rect 32768 65242 32870 65258
rect 31540 64890 31550 64980
rect 31630 64890 31640 64980
rect 31540 64880 31640 64890
rect 32770 64980 32870 65242
rect 32770 64890 32780 64980
rect 32860 64890 32870 64980
rect 32770 64880 32870 64890
rect 33810 62770 35810 65610
rect 33800 59270 35810 62770
rect 31540 56182 31640 56200
rect 32770 56198 32870 56200
rect 30824 56070 31406 56071
rect 30824 55830 30825 56070
rect 28600 55730 30825 55830
rect 28600 45950 30600 55730
rect 30824 55490 30825 55730
rect 31405 55490 31406 56070
rect 30824 55489 31406 55490
rect 31540 55378 31560 56182
rect 31624 55378 31640 56182
rect 31540 55100 31640 55378
rect 32768 56182 32870 56198
rect 32768 55378 32784 56182
rect 32848 55378 32870 56182
rect 33002 56070 33584 56071
rect 33002 55490 33003 56070
rect 33583 55830 33584 56070
rect 33810 55830 35810 59270
rect 33583 55730 35810 55830
rect 33583 55490 33584 55730
rect 33002 55489 33584 55490
rect 32768 55362 32870 55378
rect 31540 55010 31550 55100
rect 31630 55010 31640 55100
rect 31540 55000 31640 55010
rect 32770 55100 32870 55362
rect 32770 55010 32780 55100
rect 32860 55010 32870 55100
rect 32770 55000 32870 55010
rect 33810 52890 35810 55730
rect 33800 49390 35810 52890
rect 31540 46302 31640 46320
rect 32770 46318 32870 46320
rect 30824 46190 31406 46191
rect 30824 45950 30825 46190
rect 28600 45850 30825 45950
rect 28600 36070 30600 45850
rect 30824 45610 30825 45850
rect 31405 45610 31406 46190
rect 30824 45609 31406 45610
rect 31540 45498 31560 46302
rect 31624 45498 31640 46302
rect 31540 45220 31640 45498
rect 32768 46302 32870 46318
rect 32768 45498 32784 46302
rect 32848 45498 32870 46302
rect 33002 46190 33584 46191
rect 33002 45610 33003 46190
rect 33583 45950 33584 46190
rect 33810 45950 35810 49390
rect 33583 45850 35810 45950
rect 33583 45610 33584 45850
rect 33002 45609 33584 45610
rect 32768 45482 32870 45498
rect 31540 45130 31550 45220
rect 31630 45130 31640 45220
rect 31540 45120 31640 45130
rect 32770 45220 32870 45482
rect 32770 45130 32780 45220
rect 32860 45130 32870 45220
rect 32770 45120 32870 45130
rect 33810 43010 35810 45850
rect 33800 39510 35810 43010
rect 31540 36422 31640 36440
rect 32770 36438 32870 36440
rect 30824 36310 31406 36311
rect 30824 36070 30825 36310
rect 28600 35970 30825 36070
rect 28600 26190 30600 35970
rect 30824 35730 30825 35970
rect 31405 35730 31406 36310
rect 30824 35729 31406 35730
rect 31540 35618 31560 36422
rect 31624 35618 31640 36422
rect 31540 35340 31640 35618
rect 32768 36422 32870 36438
rect 32768 35618 32784 36422
rect 32848 35618 32870 36422
rect 33002 36310 33584 36311
rect 33002 35730 33003 36310
rect 33583 36070 33584 36310
rect 33810 36070 35810 39510
rect 33583 35970 35810 36070
rect 33583 35730 33584 35970
rect 33002 35729 33584 35730
rect 32768 35602 32870 35618
rect 31540 35250 31550 35340
rect 31630 35250 31640 35340
rect 31540 35240 31640 35250
rect 32770 35340 32870 35602
rect 32770 35250 32780 35340
rect 32860 35250 32870 35340
rect 32770 35240 32870 35250
rect 33810 33130 35810 35970
rect 33800 29630 35810 33130
rect 31540 26542 31640 26560
rect 32770 26558 32870 26560
rect 30824 26430 31406 26431
rect 30824 26190 30825 26430
rect 28600 26090 30825 26190
rect 28600 16310 30600 26090
rect 30824 25850 30825 26090
rect 31405 25850 31406 26430
rect 30824 25849 31406 25850
rect 31540 25738 31560 26542
rect 31624 25738 31640 26542
rect 31540 25460 31640 25738
rect 32768 26542 32870 26558
rect 32768 25738 32784 26542
rect 32848 25738 32870 26542
rect 33002 26430 33584 26431
rect 33002 25850 33003 26430
rect 33583 26190 33584 26430
rect 33810 26190 35810 29630
rect 33583 26090 35810 26190
rect 33583 25850 33584 26090
rect 33002 25849 33584 25850
rect 32768 25722 32870 25738
rect 31540 25370 31550 25460
rect 31630 25370 31640 25460
rect 31540 25360 31640 25370
rect 32770 25460 32870 25722
rect 32770 25370 32780 25460
rect 32860 25370 32870 25460
rect 32770 25360 32870 25370
rect 33810 23250 35810 26090
rect 33800 19750 35810 23250
rect 31540 16662 31640 16680
rect 32770 16678 32870 16680
rect 30824 16550 31406 16551
rect 30824 16310 30825 16550
rect 28600 16210 30825 16310
rect 28600 6430 30600 16210
rect 30824 15970 30825 16210
rect 31405 15970 31406 16550
rect 30824 15969 31406 15970
rect 31540 15858 31560 16662
rect 31624 15858 31640 16662
rect 31540 15580 31640 15858
rect 32768 16662 32870 16678
rect 32768 15858 32784 16662
rect 32848 15858 32870 16662
rect 33002 16550 33584 16551
rect 33002 15970 33003 16550
rect 33583 16310 33584 16550
rect 33810 16310 35810 19750
rect 33583 16210 35810 16310
rect 33583 15970 33584 16210
rect 33002 15969 33584 15970
rect 32768 15842 32870 15858
rect 31540 15490 31550 15580
rect 31630 15490 31640 15580
rect 31540 15480 31640 15490
rect 32770 15580 32870 15842
rect 32770 15490 32780 15580
rect 32860 15490 32870 15580
rect 32770 15480 32870 15490
rect 33810 13370 35810 16210
rect 33800 9870 35810 13370
rect 31540 6782 31640 6800
rect 32770 6798 32870 6800
rect 30824 6670 31406 6671
rect 30824 6430 30825 6670
rect 28600 6330 30825 6430
rect 28600 -10 30600 6330
rect 30824 6090 30825 6330
rect 31405 6090 31406 6670
rect 30824 6089 31406 6090
rect 31540 5978 31560 6782
rect 31624 5978 31640 6782
rect 31540 5700 31640 5978
rect 32768 6782 32870 6798
rect 32768 5978 32784 6782
rect 32848 5978 32870 6782
rect 33002 6670 33584 6671
rect 33002 6090 33003 6670
rect 33583 6430 33584 6670
rect 33810 6430 35810 9870
rect 33583 6330 35810 6430
rect 33583 6090 33584 6330
rect 33002 6089 33584 6090
rect 32768 5962 32870 5978
rect 31540 5610 31550 5700
rect 31630 5610 31640 5700
rect 31540 5600 31640 5610
rect 32770 5700 32870 5962
rect 32770 5610 32780 5700
rect 32860 5610 32870 5700
rect 32770 5600 32870 5610
rect 33810 3490 35810 6330
rect 33800 -10 35810 3490
rect 37800 103780 39800 110790
rect 37800 101800 37810 103780
rect 39790 101800 39800 103780
rect 37800 65710 39800 101800
rect 43010 109790 45010 110790
rect 43010 107810 43020 109790
rect 45000 107810 45010 109790
rect 40740 66062 40840 66080
rect 41970 66078 42070 66080
rect 40024 65950 40606 65951
rect 40024 65710 40025 65950
rect 37800 65610 40025 65710
rect 37800 55830 39800 65610
rect 40024 65370 40025 65610
rect 40605 65370 40606 65950
rect 40024 65369 40606 65370
rect 40740 65258 40760 66062
rect 40824 65258 40840 66062
rect 40740 64980 40840 65258
rect 41968 66062 42070 66078
rect 41968 65258 41984 66062
rect 42048 65258 42070 66062
rect 42202 65950 42784 65951
rect 42202 65370 42203 65950
rect 42783 65710 42784 65950
rect 43010 65710 45010 107810
rect 42783 65610 45010 65710
rect 42783 65370 42784 65610
rect 42202 65369 42784 65370
rect 41968 65242 42070 65258
rect 40740 64890 40750 64980
rect 40830 64890 40840 64980
rect 40740 64880 40840 64890
rect 41970 64980 42070 65242
rect 41970 64890 41980 64980
rect 42060 64890 42070 64980
rect 41970 64880 42070 64890
rect 43010 62770 45010 65610
rect 43000 59270 45010 62770
rect 40740 56182 40840 56200
rect 41970 56198 42070 56200
rect 40024 56070 40606 56071
rect 40024 55830 40025 56070
rect 37800 55730 40025 55830
rect 37800 45950 39800 55730
rect 40024 55490 40025 55730
rect 40605 55490 40606 56070
rect 40024 55489 40606 55490
rect 40740 55378 40760 56182
rect 40824 55378 40840 56182
rect 40740 55100 40840 55378
rect 41968 56182 42070 56198
rect 41968 55378 41984 56182
rect 42048 55378 42070 56182
rect 42202 56070 42784 56071
rect 42202 55490 42203 56070
rect 42783 55830 42784 56070
rect 43010 55830 45010 59270
rect 42783 55730 45010 55830
rect 42783 55490 42784 55730
rect 42202 55489 42784 55490
rect 41968 55362 42070 55378
rect 40740 55010 40750 55100
rect 40830 55010 40840 55100
rect 40740 55000 40840 55010
rect 41970 55100 42070 55362
rect 41970 55010 41980 55100
rect 42060 55010 42070 55100
rect 41970 55000 42070 55010
rect 43010 52890 45010 55730
rect 43000 49390 45010 52890
rect 40740 46302 40840 46320
rect 41970 46318 42070 46320
rect 40024 46190 40606 46191
rect 40024 45950 40025 46190
rect 37800 45850 40025 45950
rect 37800 36070 39800 45850
rect 40024 45610 40025 45850
rect 40605 45610 40606 46190
rect 40024 45609 40606 45610
rect 40740 45498 40760 46302
rect 40824 45498 40840 46302
rect 40740 45220 40840 45498
rect 41968 46302 42070 46318
rect 41968 45498 41984 46302
rect 42048 45498 42070 46302
rect 42202 46190 42784 46191
rect 42202 45610 42203 46190
rect 42783 45950 42784 46190
rect 43010 45950 45010 49390
rect 42783 45850 45010 45950
rect 42783 45610 42784 45850
rect 42202 45609 42784 45610
rect 41968 45482 42070 45498
rect 40740 45130 40750 45220
rect 40830 45130 40840 45220
rect 40740 45120 40840 45130
rect 41970 45220 42070 45482
rect 41970 45130 41980 45220
rect 42060 45130 42070 45220
rect 41970 45120 42070 45130
rect 43010 43010 45010 45850
rect 43000 39510 45010 43010
rect 40740 36422 40840 36440
rect 41970 36438 42070 36440
rect 40024 36310 40606 36311
rect 40024 36070 40025 36310
rect 37800 35970 40025 36070
rect 37800 26190 39800 35970
rect 40024 35730 40025 35970
rect 40605 35730 40606 36310
rect 40024 35729 40606 35730
rect 40740 35618 40760 36422
rect 40824 35618 40840 36422
rect 40740 35340 40840 35618
rect 41968 36422 42070 36438
rect 41968 35618 41984 36422
rect 42048 35618 42070 36422
rect 42202 36310 42784 36311
rect 42202 35730 42203 36310
rect 42783 36070 42784 36310
rect 43010 36070 45010 39510
rect 42783 35970 45010 36070
rect 42783 35730 42784 35970
rect 42202 35729 42784 35730
rect 41968 35602 42070 35618
rect 40740 35250 40750 35340
rect 40830 35250 40840 35340
rect 40740 35240 40840 35250
rect 41970 35340 42070 35602
rect 41970 35250 41980 35340
rect 42060 35250 42070 35340
rect 41970 35240 42070 35250
rect 43010 33130 45010 35970
rect 43000 29630 45010 33130
rect 40740 26542 40840 26560
rect 41970 26558 42070 26560
rect 40024 26430 40606 26431
rect 40024 26190 40025 26430
rect 37800 26090 40025 26190
rect 37800 16310 39800 26090
rect 40024 25850 40025 26090
rect 40605 25850 40606 26430
rect 40024 25849 40606 25850
rect 40740 25738 40760 26542
rect 40824 25738 40840 26542
rect 40740 25460 40840 25738
rect 41968 26542 42070 26558
rect 41968 25738 41984 26542
rect 42048 25738 42070 26542
rect 42202 26430 42784 26431
rect 42202 25850 42203 26430
rect 42783 26190 42784 26430
rect 43010 26190 45010 29630
rect 42783 26090 45010 26190
rect 42783 25850 42784 26090
rect 42202 25849 42784 25850
rect 41968 25722 42070 25738
rect 40740 25370 40750 25460
rect 40830 25370 40840 25460
rect 40740 25360 40840 25370
rect 41970 25460 42070 25722
rect 41970 25370 41980 25460
rect 42060 25370 42070 25460
rect 41970 25360 42070 25370
rect 43010 23250 45010 26090
rect 43000 19750 45010 23250
rect 40740 16662 40840 16680
rect 41970 16678 42070 16680
rect 40024 16550 40606 16551
rect 40024 16310 40025 16550
rect 37800 16210 40025 16310
rect 37800 6430 39800 16210
rect 40024 15970 40025 16210
rect 40605 15970 40606 16550
rect 40024 15969 40606 15970
rect 40740 15858 40760 16662
rect 40824 15858 40840 16662
rect 40740 15580 40840 15858
rect 41968 16662 42070 16678
rect 41968 15858 41984 16662
rect 42048 15858 42070 16662
rect 42202 16550 42784 16551
rect 42202 15970 42203 16550
rect 42783 16310 42784 16550
rect 43010 16310 45010 19750
rect 42783 16210 45010 16310
rect 42783 15970 42784 16210
rect 42202 15969 42784 15970
rect 41968 15842 42070 15858
rect 40740 15490 40750 15580
rect 40830 15490 40840 15580
rect 40740 15480 40840 15490
rect 41970 15580 42070 15842
rect 41970 15490 41980 15580
rect 42060 15490 42070 15580
rect 41970 15480 42070 15490
rect 43010 13370 45010 16210
rect 43000 9870 45010 13370
rect 40740 6782 40840 6800
rect 41970 6798 42070 6800
rect 40024 6670 40606 6671
rect 40024 6430 40025 6670
rect 37800 6330 40025 6430
rect 37800 -10 39800 6330
rect 40024 6090 40025 6330
rect 40605 6090 40606 6670
rect 40024 6089 40606 6090
rect 40740 5978 40760 6782
rect 40824 5978 40840 6782
rect 40740 5700 40840 5978
rect 41968 6782 42070 6798
rect 41968 5978 41984 6782
rect 42048 5978 42070 6782
rect 42202 6670 42784 6671
rect 42202 6090 42203 6670
rect 42783 6430 42784 6670
rect 43010 6430 45010 9870
rect 42783 6330 45010 6430
rect 42783 6090 42784 6330
rect 42202 6089 42784 6090
rect 41968 5962 42070 5978
rect 40740 5610 40750 5700
rect 40830 5610 40840 5700
rect 40740 5600 40840 5610
rect 41970 5700 42070 5962
rect 41970 5610 41980 5700
rect 42060 5610 42070 5700
rect 41970 5600 42070 5610
rect 43010 3490 45010 6330
rect 43000 -10 45010 3490
rect 47000 103780 49000 110790
rect 47000 101800 47010 103780
rect 48990 101800 49000 103780
rect 47000 65710 49000 101800
rect 52210 109790 54210 110790
rect 52210 107810 52220 109790
rect 54200 107810 54210 109790
rect 49940 66062 50040 66080
rect 51170 66078 51270 66080
rect 49224 65950 49806 65951
rect 49224 65710 49225 65950
rect 47000 65610 49225 65710
rect 47000 55830 49000 65610
rect 49224 65370 49225 65610
rect 49805 65370 49806 65950
rect 49224 65369 49806 65370
rect 49940 65258 49960 66062
rect 50024 65258 50040 66062
rect 49940 64980 50040 65258
rect 51168 66062 51270 66078
rect 51168 65258 51184 66062
rect 51248 65258 51270 66062
rect 51402 65950 51984 65951
rect 51402 65370 51403 65950
rect 51983 65710 51984 65950
rect 52210 65710 54210 107810
rect 51983 65610 54210 65710
rect 51983 65370 51984 65610
rect 51402 65369 51984 65370
rect 51168 65242 51270 65258
rect 49940 64890 49950 64980
rect 50030 64890 50040 64980
rect 49940 64880 50040 64890
rect 51170 64980 51270 65242
rect 51170 64890 51180 64980
rect 51260 64890 51270 64980
rect 51170 64880 51270 64890
rect 52210 62770 54210 65610
rect 52200 59270 54210 62770
rect 49940 56182 50040 56200
rect 51170 56198 51270 56200
rect 49224 56070 49806 56071
rect 49224 55830 49225 56070
rect 47000 55730 49225 55830
rect 47000 45950 49000 55730
rect 49224 55490 49225 55730
rect 49805 55490 49806 56070
rect 49224 55489 49806 55490
rect 49940 55378 49960 56182
rect 50024 55378 50040 56182
rect 49940 55100 50040 55378
rect 51168 56182 51270 56198
rect 51168 55378 51184 56182
rect 51248 55378 51270 56182
rect 51402 56070 51984 56071
rect 51402 55490 51403 56070
rect 51983 55830 51984 56070
rect 52210 55830 54210 59270
rect 51983 55730 54210 55830
rect 51983 55490 51984 55730
rect 51402 55489 51984 55490
rect 51168 55362 51270 55378
rect 49940 55010 49950 55100
rect 50030 55010 50040 55100
rect 49940 55000 50040 55010
rect 51170 55100 51270 55362
rect 51170 55010 51180 55100
rect 51260 55010 51270 55100
rect 51170 55000 51270 55010
rect 52210 52890 54210 55730
rect 52200 49390 54210 52890
rect 49940 46302 50040 46320
rect 51170 46318 51270 46320
rect 49224 46190 49806 46191
rect 49224 45950 49225 46190
rect 47000 45850 49225 45950
rect 47000 36070 49000 45850
rect 49224 45610 49225 45850
rect 49805 45610 49806 46190
rect 49224 45609 49806 45610
rect 49940 45498 49960 46302
rect 50024 45498 50040 46302
rect 49940 45220 50040 45498
rect 51168 46302 51270 46318
rect 51168 45498 51184 46302
rect 51248 45498 51270 46302
rect 51402 46190 51984 46191
rect 51402 45610 51403 46190
rect 51983 45950 51984 46190
rect 52210 45950 54210 49390
rect 51983 45850 54210 45950
rect 51983 45610 51984 45850
rect 51402 45609 51984 45610
rect 51168 45482 51270 45498
rect 49940 45130 49950 45220
rect 50030 45130 50040 45220
rect 49940 45120 50040 45130
rect 51170 45220 51270 45482
rect 51170 45130 51180 45220
rect 51260 45130 51270 45220
rect 51170 45120 51270 45130
rect 52210 43010 54210 45850
rect 52200 39510 54210 43010
rect 49940 36422 50040 36440
rect 51170 36438 51270 36440
rect 49224 36310 49806 36311
rect 49224 36070 49225 36310
rect 47000 35970 49225 36070
rect 47000 26190 49000 35970
rect 49224 35730 49225 35970
rect 49805 35730 49806 36310
rect 49224 35729 49806 35730
rect 49940 35618 49960 36422
rect 50024 35618 50040 36422
rect 49940 35340 50040 35618
rect 51168 36422 51270 36438
rect 51168 35618 51184 36422
rect 51248 35618 51270 36422
rect 51402 36310 51984 36311
rect 51402 35730 51403 36310
rect 51983 36070 51984 36310
rect 52210 36070 54210 39510
rect 51983 35970 54210 36070
rect 51983 35730 51984 35970
rect 51402 35729 51984 35730
rect 51168 35602 51270 35618
rect 49940 35250 49950 35340
rect 50030 35250 50040 35340
rect 49940 35240 50040 35250
rect 51170 35340 51270 35602
rect 51170 35250 51180 35340
rect 51260 35250 51270 35340
rect 51170 35240 51270 35250
rect 52210 33130 54210 35970
rect 52200 29630 54210 33130
rect 49940 26542 50040 26560
rect 51170 26558 51270 26560
rect 49224 26430 49806 26431
rect 49224 26190 49225 26430
rect 47000 26090 49225 26190
rect 47000 16310 49000 26090
rect 49224 25850 49225 26090
rect 49805 25850 49806 26430
rect 49224 25849 49806 25850
rect 49940 25738 49960 26542
rect 50024 25738 50040 26542
rect 49940 25460 50040 25738
rect 51168 26542 51270 26558
rect 51168 25738 51184 26542
rect 51248 25738 51270 26542
rect 51402 26430 51984 26431
rect 51402 25850 51403 26430
rect 51983 26190 51984 26430
rect 52210 26190 54210 29630
rect 51983 26090 54210 26190
rect 51983 25850 51984 26090
rect 51402 25849 51984 25850
rect 51168 25722 51270 25738
rect 49940 25370 49950 25460
rect 50030 25370 50040 25460
rect 49940 25360 50040 25370
rect 51170 25460 51270 25722
rect 51170 25370 51180 25460
rect 51260 25370 51270 25460
rect 51170 25360 51270 25370
rect 52210 23250 54210 26090
rect 52200 19750 54210 23250
rect 49940 16662 50040 16680
rect 51170 16678 51270 16680
rect 49224 16550 49806 16551
rect 49224 16310 49225 16550
rect 47000 16210 49225 16310
rect 47000 6430 49000 16210
rect 49224 15970 49225 16210
rect 49805 15970 49806 16550
rect 49224 15969 49806 15970
rect 49940 15858 49960 16662
rect 50024 15858 50040 16662
rect 49940 15580 50040 15858
rect 51168 16662 51270 16678
rect 51168 15858 51184 16662
rect 51248 15858 51270 16662
rect 51402 16550 51984 16551
rect 51402 15970 51403 16550
rect 51983 16310 51984 16550
rect 52210 16310 54210 19750
rect 51983 16210 54210 16310
rect 51983 15970 51984 16210
rect 51402 15969 51984 15970
rect 51168 15842 51270 15858
rect 49940 15490 49950 15580
rect 50030 15490 50040 15580
rect 49940 15480 50040 15490
rect 51170 15580 51270 15842
rect 51170 15490 51180 15580
rect 51260 15490 51270 15580
rect 51170 15480 51270 15490
rect 52210 13370 54210 16210
rect 52200 9870 54210 13370
rect 49940 6782 50040 6800
rect 51170 6798 51270 6800
rect 49224 6670 49806 6671
rect 49224 6430 49225 6670
rect 47000 6330 49225 6430
rect 47000 -10 49000 6330
rect 49224 6090 49225 6330
rect 49805 6090 49806 6670
rect 49224 6089 49806 6090
rect 49940 5978 49960 6782
rect 50024 5978 50040 6782
rect 49940 5700 50040 5978
rect 51168 6782 51270 6798
rect 51168 5978 51184 6782
rect 51248 5978 51270 6782
rect 51402 6670 51984 6671
rect 51402 6090 51403 6670
rect 51983 6430 51984 6670
rect 52210 6430 54210 9870
rect 51983 6330 54210 6430
rect 51983 6090 51984 6330
rect 51402 6089 51984 6090
rect 51168 5962 51270 5978
rect 49940 5610 49950 5700
rect 50030 5610 50040 5700
rect 49940 5600 50040 5610
rect 51170 5700 51270 5962
rect 51170 5610 51180 5700
rect 51260 5610 51270 5700
rect 51170 5600 51270 5610
rect 52210 3490 54210 6330
rect 52200 -10 54210 3490
rect 56200 103780 58200 110790
rect 56200 101800 56210 103780
rect 58190 101800 58200 103780
rect 56200 65710 58200 101800
rect 61410 109780 63410 110790
rect 61410 107800 61420 109780
rect 63400 107800 63410 109780
rect 59140 66062 59240 66080
rect 60370 66078 60470 66080
rect 58424 65950 59006 65951
rect 58424 65710 58425 65950
rect 56200 65610 58425 65710
rect 56200 55830 58200 65610
rect 58424 65370 58425 65610
rect 59005 65370 59006 65950
rect 58424 65369 59006 65370
rect 59140 65258 59160 66062
rect 59224 65258 59240 66062
rect 59140 64980 59240 65258
rect 60368 66062 60470 66078
rect 60368 65258 60384 66062
rect 60448 65258 60470 66062
rect 60602 65950 61184 65951
rect 60602 65370 60603 65950
rect 61183 65710 61184 65950
rect 61410 65710 63410 107800
rect 61183 65610 63410 65710
rect 61183 65370 61184 65610
rect 60602 65369 61184 65370
rect 60368 65242 60470 65258
rect 59140 64890 59150 64980
rect 59230 64890 59240 64980
rect 59140 64880 59240 64890
rect 60370 64980 60470 65242
rect 60370 64890 60380 64980
rect 60460 64890 60470 64980
rect 60370 64880 60470 64890
rect 61410 62770 63410 65610
rect 61400 59270 63410 62770
rect 59140 56182 59240 56200
rect 60370 56198 60470 56200
rect 58424 56070 59006 56071
rect 58424 55830 58425 56070
rect 56200 55730 58425 55830
rect 56200 45950 58200 55730
rect 58424 55490 58425 55730
rect 59005 55490 59006 56070
rect 58424 55489 59006 55490
rect 59140 55378 59160 56182
rect 59224 55378 59240 56182
rect 59140 55100 59240 55378
rect 60368 56182 60470 56198
rect 60368 55378 60384 56182
rect 60448 55378 60470 56182
rect 60602 56070 61184 56071
rect 60602 55490 60603 56070
rect 61183 55830 61184 56070
rect 61410 55830 63410 59270
rect 61183 55730 63410 55830
rect 61183 55490 61184 55730
rect 60602 55489 61184 55490
rect 60368 55362 60470 55378
rect 59140 55010 59150 55100
rect 59230 55010 59240 55100
rect 59140 55000 59240 55010
rect 60370 55100 60470 55362
rect 60370 55010 60380 55100
rect 60460 55010 60470 55100
rect 60370 55000 60470 55010
rect 61410 52890 63410 55730
rect 61400 49390 63410 52890
rect 59140 46302 59240 46320
rect 60370 46318 60470 46320
rect 58424 46190 59006 46191
rect 58424 45950 58425 46190
rect 56200 45850 58425 45950
rect 56200 36070 58200 45850
rect 58424 45610 58425 45850
rect 59005 45610 59006 46190
rect 58424 45609 59006 45610
rect 59140 45498 59160 46302
rect 59224 45498 59240 46302
rect 59140 45220 59240 45498
rect 60368 46302 60470 46318
rect 60368 45498 60384 46302
rect 60448 45498 60470 46302
rect 60602 46190 61184 46191
rect 60602 45610 60603 46190
rect 61183 45950 61184 46190
rect 61410 45950 63410 49390
rect 61183 45850 63410 45950
rect 61183 45610 61184 45850
rect 60602 45609 61184 45610
rect 60368 45482 60470 45498
rect 59140 45130 59150 45220
rect 59230 45130 59240 45220
rect 59140 45120 59240 45130
rect 60370 45220 60470 45482
rect 60370 45130 60380 45220
rect 60460 45130 60470 45220
rect 60370 45120 60470 45130
rect 61410 43010 63410 45850
rect 61400 39510 63410 43010
rect 59140 36422 59240 36440
rect 60370 36438 60470 36440
rect 58424 36310 59006 36311
rect 58424 36070 58425 36310
rect 56200 35970 58425 36070
rect 56200 26190 58200 35970
rect 58424 35730 58425 35970
rect 59005 35730 59006 36310
rect 58424 35729 59006 35730
rect 59140 35618 59160 36422
rect 59224 35618 59240 36422
rect 59140 35340 59240 35618
rect 60368 36422 60470 36438
rect 60368 35618 60384 36422
rect 60448 35618 60470 36422
rect 60602 36310 61184 36311
rect 60602 35730 60603 36310
rect 61183 36070 61184 36310
rect 61410 36070 63410 39510
rect 61183 35970 63410 36070
rect 61183 35730 61184 35970
rect 60602 35729 61184 35730
rect 60368 35602 60470 35618
rect 59140 35250 59150 35340
rect 59230 35250 59240 35340
rect 59140 35240 59240 35250
rect 60370 35340 60470 35602
rect 60370 35250 60380 35340
rect 60460 35250 60470 35340
rect 60370 35240 60470 35250
rect 61410 33130 63410 35970
rect 61400 29630 63410 33130
rect 59140 26542 59240 26560
rect 60370 26558 60470 26560
rect 58424 26430 59006 26431
rect 58424 26190 58425 26430
rect 56200 26090 58425 26190
rect 56200 16310 58200 26090
rect 58424 25850 58425 26090
rect 59005 25850 59006 26430
rect 58424 25849 59006 25850
rect 59140 25738 59160 26542
rect 59224 25738 59240 26542
rect 59140 25460 59240 25738
rect 60368 26542 60470 26558
rect 60368 25738 60384 26542
rect 60448 25738 60470 26542
rect 60602 26430 61184 26431
rect 60602 25850 60603 26430
rect 61183 26190 61184 26430
rect 61410 26190 63410 29630
rect 61183 26090 63410 26190
rect 61183 25850 61184 26090
rect 60602 25849 61184 25850
rect 60368 25722 60470 25738
rect 59140 25370 59150 25460
rect 59230 25370 59240 25460
rect 59140 25360 59240 25370
rect 60370 25460 60470 25722
rect 60370 25370 60380 25460
rect 60460 25370 60470 25460
rect 60370 25360 60470 25370
rect 61410 23250 63410 26090
rect 61400 19750 63410 23250
rect 59140 16662 59240 16680
rect 60370 16678 60470 16680
rect 58424 16550 59006 16551
rect 58424 16310 58425 16550
rect 56200 16210 58425 16310
rect 56200 6430 58200 16210
rect 58424 15970 58425 16210
rect 59005 15970 59006 16550
rect 58424 15969 59006 15970
rect 59140 15858 59160 16662
rect 59224 15858 59240 16662
rect 59140 15580 59240 15858
rect 60368 16662 60470 16678
rect 60368 15858 60384 16662
rect 60448 15858 60470 16662
rect 60602 16550 61184 16551
rect 60602 15970 60603 16550
rect 61183 16310 61184 16550
rect 61410 16310 63410 19750
rect 61183 16210 63410 16310
rect 61183 15970 61184 16210
rect 60602 15969 61184 15970
rect 60368 15842 60470 15858
rect 59140 15490 59150 15580
rect 59230 15490 59240 15580
rect 59140 15480 59240 15490
rect 60370 15580 60470 15842
rect 60370 15490 60380 15580
rect 60460 15490 60470 15580
rect 60370 15480 60470 15490
rect 61410 13370 63410 16210
rect 61400 9870 63410 13370
rect 59140 6782 59240 6800
rect 60370 6798 60470 6800
rect 58424 6670 59006 6671
rect 58424 6430 58425 6670
rect 56200 6330 58425 6430
rect 56200 -10 58200 6330
rect 58424 6090 58425 6330
rect 59005 6090 59006 6670
rect 58424 6089 59006 6090
rect 59140 5978 59160 6782
rect 59224 5978 59240 6782
rect 59140 5700 59240 5978
rect 60368 6782 60470 6798
rect 60368 5978 60384 6782
rect 60448 5978 60470 6782
rect 60602 6670 61184 6671
rect 60602 6090 60603 6670
rect 61183 6430 61184 6670
rect 61410 6430 63410 9870
rect 61183 6330 63410 6430
rect 61183 6090 61184 6330
rect 60602 6089 61184 6090
rect 60368 5962 60470 5978
rect 59140 5610 59150 5700
rect 59230 5610 59240 5700
rect 59140 5600 59240 5610
rect 60370 5700 60470 5962
rect 60370 5610 60380 5700
rect 60460 5610 60470 5700
rect 60370 5600 60470 5610
rect 61410 3490 63410 6330
rect 61400 -10 63410 3490
rect 65400 103780 67400 110790
rect 65400 101800 65410 103780
rect 67390 101800 67400 103780
rect 65400 65710 67400 101800
rect 70610 109780 72610 110790
rect 70610 107800 70620 109780
rect 72600 107800 72610 109780
rect 68340 66062 68440 66080
rect 69570 66078 69670 66080
rect 67624 65950 68206 65951
rect 67624 65710 67625 65950
rect 65400 65610 67625 65710
rect 65400 55830 67400 65610
rect 67624 65370 67625 65610
rect 68205 65370 68206 65950
rect 67624 65369 68206 65370
rect 68340 65258 68360 66062
rect 68424 65258 68440 66062
rect 68340 64980 68440 65258
rect 69568 66062 69670 66078
rect 69568 65258 69584 66062
rect 69648 65258 69670 66062
rect 69802 65950 70384 65951
rect 69802 65370 69803 65950
rect 70383 65710 70384 65950
rect 70610 65710 72610 107800
rect 70383 65610 72610 65710
rect 70383 65370 70384 65610
rect 69802 65369 70384 65370
rect 69568 65242 69670 65258
rect 68340 64890 68350 64980
rect 68430 64890 68440 64980
rect 68340 64880 68440 64890
rect 69570 64980 69670 65242
rect 69570 64890 69580 64980
rect 69660 64890 69670 64980
rect 69570 64880 69670 64890
rect 70610 62770 72610 65610
rect 70600 59270 72610 62770
rect 68340 56182 68440 56200
rect 69570 56198 69670 56200
rect 67624 56070 68206 56071
rect 67624 55830 67625 56070
rect 65400 55730 67625 55830
rect 65400 45950 67400 55730
rect 67624 55490 67625 55730
rect 68205 55490 68206 56070
rect 67624 55489 68206 55490
rect 68340 55378 68360 56182
rect 68424 55378 68440 56182
rect 68340 55100 68440 55378
rect 69568 56182 69670 56198
rect 69568 55378 69584 56182
rect 69648 55378 69670 56182
rect 69802 56070 70384 56071
rect 69802 55490 69803 56070
rect 70383 55830 70384 56070
rect 70610 55830 72610 59270
rect 70383 55730 72610 55830
rect 70383 55490 70384 55730
rect 69802 55489 70384 55490
rect 69568 55362 69670 55378
rect 68340 55010 68350 55100
rect 68430 55010 68440 55100
rect 68340 55000 68440 55010
rect 69570 55100 69670 55362
rect 69570 55010 69580 55100
rect 69660 55010 69670 55100
rect 69570 55000 69670 55010
rect 70610 52890 72610 55730
rect 70600 49390 72610 52890
rect 68340 46302 68440 46320
rect 69570 46318 69670 46320
rect 67624 46190 68206 46191
rect 67624 45950 67625 46190
rect 65400 45850 67625 45950
rect 65400 36070 67400 45850
rect 67624 45610 67625 45850
rect 68205 45610 68206 46190
rect 67624 45609 68206 45610
rect 68340 45498 68360 46302
rect 68424 45498 68440 46302
rect 68340 45220 68440 45498
rect 69568 46302 69670 46318
rect 69568 45498 69584 46302
rect 69648 45498 69670 46302
rect 69802 46190 70384 46191
rect 69802 45610 69803 46190
rect 70383 45950 70384 46190
rect 70610 45950 72610 49390
rect 70383 45850 72610 45950
rect 70383 45610 70384 45850
rect 69802 45609 70384 45610
rect 69568 45482 69670 45498
rect 68340 45130 68350 45220
rect 68430 45130 68440 45220
rect 68340 45120 68440 45130
rect 69570 45220 69670 45482
rect 69570 45130 69580 45220
rect 69660 45130 69670 45220
rect 69570 45120 69670 45130
rect 70610 43010 72610 45850
rect 70600 39510 72610 43010
rect 68340 36422 68440 36440
rect 69570 36438 69670 36440
rect 67624 36310 68206 36311
rect 67624 36070 67625 36310
rect 65400 35970 67625 36070
rect 65400 26190 67400 35970
rect 67624 35730 67625 35970
rect 68205 35730 68206 36310
rect 67624 35729 68206 35730
rect 68340 35618 68360 36422
rect 68424 35618 68440 36422
rect 68340 35340 68440 35618
rect 69568 36422 69670 36438
rect 69568 35618 69584 36422
rect 69648 35618 69670 36422
rect 69802 36310 70384 36311
rect 69802 35730 69803 36310
rect 70383 36070 70384 36310
rect 70610 36070 72610 39510
rect 70383 35970 72610 36070
rect 70383 35730 70384 35970
rect 69802 35729 70384 35730
rect 69568 35602 69670 35618
rect 68340 35250 68350 35340
rect 68430 35250 68440 35340
rect 68340 35240 68440 35250
rect 69570 35340 69670 35602
rect 69570 35250 69580 35340
rect 69660 35250 69670 35340
rect 69570 35240 69670 35250
rect 70610 33130 72610 35970
rect 70600 29630 72610 33130
rect 68340 26542 68440 26560
rect 69570 26558 69670 26560
rect 67624 26430 68206 26431
rect 67624 26190 67625 26430
rect 65400 26090 67625 26190
rect 65400 16310 67400 26090
rect 67624 25850 67625 26090
rect 68205 25850 68206 26430
rect 67624 25849 68206 25850
rect 68340 25738 68360 26542
rect 68424 25738 68440 26542
rect 68340 25460 68440 25738
rect 69568 26542 69670 26558
rect 69568 25738 69584 26542
rect 69648 25738 69670 26542
rect 69802 26430 70384 26431
rect 69802 25850 69803 26430
rect 70383 26190 70384 26430
rect 70610 26190 72610 29630
rect 70383 26090 72610 26190
rect 70383 25850 70384 26090
rect 69802 25849 70384 25850
rect 69568 25722 69670 25738
rect 68340 25370 68350 25460
rect 68430 25370 68440 25460
rect 68340 25360 68440 25370
rect 69570 25460 69670 25722
rect 69570 25370 69580 25460
rect 69660 25370 69670 25460
rect 69570 25360 69670 25370
rect 70610 23250 72610 26090
rect 70600 19750 72610 23250
rect 68340 16662 68440 16680
rect 69570 16678 69670 16680
rect 67624 16550 68206 16551
rect 67624 16310 67625 16550
rect 65400 16210 67625 16310
rect 65400 6430 67400 16210
rect 67624 15970 67625 16210
rect 68205 15970 68206 16550
rect 67624 15969 68206 15970
rect 68340 15858 68360 16662
rect 68424 15858 68440 16662
rect 68340 15580 68440 15858
rect 69568 16662 69670 16678
rect 69568 15858 69584 16662
rect 69648 15858 69670 16662
rect 69802 16550 70384 16551
rect 69802 15970 69803 16550
rect 70383 16310 70384 16550
rect 70610 16310 72610 19750
rect 70383 16210 72610 16310
rect 70383 15970 70384 16210
rect 69802 15969 70384 15970
rect 69568 15842 69670 15858
rect 68340 15490 68350 15580
rect 68430 15490 68440 15580
rect 68340 15480 68440 15490
rect 69570 15580 69670 15842
rect 69570 15490 69580 15580
rect 69660 15490 69670 15580
rect 69570 15480 69670 15490
rect 70610 13370 72610 16210
rect 70600 9870 72610 13370
rect 68340 6782 68440 6800
rect 69570 6798 69670 6800
rect 67624 6670 68206 6671
rect 67624 6430 67625 6670
rect 65400 6330 67625 6430
rect 65400 -10 67400 6330
rect 67624 6090 67625 6330
rect 68205 6090 68206 6670
rect 67624 6089 68206 6090
rect 68340 5978 68360 6782
rect 68424 5978 68440 6782
rect 68340 5700 68440 5978
rect 69568 6782 69670 6798
rect 69568 5978 69584 6782
rect 69648 5978 69670 6782
rect 69802 6670 70384 6671
rect 69802 6090 69803 6670
rect 70383 6430 70384 6670
rect 70610 6430 72610 9870
rect 70383 6330 72610 6430
rect 70383 6090 70384 6330
rect 69802 6089 70384 6090
rect 69568 5962 69670 5978
rect 68340 5610 68350 5700
rect 68430 5610 68440 5700
rect 68340 5600 68440 5610
rect 69570 5700 69670 5962
rect 69570 5610 69580 5700
rect 69660 5610 69670 5700
rect 69570 5600 69670 5610
rect 70610 3490 72610 6330
rect 70600 -10 72610 3490
<< res0p35 >>
rect 4174 95316 4248 95520
rect 4912 95316 4986 95520
rect 4174 85436 4248 85640
rect 4912 85436 4986 85640
rect 13374 85436 13448 85640
rect 14112 85436 14186 85640
rect 4174 75556 4248 75760
rect 4912 75556 4986 75760
rect 13374 75556 13448 75760
rect 14112 75556 14186 75760
rect 22574 75556 22648 75760
rect 23312 75556 23386 75760
rect 31774 75556 31848 75760
rect 32512 75556 32586 75760
rect 4174 65676 4248 65880
rect 4912 65676 4986 65880
rect 13374 65676 13448 65880
rect 14112 65676 14186 65880
rect 22574 65676 22648 65880
rect 23312 65676 23386 65880
rect 31774 65676 31848 65880
rect 32512 65676 32586 65880
rect 40974 65676 41048 65880
rect 41712 65676 41786 65880
rect 50174 65676 50248 65880
rect 50912 65676 50986 65880
rect 59374 65676 59448 65880
rect 60112 65676 60186 65880
rect 68574 65676 68648 65880
rect 69312 65676 69386 65880
rect 4174 55796 4248 56000
rect 4912 55796 4986 56000
rect 13374 55796 13448 56000
rect 14112 55796 14186 56000
rect 22574 55796 22648 56000
rect 23312 55796 23386 56000
rect 31774 55796 31848 56000
rect 32512 55796 32586 56000
rect 40974 55796 41048 56000
rect 41712 55796 41786 56000
rect 50174 55796 50248 56000
rect 50912 55796 50986 56000
rect 59374 55796 59448 56000
rect 60112 55796 60186 56000
rect 68574 55796 68648 56000
rect 69312 55796 69386 56000
rect 4174 45916 4248 46120
rect 4912 45916 4986 46120
rect 13374 45916 13448 46120
rect 14112 45916 14186 46120
rect 22574 45916 22648 46120
rect 23312 45916 23386 46120
rect 31774 45916 31848 46120
rect 32512 45916 32586 46120
rect 40974 45916 41048 46120
rect 41712 45916 41786 46120
rect 50174 45916 50248 46120
rect 50912 45916 50986 46120
rect 59374 45916 59448 46120
rect 60112 45916 60186 46120
rect 68574 45916 68648 46120
rect 69312 45916 69386 46120
rect 4174 36036 4248 36240
rect 4912 36036 4986 36240
rect 13374 36036 13448 36240
rect 14112 36036 14186 36240
rect 22574 36036 22648 36240
rect 23312 36036 23386 36240
rect 31774 36036 31848 36240
rect 32512 36036 32586 36240
rect 40974 36036 41048 36240
rect 41712 36036 41786 36240
rect 50174 36036 50248 36240
rect 50912 36036 50986 36240
rect 59374 36036 59448 36240
rect 60112 36036 60186 36240
rect 68574 36036 68648 36240
rect 69312 36036 69386 36240
rect 4174 26156 4248 26360
rect 4912 26156 4986 26360
rect 13374 26156 13448 26360
rect 14112 26156 14186 26360
rect 22574 26156 22648 26360
rect 23312 26156 23386 26360
rect 31774 26156 31848 26360
rect 32512 26156 32586 26360
rect 40974 26156 41048 26360
rect 41712 26156 41786 26360
rect 50174 26156 50248 26360
rect 50912 26156 50986 26360
rect 59374 26156 59448 26360
rect 60112 26156 60186 26360
rect 68574 26156 68648 26360
rect 69312 26156 69386 26360
rect 4174 16276 4248 16480
rect 4912 16276 4986 16480
rect 13374 16276 13448 16480
rect 14112 16276 14186 16480
rect 22574 16276 22648 16480
rect 23312 16276 23386 16480
rect 31774 16276 31848 16480
rect 32512 16276 32586 16480
rect 40974 16276 41048 16480
rect 41712 16276 41786 16480
rect 50174 16276 50248 16480
rect 50912 16276 50986 16480
rect 59374 16276 59448 16480
rect 60112 16276 60186 16480
rect 68574 16276 68648 16480
rect 69312 16276 69386 16480
rect 4174 6396 4248 6600
rect 4912 6396 4986 6600
rect 13374 6396 13448 6600
rect 14112 6396 14186 6600
rect 22574 6396 22648 6600
rect 23312 6396 23386 6600
rect 31774 6396 31848 6600
rect 32512 6396 32586 6600
rect 40974 6396 41048 6600
rect 41712 6396 41786 6600
rect 50174 6396 50248 6600
rect 50912 6396 50986 6600
rect 59374 6396 59448 6600
rect 60112 6396 60186 6600
rect 68574 6396 68648 6600
rect 69312 6396 69386 6600
<< labels >>
flabel metal3 -9760 102720 -9760 102720 3 FreeSans 2400 0 0 0 OUT_P
port 1 e
flabel metal3 82600 108800 82600 108800 7 FreeSans 2400 0 0 0 OUT_N
port 2 w
flabel metal2 82600 93460 82600 93460 7 FreeSans 2400 0 0 0 bit0
port 3 w
flabel metal2 82600 83500 82600 83500 7 FreeSans 2400 0 0 0 bit1
port 4 w
flabel metal2 82600 73590 82600 73590 7 FreeSans 2400 0 0 0 bit2
port 5 w
flabel metal2 82600 63750 82600 63750 7 FreeSans 2400 0 0 0 bit3
port 6 w
flabel metal2 82600 43930 82600 43930 7 FreeSans 2400 0 0 0 bit4
port 7 w
flabel metal2 82600 4390 82600 4390 7 FreeSans 2400 0 0 0 bit5
port 8 w
flabel metal2 -5980 110790 -5980 110790 5 FreeSans 2400 0 0 0 VDD
port 9 s
flabel metal1 -2890 110790 -2890 110790 5 FreeSans 2400 0 0 0 GND
port 10 s
flabel metal1 -610 5890 -610 5890 1 FreeSans 400 0 0 0 inv_1_0/OUT
flabel metal2 -110 5840 -110 5840 1 FreeSans 400 0 0 0 inv_1_0/ON
flabel metal2 -5820 9870 -5820 9870 5 FreeSans 2400 0 0 0 inv_1_0/VDD
flabel metal1 -2820 9870 -2820 9870 5 FreeSans 2400 0 0 0 inv_1_0/GND
flabel metal2 9200 14330 9200 14330 7 FreeSans 2400 0 0 0 cell_unit_8/ON
flabel metal1 9200 17690 9200 17690 7 FreeSans 2400 0 0 0 cell_unit_8/V_bias
flabel metal4 1950 19750 1950 19750 5 FreeSans 2400 0 0 0 cell_unit_8/OUT_P
flabel metal4 7210 19750 7210 19750 5 FreeSans 2400 0 0 0 cell_unit_8/OUT_N
flabel metal1 9200 11870 9200 11870 7 FreeSans 2400 0 0 0 cell_unit_8/GND
flabel metal2 4328 16112 4348 16240 7 FreeSans 300 180 0 0 cell_unit_8/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 15934 4348 16062 7 FreeSans 300 180 0 0 cell_unit_8/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 16278 4681 16344 0 FreeSans 300 0 0 0 cell_unit_8/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 15934 4412 15950 3 FreeSans 300 90 0 0 cell_unit_8/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 15830 4681 15896 0 FreeSans 300 0 0 0 cell_unit_8/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 15934 4806 15950 3 FreeSans 300 90 0 0 cell_unit_8/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 9200 4450 9200 4450 7 FreeSans 2400 0 0 0 cell_unit_0/ON
flabel metal1 9200 7810 9200 7810 7 FreeSans 2400 0 0 0 cell_unit_0/V_bias
flabel metal4 1950 9870 1950 9870 5 FreeSans 2400 0 0 0 cell_unit_0/OUT_P
flabel metal4 7210 9870 7210 9870 5 FreeSans 2400 0 0 0 cell_unit_0/OUT_N
flabel metal1 9200 1990 9200 1990 7 FreeSans 2400 0 0 0 cell_unit_0/GND
flabel metal2 4328 6232 4348 6360 7 FreeSans 300 180 0 0 cell_unit_0/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 6054 4348 6182 7 FreeSans 300 180 0 0 cell_unit_0/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 6398 4681 6464 0 FreeSans 300 0 0 0 cell_unit_0/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 6054 4412 6070 3 FreeSans 300 90 0 0 cell_unit_0/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 5950 4681 6016 0 FreeSans 300 0 0 0 cell_unit_0/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 6054 4806 6070 3 FreeSans 300 90 0 0 cell_unit_0/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 14330 18400 14330 7 FreeSans 2400 0 0 0 cell_unit_11/ON
flabel metal1 18400 17690 18400 17690 7 FreeSans 2400 0 0 0 cell_unit_11/V_bias
flabel metal4 11150 19750 11150 19750 5 FreeSans 2400 0 0 0 cell_unit_11/OUT_P
flabel metal4 16410 19750 16410 19750 5 FreeSans 2400 0 0 0 cell_unit_11/OUT_N
flabel metal1 18400 11870 18400 11870 7 FreeSans 2400 0 0 0 cell_unit_11/GND
flabel metal2 13528 16112 13548 16240 7 FreeSans 300 180 0 0 cell_unit_11/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 15934 13548 16062 7 FreeSans 300 180 0 0 cell_unit_11/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 16278 13881 16344 0 FreeSans 300 0 0 0 cell_unit_11/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 15934 13612 15950 3 FreeSans 300 90 0 0 cell_unit_11/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 15830 13881 15896 0 FreeSans 300 0 0 0 cell_unit_11/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 15934 14006 15950 3 FreeSans 300 90 0 0 cell_unit_11/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 4450 18400 4450 7 FreeSans 2400 0 0 0 cell_unit_1/ON
flabel metal1 18400 7810 18400 7810 7 FreeSans 2400 0 0 0 cell_unit_1/V_bias
flabel metal4 11150 9870 11150 9870 5 FreeSans 2400 0 0 0 cell_unit_1/OUT_P
flabel metal4 16410 9870 16410 9870 5 FreeSans 2400 0 0 0 cell_unit_1/OUT_N
flabel metal1 18400 1990 18400 1990 7 FreeSans 2400 0 0 0 cell_unit_1/GND
flabel metal2 13528 6232 13548 6360 7 FreeSans 300 180 0 0 cell_unit_1/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 6054 13548 6182 7 FreeSans 300 180 0 0 cell_unit_1/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 6398 13881 6464 0 FreeSans 300 0 0 0 cell_unit_1/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 6054 13612 6070 3 FreeSans 300 90 0 0 cell_unit_1/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 5950 13881 6016 0 FreeSans 300 0 0 0 cell_unit_1/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 6054 14006 6070 3 FreeSans 300 90 0 0 cell_unit_1/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 14330 27600 14330 7 FreeSans 2400 0 0 0 cell_unit_12/ON
flabel metal1 27600 17690 27600 17690 7 FreeSans 2400 0 0 0 cell_unit_12/V_bias
flabel metal4 20350 19750 20350 19750 5 FreeSans 2400 0 0 0 cell_unit_12/OUT_P
flabel metal4 25610 19750 25610 19750 5 FreeSans 2400 0 0 0 cell_unit_12/OUT_N
flabel metal1 27600 11870 27600 11870 7 FreeSans 2400 0 0 0 cell_unit_12/GND
flabel metal2 22728 16112 22748 16240 7 FreeSans 300 180 0 0 cell_unit_12/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 15934 22748 16062 7 FreeSans 300 180 0 0 cell_unit_12/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 16278 23081 16344 0 FreeSans 300 0 0 0 cell_unit_12/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 15934 22812 15950 3 FreeSans 300 90 0 0 cell_unit_12/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 15830 23081 15896 0 FreeSans 300 0 0 0 cell_unit_12/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 15934 23206 15950 3 FreeSans 300 90 0 0 cell_unit_12/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 4450 27600 4450 7 FreeSans 2400 0 0 0 cell_unit_2/ON
flabel metal1 27600 7810 27600 7810 7 FreeSans 2400 0 0 0 cell_unit_2/V_bias
flabel metal4 20350 9870 20350 9870 5 FreeSans 2400 0 0 0 cell_unit_2/OUT_P
flabel metal4 25610 9870 25610 9870 5 FreeSans 2400 0 0 0 cell_unit_2/OUT_N
flabel metal1 27600 1990 27600 1990 7 FreeSans 2400 0 0 0 cell_unit_2/GND
flabel metal2 22728 6232 22748 6360 7 FreeSans 300 180 0 0 cell_unit_2/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 6054 22748 6182 7 FreeSans 300 180 0 0 cell_unit_2/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 6398 23081 6464 0 FreeSans 300 0 0 0 cell_unit_2/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 6054 22812 6070 3 FreeSans 300 90 0 0 cell_unit_2/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 5950 23081 6016 0 FreeSans 300 0 0 0 cell_unit_2/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 6054 23206 6070 3 FreeSans 300 90 0 0 cell_unit_2/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 14330 36800 14330 7 FreeSans 2400 0 0 0 cell_unit_13/ON
flabel metal1 36800 17690 36800 17690 7 FreeSans 2400 0 0 0 cell_unit_13/V_bias
flabel metal4 29550 19750 29550 19750 5 FreeSans 2400 0 0 0 cell_unit_13/OUT_P
flabel metal4 34810 19750 34810 19750 5 FreeSans 2400 0 0 0 cell_unit_13/OUT_N
flabel metal1 36800 11870 36800 11870 7 FreeSans 2400 0 0 0 cell_unit_13/GND
flabel metal2 31928 16112 31948 16240 7 FreeSans 300 180 0 0 cell_unit_13/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 15934 31948 16062 7 FreeSans 300 180 0 0 cell_unit_13/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 16278 32281 16344 0 FreeSans 300 0 0 0 cell_unit_13/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 15934 32012 15950 3 FreeSans 300 90 0 0 cell_unit_13/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 15830 32281 15896 0 FreeSans 300 0 0 0 cell_unit_13/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 15934 32406 15950 3 FreeSans 300 90 0 0 cell_unit_13/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 4450 36800 4450 7 FreeSans 2400 0 0 0 cell_unit_3/ON
flabel metal1 36800 7810 36800 7810 7 FreeSans 2400 0 0 0 cell_unit_3/V_bias
flabel metal4 29550 9870 29550 9870 5 FreeSans 2400 0 0 0 cell_unit_3/OUT_P
flabel metal4 34810 9870 34810 9870 5 FreeSans 2400 0 0 0 cell_unit_3/OUT_N
flabel metal1 36800 1990 36800 1990 7 FreeSans 2400 0 0 0 cell_unit_3/GND
flabel metal2 31928 6232 31948 6360 7 FreeSans 300 180 0 0 cell_unit_3/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 6054 31948 6182 7 FreeSans 300 180 0 0 cell_unit_3/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 6398 32281 6464 0 FreeSans 300 0 0 0 cell_unit_3/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 6054 32012 6070 3 FreeSans 300 90 0 0 cell_unit_3/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 5950 32281 6016 0 FreeSans 300 0 0 0 cell_unit_3/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 6054 32406 6070 3 FreeSans 300 90 0 0 cell_unit_3/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 14330 55200 14330 7 FreeSans 2400 0 0 0 cell_unit_15/ON
flabel metal1 55200 17690 55200 17690 7 FreeSans 2400 0 0 0 cell_unit_15/V_bias
flabel metal4 47950 19750 47950 19750 5 FreeSans 2400 0 0 0 cell_unit_15/OUT_P
flabel metal4 53210 19750 53210 19750 5 FreeSans 2400 0 0 0 cell_unit_15/OUT_N
flabel metal1 55200 11870 55200 11870 7 FreeSans 2400 0 0 0 cell_unit_15/GND
flabel metal2 50328 16112 50348 16240 7 FreeSans 300 180 0 0 cell_unit_15/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 15934 50348 16062 7 FreeSans 300 180 0 0 cell_unit_15/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 16278 50681 16344 0 FreeSans 300 0 0 0 cell_unit_15/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 15934 50412 15950 3 FreeSans 300 90 0 0 cell_unit_15/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 15830 50681 15896 0 FreeSans 300 0 0 0 cell_unit_15/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 15934 50806 15950 3 FreeSans 300 90 0 0 cell_unit_15/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 14330 46000 14330 7 FreeSans 2400 0 0 0 cell_unit_14/ON
flabel metal1 46000 17690 46000 17690 7 FreeSans 2400 0 0 0 cell_unit_14/V_bias
flabel metal4 38750 19750 38750 19750 5 FreeSans 2400 0 0 0 cell_unit_14/OUT_P
flabel metal4 44010 19750 44010 19750 5 FreeSans 2400 0 0 0 cell_unit_14/OUT_N
flabel metal1 46000 11870 46000 11870 7 FreeSans 2400 0 0 0 cell_unit_14/GND
flabel metal2 41128 16112 41148 16240 7 FreeSans 300 180 0 0 cell_unit_14/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 15934 41148 16062 7 FreeSans 300 180 0 0 cell_unit_14/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 16278 41481 16344 0 FreeSans 300 0 0 0 cell_unit_14/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 15934 41212 15950 3 FreeSans 300 90 0 0 cell_unit_14/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 15830 41481 15896 0 FreeSans 300 0 0 0 cell_unit_14/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 15934 41606 15950 3 FreeSans 300 90 0 0 cell_unit_14/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 4450 55200 4450 7 FreeSans 2400 0 0 0 cell_unit_5/ON
flabel metal1 55200 7810 55200 7810 7 FreeSans 2400 0 0 0 cell_unit_5/V_bias
flabel metal4 47950 9870 47950 9870 5 FreeSans 2400 0 0 0 cell_unit_5/OUT_P
flabel metal4 53210 9870 53210 9870 5 FreeSans 2400 0 0 0 cell_unit_5/OUT_N
flabel metal1 55200 1990 55200 1990 7 FreeSans 2400 0 0 0 cell_unit_5/GND
flabel metal2 50328 6232 50348 6360 7 FreeSans 300 180 0 0 cell_unit_5/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 6054 50348 6182 7 FreeSans 300 180 0 0 cell_unit_5/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 6398 50681 6464 0 FreeSans 300 0 0 0 cell_unit_5/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 6054 50412 6070 3 FreeSans 300 90 0 0 cell_unit_5/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 5950 50681 6016 0 FreeSans 300 0 0 0 cell_unit_5/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 6054 50806 6070 3 FreeSans 300 90 0 0 cell_unit_5/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 4450 46000 4450 7 FreeSans 2400 0 0 0 cell_unit_4/ON
flabel metal1 46000 7810 46000 7810 7 FreeSans 2400 0 0 0 cell_unit_4/V_bias
flabel metal4 38750 9870 38750 9870 5 FreeSans 2400 0 0 0 cell_unit_4/OUT_P
flabel metal4 44010 9870 44010 9870 5 FreeSans 2400 0 0 0 cell_unit_4/OUT_N
flabel metal1 46000 1990 46000 1990 7 FreeSans 2400 0 0 0 cell_unit_4/GND
flabel metal2 41128 6232 41148 6360 7 FreeSans 300 180 0 0 cell_unit_4/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 6054 41148 6182 7 FreeSans 300 180 0 0 cell_unit_4/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 6398 41481 6464 0 FreeSans 300 0 0 0 cell_unit_4/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 6054 41212 6070 3 FreeSans 300 90 0 0 cell_unit_4/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 5950 41481 6016 0 FreeSans 300 0 0 0 cell_unit_4/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 6054 41606 6070 3 FreeSans 300 90 0 0 cell_unit_4/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 14330 64400 14330 7 FreeSans 2400 0 0 0 cell_unit_16/ON
flabel metal1 64400 17690 64400 17690 7 FreeSans 2400 0 0 0 cell_unit_16/V_bias
flabel metal4 57150 19750 57150 19750 5 FreeSans 2400 0 0 0 cell_unit_16/OUT_P
flabel metal4 62410 19750 62410 19750 5 FreeSans 2400 0 0 0 cell_unit_16/OUT_N
flabel metal1 64400 11870 64400 11870 7 FreeSans 2400 0 0 0 cell_unit_16/GND
flabel metal2 59528 16112 59548 16240 7 FreeSans 300 180 0 0 cell_unit_16/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 15934 59548 16062 7 FreeSans 300 180 0 0 cell_unit_16/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 16278 59881 16344 0 FreeSans 300 0 0 0 cell_unit_16/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 15934 59612 15950 3 FreeSans 300 90 0 0 cell_unit_16/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 15830 59881 15896 0 FreeSans 300 0 0 0 cell_unit_16/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 15934 60006 15950 3 FreeSans 300 90 0 0 cell_unit_16/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 4450 64400 4450 7 FreeSans 2400 0 0 0 cell_unit_6/ON
flabel metal1 64400 7810 64400 7810 7 FreeSans 2400 0 0 0 cell_unit_6/V_bias
flabel metal4 57150 9870 57150 9870 5 FreeSans 2400 0 0 0 cell_unit_6/OUT_P
flabel metal4 62410 9870 62410 9870 5 FreeSans 2400 0 0 0 cell_unit_6/OUT_N
flabel metal1 64400 1990 64400 1990 7 FreeSans 2400 0 0 0 cell_unit_6/GND
flabel metal2 59528 6232 59548 6360 7 FreeSans 300 180 0 0 cell_unit_6/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 6054 59548 6182 7 FreeSans 300 180 0 0 cell_unit_6/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 6398 59881 6464 0 FreeSans 300 0 0 0 cell_unit_6/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 6054 59612 6070 3 FreeSans 300 90 0 0 cell_unit_6/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 5950 59881 6016 0 FreeSans 300 0 0 0 cell_unit_6/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 6054 60006 6070 3 FreeSans 300 90 0 0 cell_unit_6/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 14330 73600 14330 7 FreeSans 2400 0 0 0 cell_unit_17/ON
flabel metal1 73600 17690 73600 17690 7 FreeSans 2400 0 0 0 cell_unit_17/V_bias
flabel metal4 66350 19750 66350 19750 5 FreeSans 2400 0 0 0 cell_unit_17/OUT_P
flabel metal4 71610 19750 71610 19750 5 FreeSans 2400 0 0 0 cell_unit_17/OUT_N
flabel metal1 73600 11870 73600 11870 7 FreeSans 2400 0 0 0 cell_unit_17/GND
flabel metal2 68728 16112 68748 16240 7 FreeSans 300 180 0 0 cell_unit_17/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 15934 68748 16062 7 FreeSans 300 180 0 0 cell_unit_17/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 16278 69081 16344 0 FreeSans 300 0 0 0 cell_unit_17/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 15934 68812 15950 3 FreeSans 300 90 0 0 cell_unit_17/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 15830 69081 15896 0 FreeSans 300 0 0 0 cell_unit_17/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 15934 69206 15950 3 FreeSans 300 90 0 0 cell_unit_17/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 4450 73600 4450 7 FreeSans 2400 0 0 0 cell_unit_7/ON
flabel metal1 73600 7810 73600 7810 7 FreeSans 2400 0 0 0 cell_unit_7/V_bias
flabel metal4 66350 9870 66350 9870 5 FreeSans 2400 0 0 0 cell_unit_7/OUT_P
flabel metal4 71610 9870 71610 9870 5 FreeSans 2400 0 0 0 cell_unit_7/OUT_N
flabel metal1 73600 1990 73600 1990 7 FreeSans 2400 0 0 0 cell_unit_7/GND
flabel metal2 68728 6232 68748 6360 7 FreeSans 300 180 0 0 cell_unit_7/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 6054 68748 6182 7 FreeSans 300 180 0 0 cell_unit_7/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 6398 69081 6464 0 FreeSans 300 0 0 0 cell_unit_7/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 6054 68812 6070 3 FreeSans 300 90 0 0 cell_unit_7/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 5950 69081 6016 0 FreeSans 300 0 0 0 cell_unit_7/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 6054 69206 6070 3 FreeSans 300 90 0 0 cell_unit_7/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 9200 24210 9200 24210 7 FreeSans 2400 0 0 0 cell_unit_9/ON
flabel metal1 9200 27570 9200 27570 7 FreeSans 2400 0 0 0 cell_unit_9/V_bias
flabel metal4 1950 29630 1950 29630 5 FreeSans 2400 0 0 0 cell_unit_9/OUT_P
flabel metal4 7210 29630 7210 29630 5 FreeSans 2400 0 0 0 cell_unit_9/OUT_N
flabel metal1 9200 21750 9200 21750 7 FreeSans 2400 0 0 0 cell_unit_9/GND
flabel metal2 4328 25992 4348 26120 7 FreeSans 300 180 0 0 cell_unit_9/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 25814 4348 25942 7 FreeSans 300 180 0 0 cell_unit_9/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 26158 4681 26224 0 FreeSans 300 0 0 0 cell_unit_9/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 25814 4412 25830 3 FreeSans 300 90 0 0 cell_unit_9/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 25710 4681 25776 0 FreeSans 300 0 0 0 cell_unit_9/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 25814 4806 25830 3 FreeSans 300 90 0 0 cell_unit_9/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 24210 18400 24210 7 FreeSans 2400 0 0 0 cell_unit_18/ON
flabel metal1 18400 27570 18400 27570 7 FreeSans 2400 0 0 0 cell_unit_18/V_bias
flabel metal4 11150 29630 11150 29630 5 FreeSans 2400 0 0 0 cell_unit_18/OUT_P
flabel metal4 16410 29630 16410 29630 5 FreeSans 2400 0 0 0 cell_unit_18/OUT_N
flabel metal1 18400 21750 18400 21750 7 FreeSans 2400 0 0 0 cell_unit_18/GND
flabel metal2 13528 25992 13548 26120 7 FreeSans 300 180 0 0 cell_unit_18/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 25814 13548 25942 7 FreeSans 300 180 0 0 cell_unit_18/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 26158 13881 26224 0 FreeSans 300 0 0 0 cell_unit_18/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 25814 13612 25830 3 FreeSans 300 90 0 0 cell_unit_18/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 25710 13881 25776 0 FreeSans 300 0 0 0 cell_unit_18/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 25814 14006 25830 3 FreeSans 300 90 0 0 cell_unit_18/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 24210 27600 24210 7 FreeSans 2400 0 0 0 cell_unit_19/ON
flabel metal1 27600 27570 27600 27570 7 FreeSans 2400 0 0 0 cell_unit_19/V_bias
flabel metal4 20350 29630 20350 29630 5 FreeSans 2400 0 0 0 cell_unit_19/OUT_P
flabel metal4 25610 29630 25610 29630 5 FreeSans 2400 0 0 0 cell_unit_19/OUT_N
flabel metal1 27600 21750 27600 21750 7 FreeSans 2400 0 0 0 cell_unit_19/GND
flabel metal2 22728 25992 22748 26120 7 FreeSans 300 180 0 0 cell_unit_19/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 25814 22748 25942 7 FreeSans 300 180 0 0 cell_unit_19/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 26158 23081 26224 0 FreeSans 300 0 0 0 cell_unit_19/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 25814 22812 25830 3 FreeSans 300 90 0 0 cell_unit_19/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 25710 23081 25776 0 FreeSans 300 0 0 0 cell_unit_19/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 25814 23206 25830 3 FreeSans 300 90 0 0 cell_unit_19/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 24210 36800 24210 7 FreeSans 2400 0 0 0 cell_unit_20/ON
flabel metal1 36800 27570 36800 27570 7 FreeSans 2400 0 0 0 cell_unit_20/V_bias
flabel metal4 29550 29630 29550 29630 5 FreeSans 2400 0 0 0 cell_unit_20/OUT_P
flabel metal4 34810 29630 34810 29630 5 FreeSans 2400 0 0 0 cell_unit_20/OUT_N
flabel metal1 36800 21750 36800 21750 7 FreeSans 2400 0 0 0 cell_unit_20/GND
flabel metal2 31928 25992 31948 26120 7 FreeSans 300 180 0 0 cell_unit_20/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 25814 31948 25942 7 FreeSans 300 180 0 0 cell_unit_20/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 26158 32281 26224 0 FreeSans 300 0 0 0 cell_unit_20/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 25814 32012 25830 3 FreeSans 300 90 0 0 cell_unit_20/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 25710 32281 25776 0 FreeSans 300 0 0 0 cell_unit_20/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 25814 32406 25830 3 FreeSans 300 90 0 0 cell_unit_20/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 24210 55200 24210 7 FreeSans 2400 0 0 0 cell_unit_22/ON
flabel metal1 55200 27570 55200 27570 7 FreeSans 2400 0 0 0 cell_unit_22/V_bias
flabel metal4 47950 29630 47950 29630 5 FreeSans 2400 0 0 0 cell_unit_22/OUT_P
flabel metal4 53210 29630 53210 29630 5 FreeSans 2400 0 0 0 cell_unit_22/OUT_N
flabel metal1 55200 21750 55200 21750 7 FreeSans 2400 0 0 0 cell_unit_22/GND
flabel metal2 50328 25992 50348 26120 7 FreeSans 300 180 0 0 cell_unit_22/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 25814 50348 25942 7 FreeSans 300 180 0 0 cell_unit_22/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 26158 50681 26224 0 FreeSans 300 0 0 0 cell_unit_22/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 25814 50412 25830 3 FreeSans 300 90 0 0 cell_unit_22/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 25710 50681 25776 0 FreeSans 300 0 0 0 cell_unit_22/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 25814 50806 25830 3 FreeSans 300 90 0 0 cell_unit_22/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 24210 46000 24210 7 FreeSans 2400 0 0 0 cell_unit_21/ON
flabel metal1 46000 27570 46000 27570 7 FreeSans 2400 0 0 0 cell_unit_21/V_bias
flabel metal4 38750 29630 38750 29630 5 FreeSans 2400 0 0 0 cell_unit_21/OUT_P
flabel metal4 44010 29630 44010 29630 5 FreeSans 2400 0 0 0 cell_unit_21/OUT_N
flabel metal1 46000 21750 46000 21750 7 FreeSans 2400 0 0 0 cell_unit_21/GND
flabel metal2 41128 25992 41148 26120 7 FreeSans 300 180 0 0 cell_unit_21/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 25814 41148 25942 7 FreeSans 300 180 0 0 cell_unit_21/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 26158 41481 26224 0 FreeSans 300 0 0 0 cell_unit_21/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 25814 41212 25830 3 FreeSans 300 90 0 0 cell_unit_21/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 25710 41481 25776 0 FreeSans 300 0 0 0 cell_unit_21/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 25814 41606 25830 3 FreeSans 300 90 0 0 cell_unit_21/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 24210 64400 24210 7 FreeSans 2400 0 0 0 cell_unit_23/ON
flabel metal1 64400 27570 64400 27570 7 FreeSans 2400 0 0 0 cell_unit_23/V_bias
flabel metal4 57150 29630 57150 29630 5 FreeSans 2400 0 0 0 cell_unit_23/OUT_P
flabel metal4 62410 29630 62410 29630 5 FreeSans 2400 0 0 0 cell_unit_23/OUT_N
flabel metal1 64400 21750 64400 21750 7 FreeSans 2400 0 0 0 cell_unit_23/GND
flabel metal2 59528 25992 59548 26120 7 FreeSans 300 180 0 0 cell_unit_23/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 25814 59548 25942 7 FreeSans 300 180 0 0 cell_unit_23/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 26158 59881 26224 0 FreeSans 300 0 0 0 cell_unit_23/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 25814 59612 25830 3 FreeSans 300 90 0 0 cell_unit_23/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 25710 59881 25776 0 FreeSans 300 0 0 0 cell_unit_23/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 25814 60006 25830 3 FreeSans 300 90 0 0 cell_unit_23/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 24210 73600 24210 7 FreeSans 2400 0 0 0 cell_unit_24/ON
flabel metal1 73600 27570 73600 27570 7 FreeSans 2400 0 0 0 cell_unit_24/V_bias
flabel metal4 66350 29630 66350 29630 5 FreeSans 2400 0 0 0 cell_unit_24/OUT_P
flabel metal4 71610 29630 71610 29630 5 FreeSans 2400 0 0 0 cell_unit_24/OUT_N
flabel metal1 73600 21750 73600 21750 7 FreeSans 2400 0 0 0 cell_unit_24/GND
flabel metal2 68728 25992 68748 26120 7 FreeSans 300 180 0 0 cell_unit_24/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 25814 68748 25942 7 FreeSans 300 180 0 0 cell_unit_24/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 26158 69081 26224 0 FreeSans 300 0 0 0 cell_unit_24/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 25814 68812 25830 3 FreeSans 300 90 0 0 cell_unit_24/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 25710 69081 25776 0 FreeSans 300 0 0 0 cell_unit_24/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 25814 69206 25830 3 FreeSans 300 90 0 0 cell_unit_24/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 9200 34090 9200 34090 7 FreeSans 2400 0 0 0 cell_unit_10/ON
flabel metal1 9200 37450 9200 37450 7 FreeSans 2400 0 0 0 cell_unit_10/V_bias
flabel metal4 1950 39510 1950 39510 5 FreeSans 2400 0 0 0 cell_unit_10/OUT_P
flabel metal4 7210 39510 7210 39510 5 FreeSans 2400 0 0 0 cell_unit_10/OUT_N
flabel metal1 9200 31630 9200 31630 7 FreeSans 2400 0 0 0 cell_unit_10/GND
flabel metal2 4328 35872 4348 36000 7 FreeSans 300 180 0 0 cell_unit_10/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 35694 4348 35822 7 FreeSans 300 180 0 0 cell_unit_10/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 36038 4681 36104 0 FreeSans 300 0 0 0 cell_unit_10/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 35694 4412 35710 3 FreeSans 300 90 0 0 cell_unit_10/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 35590 4681 35656 0 FreeSans 300 0 0 0 cell_unit_10/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 35694 4806 35710 3 FreeSans 300 90 0 0 cell_unit_10/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 34090 18400 34090 7 FreeSans 2400 0 0 0 cell_unit_25/ON
flabel metal1 18400 37450 18400 37450 7 FreeSans 2400 0 0 0 cell_unit_25/V_bias
flabel metal4 11150 39510 11150 39510 5 FreeSans 2400 0 0 0 cell_unit_25/OUT_P
flabel metal4 16410 39510 16410 39510 5 FreeSans 2400 0 0 0 cell_unit_25/OUT_N
flabel metal1 18400 31630 18400 31630 7 FreeSans 2400 0 0 0 cell_unit_25/GND
flabel metal2 13528 35872 13548 36000 7 FreeSans 300 180 0 0 cell_unit_25/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 35694 13548 35822 7 FreeSans 300 180 0 0 cell_unit_25/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 36038 13881 36104 0 FreeSans 300 0 0 0 cell_unit_25/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 35694 13612 35710 3 FreeSans 300 90 0 0 cell_unit_25/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 35590 13881 35656 0 FreeSans 300 0 0 0 cell_unit_25/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 35694 14006 35710 3 FreeSans 300 90 0 0 cell_unit_25/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 34090 27600 34090 7 FreeSans 2400 0 0 0 cell_unit_26/ON
flabel metal1 27600 37450 27600 37450 7 FreeSans 2400 0 0 0 cell_unit_26/V_bias
flabel metal4 20350 39510 20350 39510 5 FreeSans 2400 0 0 0 cell_unit_26/OUT_P
flabel metal4 25610 39510 25610 39510 5 FreeSans 2400 0 0 0 cell_unit_26/OUT_N
flabel metal1 27600 31630 27600 31630 7 FreeSans 2400 0 0 0 cell_unit_26/GND
flabel metal2 22728 35872 22748 36000 7 FreeSans 300 180 0 0 cell_unit_26/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 35694 22748 35822 7 FreeSans 300 180 0 0 cell_unit_26/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 36038 23081 36104 0 FreeSans 300 0 0 0 cell_unit_26/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 35694 22812 35710 3 FreeSans 300 90 0 0 cell_unit_26/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 35590 23081 35656 0 FreeSans 300 0 0 0 cell_unit_26/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 35694 23206 35710 3 FreeSans 300 90 0 0 cell_unit_26/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 34090 36800 34090 7 FreeSans 2400 0 0 0 cell_unit_27/ON
flabel metal1 36800 37450 36800 37450 7 FreeSans 2400 0 0 0 cell_unit_27/V_bias
flabel metal4 29550 39510 29550 39510 5 FreeSans 2400 0 0 0 cell_unit_27/OUT_P
flabel metal4 34810 39510 34810 39510 5 FreeSans 2400 0 0 0 cell_unit_27/OUT_N
flabel metal1 36800 31630 36800 31630 7 FreeSans 2400 0 0 0 cell_unit_27/GND
flabel metal2 31928 35872 31948 36000 7 FreeSans 300 180 0 0 cell_unit_27/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 35694 31948 35822 7 FreeSans 300 180 0 0 cell_unit_27/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 36038 32281 36104 0 FreeSans 300 0 0 0 cell_unit_27/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 35694 32012 35710 3 FreeSans 300 90 0 0 cell_unit_27/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 35590 32281 35656 0 FreeSans 300 0 0 0 cell_unit_27/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 35694 32406 35710 3 FreeSans 300 90 0 0 cell_unit_27/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 34090 55200 34090 7 FreeSans 2400 0 0 0 cell_unit_29/ON
flabel metal1 55200 37450 55200 37450 7 FreeSans 2400 0 0 0 cell_unit_29/V_bias
flabel metal4 47950 39510 47950 39510 5 FreeSans 2400 0 0 0 cell_unit_29/OUT_P
flabel metal4 53210 39510 53210 39510 5 FreeSans 2400 0 0 0 cell_unit_29/OUT_N
flabel metal1 55200 31630 55200 31630 7 FreeSans 2400 0 0 0 cell_unit_29/GND
flabel metal2 50328 35872 50348 36000 7 FreeSans 300 180 0 0 cell_unit_29/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 35694 50348 35822 7 FreeSans 300 180 0 0 cell_unit_29/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 36038 50681 36104 0 FreeSans 300 0 0 0 cell_unit_29/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 35694 50412 35710 3 FreeSans 300 90 0 0 cell_unit_29/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 35590 50681 35656 0 FreeSans 300 0 0 0 cell_unit_29/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 35694 50806 35710 3 FreeSans 300 90 0 0 cell_unit_29/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 34090 46000 34090 7 FreeSans 2400 0 0 0 cell_unit_28/ON
flabel metal1 46000 37450 46000 37450 7 FreeSans 2400 0 0 0 cell_unit_28/V_bias
flabel metal4 38750 39510 38750 39510 5 FreeSans 2400 0 0 0 cell_unit_28/OUT_P
flabel metal4 44010 39510 44010 39510 5 FreeSans 2400 0 0 0 cell_unit_28/OUT_N
flabel metal1 46000 31630 46000 31630 7 FreeSans 2400 0 0 0 cell_unit_28/GND
flabel metal2 41128 35872 41148 36000 7 FreeSans 300 180 0 0 cell_unit_28/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 35694 41148 35822 7 FreeSans 300 180 0 0 cell_unit_28/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 36038 41481 36104 0 FreeSans 300 0 0 0 cell_unit_28/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 35694 41212 35710 3 FreeSans 300 90 0 0 cell_unit_28/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 35590 41481 35656 0 FreeSans 300 0 0 0 cell_unit_28/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 35694 41606 35710 3 FreeSans 300 90 0 0 cell_unit_28/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 34090 64400 34090 7 FreeSans 2400 0 0 0 cell_unit_30/ON
flabel metal1 64400 37450 64400 37450 7 FreeSans 2400 0 0 0 cell_unit_30/V_bias
flabel metal4 57150 39510 57150 39510 5 FreeSans 2400 0 0 0 cell_unit_30/OUT_P
flabel metal4 62410 39510 62410 39510 5 FreeSans 2400 0 0 0 cell_unit_30/OUT_N
flabel metal1 64400 31630 64400 31630 7 FreeSans 2400 0 0 0 cell_unit_30/GND
flabel metal2 59528 35872 59548 36000 7 FreeSans 300 180 0 0 cell_unit_30/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 35694 59548 35822 7 FreeSans 300 180 0 0 cell_unit_30/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 36038 59881 36104 0 FreeSans 300 0 0 0 cell_unit_30/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 35694 59612 35710 3 FreeSans 300 90 0 0 cell_unit_30/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 35590 59881 35656 0 FreeSans 300 0 0 0 cell_unit_30/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 35694 60006 35710 3 FreeSans 300 90 0 0 cell_unit_30/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 34090 73600 34090 7 FreeSans 2400 0 0 0 cell_unit_31/ON
flabel metal1 73600 37450 73600 37450 7 FreeSans 2400 0 0 0 cell_unit_31/V_bias
flabel metal4 66350 39510 66350 39510 5 FreeSans 2400 0 0 0 cell_unit_31/OUT_P
flabel metal4 71610 39510 71610 39510 5 FreeSans 2400 0 0 0 cell_unit_31/OUT_N
flabel metal1 73600 31630 73600 31630 7 FreeSans 2400 0 0 0 cell_unit_31/GND
flabel metal2 68728 35872 68748 36000 7 FreeSans 300 180 0 0 cell_unit_31/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 35694 68748 35822 7 FreeSans 300 180 0 0 cell_unit_31/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 36038 69081 36104 0 FreeSans 300 0 0 0 cell_unit_31/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 35694 68812 35710 3 FreeSans 300 90 0 0 cell_unit_31/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 35590 69081 35656 0 FreeSans 300 0 0 0 cell_unit_31/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 35694 69206 35710 3 FreeSans 300 90 0 0 cell_unit_31/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 -610 45410 -610 45410 1 FreeSans 400 0 0 0 inv_1_1/OUT
flabel metal2 -110 45360 -110 45360 1 FreeSans 400 0 0 0 inv_1_1/ON
flabel metal2 -5820 49390 -5820 49390 5 FreeSans 2400 0 0 0 inv_1_1/VDD
flabel metal1 -2820 49390 -2820 49390 5 FreeSans 2400 0 0 0 inv_1_1/GND
flabel metal2 9200 43970 9200 43970 7 FreeSans 2400 0 0 0 cell_unit_32/ON
flabel metal1 9200 47330 9200 47330 7 FreeSans 2400 0 0 0 cell_unit_32/V_bias
flabel metal4 1950 49390 1950 49390 5 FreeSans 2400 0 0 0 cell_unit_32/OUT_P
flabel metal4 7210 49390 7210 49390 5 FreeSans 2400 0 0 0 cell_unit_32/OUT_N
flabel metal1 9200 41510 9200 41510 7 FreeSans 2400 0 0 0 cell_unit_32/GND
flabel metal2 4328 45752 4348 45880 7 FreeSans 300 180 0 0 cell_unit_32/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 45574 4348 45702 7 FreeSans 300 180 0 0 cell_unit_32/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 45918 4681 45984 0 FreeSans 300 0 0 0 cell_unit_32/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 45574 4412 45590 3 FreeSans 300 90 0 0 cell_unit_32/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 45470 4681 45536 0 FreeSans 300 0 0 0 cell_unit_32/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 45574 4806 45590 3 FreeSans 300 90 0 0 cell_unit_32/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 43970 18400 43970 7 FreeSans 2400 0 0 0 cell_unit_34/ON
flabel metal1 18400 47330 18400 47330 7 FreeSans 2400 0 0 0 cell_unit_34/V_bias
flabel metal4 11150 49390 11150 49390 5 FreeSans 2400 0 0 0 cell_unit_34/OUT_P
flabel metal4 16410 49390 16410 49390 5 FreeSans 2400 0 0 0 cell_unit_34/OUT_N
flabel metal1 18400 41510 18400 41510 7 FreeSans 2400 0 0 0 cell_unit_34/GND
flabel metal2 13528 45752 13548 45880 7 FreeSans 300 180 0 0 cell_unit_34/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 45574 13548 45702 7 FreeSans 300 180 0 0 cell_unit_34/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 45918 13881 45984 0 FreeSans 300 0 0 0 cell_unit_34/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 45574 13612 45590 3 FreeSans 300 90 0 0 cell_unit_34/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 45470 13881 45536 0 FreeSans 300 0 0 0 cell_unit_34/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 45574 14006 45590 3 FreeSans 300 90 0 0 cell_unit_34/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 43970 27600 43970 7 FreeSans 2400 0 0 0 cell_unit_35/ON
flabel metal1 27600 47330 27600 47330 7 FreeSans 2400 0 0 0 cell_unit_35/V_bias
flabel metal4 20350 49390 20350 49390 5 FreeSans 2400 0 0 0 cell_unit_35/OUT_P
flabel metal4 25610 49390 25610 49390 5 FreeSans 2400 0 0 0 cell_unit_35/OUT_N
flabel metal1 27600 41510 27600 41510 7 FreeSans 2400 0 0 0 cell_unit_35/GND
flabel metal2 22728 45752 22748 45880 7 FreeSans 300 180 0 0 cell_unit_35/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 45574 22748 45702 7 FreeSans 300 180 0 0 cell_unit_35/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 45918 23081 45984 0 FreeSans 300 0 0 0 cell_unit_35/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 45574 22812 45590 3 FreeSans 300 90 0 0 cell_unit_35/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 45470 23081 45536 0 FreeSans 300 0 0 0 cell_unit_35/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 45574 23206 45590 3 FreeSans 300 90 0 0 cell_unit_35/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 43970 36800 43970 7 FreeSans 2400 0 0 0 cell_unit_36/ON
flabel metal1 36800 47330 36800 47330 7 FreeSans 2400 0 0 0 cell_unit_36/V_bias
flabel metal4 29550 49390 29550 49390 5 FreeSans 2400 0 0 0 cell_unit_36/OUT_P
flabel metal4 34810 49390 34810 49390 5 FreeSans 2400 0 0 0 cell_unit_36/OUT_N
flabel metal1 36800 41510 36800 41510 7 FreeSans 2400 0 0 0 cell_unit_36/GND
flabel metal2 31928 45752 31948 45880 7 FreeSans 300 180 0 0 cell_unit_36/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 45574 31948 45702 7 FreeSans 300 180 0 0 cell_unit_36/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 45918 32281 45984 0 FreeSans 300 0 0 0 cell_unit_36/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 45574 32012 45590 3 FreeSans 300 90 0 0 cell_unit_36/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 45470 32281 45536 0 FreeSans 300 0 0 0 cell_unit_36/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 45574 32406 45590 3 FreeSans 300 90 0 0 cell_unit_36/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 43970 55200 43970 7 FreeSans 2400 0 0 0 cell_unit_38/ON
flabel metal1 55200 47330 55200 47330 7 FreeSans 2400 0 0 0 cell_unit_38/V_bias
flabel metal4 47950 49390 47950 49390 5 FreeSans 2400 0 0 0 cell_unit_38/OUT_P
flabel metal4 53210 49390 53210 49390 5 FreeSans 2400 0 0 0 cell_unit_38/OUT_N
flabel metal1 55200 41510 55200 41510 7 FreeSans 2400 0 0 0 cell_unit_38/GND
flabel metal2 50328 45752 50348 45880 7 FreeSans 300 180 0 0 cell_unit_38/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 45574 50348 45702 7 FreeSans 300 180 0 0 cell_unit_38/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 45918 50681 45984 0 FreeSans 300 0 0 0 cell_unit_38/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 45574 50412 45590 3 FreeSans 300 90 0 0 cell_unit_38/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 45470 50681 45536 0 FreeSans 300 0 0 0 cell_unit_38/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 45574 50806 45590 3 FreeSans 300 90 0 0 cell_unit_38/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 43970 46000 43970 7 FreeSans 2400 0 0 0 cell_unit_37/ON
flabel metal1 46000 47330 46000 47330 7 FreeSans 2400 0 0 0 cell_unit_37/V_bias
flabel metal4 38750 49390 38750 49390 5 FreeSans 2400 0 0 0 cell_unit_37/OUT_P
flabel metal4 44010 49390 44010 49390 5 FreeSans 2400 0 0 0 cell_unit_37/OUT_N
flabel metal1 46000 41510 46000 41510 7 FreeSans 2400 0 0 0 cell_unit_37/GND
flabel metal2 41128 45752 41148 45880 7 FreeSans 300 180 0 0 cell_unit_37/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 45574 41148 45702 7 FreeSans 300 180 0 0 cell_unit_37/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 45918 41481 45984 0 FreeSans 300 0 0 0 cell_unit_37/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 45574 41212 45590 3 FreeSans 300 90 0 0 cell_unit_37/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 45470 41481 45536 0 FreeSans 300 0 0 0 cell_unit_37/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 45574 41606 45590 3 FreeSans 300 90 0 0 cell_unit_37/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 43970 64400 43970 7 FreeSans 2400 0 0 0 cell_unit_39/ON
flabel metal1 64400 47330 64400 47330 7 FreeSans 2400 0 0 0 cell_unit_39/V_bias
flabel metal4 57150 49390 57150 49390 5 FreeSans 2400 0 0 0 cell_unit_39/OUT_P
flabel metal4 62410 49390 62410 49390 5 FreeSans 2400 0 0 0 cell_unit_39/OUT_N
flabel metal1 64400 41510 64400 41510 7 FreeSans 2400 0 0 0 cell_unit_39/GND
flabel metal2 59528 45752 59548 45880 7 FreeSans 300 180 0 0 cell_unit_39/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 45574 59548 45702 7 FreeSans 300 180 0 0 cell_unit_39/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 45918 59881 45984 0 FreeSans 300 0 0 0 cell_unit_39/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 45574 59612 45590 3 FreeSans 300 90 0 0 cell_unit_39/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 45470 59881 45536 0 FreeSans 300 0 0 0 cell_unit_39/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 45574 60006 45590 3 FreeSans 300 90 0 0 cell_unit_39/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 43970 73600 43970 7 FreeSans 2400 0 0 0 cell_unit_40/ON
flabel metal1 73600 47330 73600 47330 7 FreeSans 2400 0 0 0 cell_unit_40/V_bias
flabel metal4 66350 49390 66350 49390 5 FreeSans 2400 0 0 0 cell_unit_40/OUT_P
flabel metal4 71610 49390 71610 49390 5 FreeSans 2400 0 0 0 cell_unit_40/OUT_N
flabel metal1 73600 41510 73600 41510 7 FreeSans 2400 0 0 0 cell_unit_40/GND
flabel metal2 68728 45752 68748 45880 7 FreeSans 300 180 0 0 cell_unit_40/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 45574 68748 45702 7 FreeSans 300 180 0 0 cell_unit_40/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 45918 69081 45984 0 FreeSans 300 0 0 0 cell_unit_40/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 45574 68812 45590 3 FreeSans 300 90 0 0 cell_unit_40/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 45470 69081 45536 0 FreeSans 300 0 0 0 cell_unit_40/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 45574 69206 45590 3 FreeSans 300 90 0 0 cell_unit_40/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 9200 53850 9200 53850 7 FreeSans 2400 0 0 0 cell_unit_33/ON
flabel metal1 9200 57210 9200 57210 7 FreeSans 2400 0 0 0 cell_unit_33/V_bias
flabel metal4 1950 59270 1950 59270 5 FreeSans 2400 0 0 0 cell_unit_33/OUT_P
flabel metal4 7210 59270 7210 59270 5 FreeSans 2400 0 0 0 cell_unit_33/OUT_N
flabel metal1 9200 51390 9200 51390 7 FreeSans 2400 0 0 0 cell_unit_33/GND
flabel metal2 4328 55632 4348 55760 7 FreeSans 300 180 0 0 cell_unit_33/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 55454 4348 55582 7 FreeSans 300 180 0 0 cell_unit_33/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 55798 4681 55864 0 FreeSans 300 0 0 0 cell_unit_33/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 55454 4412 55470 3 FreeSans 300 90 0 0 cell_unit_33/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 55350 4681 55416 0 FreeSans 300 0 0 0 cell_unit_33/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 55454 4806 55470 3 FreeSans 300 90 0 0 cell_unit_33/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 53850 18400 53850 7 FreeSans 2400 0 0 0 cell_unit_41/ON
flabel metal1 18400 57210 18400 57210 7 FreeSans 2400 0 0 0 cell_unit_41/V_bias
flabel metal4 11150 59270 11150 59270 5 FreeSans 2400 0 0 0 cell_unit_41/OUT_P
flabel metal4 16410 59270 16410 59270 5 FreeSans 2400 0 0 0 cell_unit_41/OUT_N
flabel metal1 18400 51390 18400 51390 7 FreeSans 2400 0 0 0 cell_unit_41/GND
flabel metal2 13528 55632 13548 55760 7 FreeSans 300 180 0 0 cell_unit_41/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 55454 13548 55582 7 FreeSans 300 180 0 0 cell_unit_41/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 55798 13881 55864 0 FreeSans 300 0 0 0 cell_unit_41/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 55454 13612 55470 3 FreeSans 300 90 0 0 cell_unit_41/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 55350 13881 55416 0 FreeSans 300 0 0 0 cell_unit_41/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 55454 14006 55470 3 FreeSans 300 90 0 0 cell_unit_41/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 53850 27600 53850 7 FreeSans 2400 0 0 0 cell_unit_42/ON
flabel metal1 27600 57210 27600 57210 7 FreeSans 2400 0 0 0 cell_unit_42/V_bias
flabel metal4 20350 59270 20350 59270 5 FreeSans 2400 0 0 0 cell_unit_42/OUT_P
flabel metal4 25610 59270 25610 59270 5 FreeSans 2400 0 0 0 cell_unit_42/OUT_N
flabel metal1 27600 51390 27600 51390 7 FreeSans 2400 0 0 0 cell_unit_42/GND
flabel metal2 22728 55632 22748 55760 7 FreeSans 300 180 0 0 cell_unit_42/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 55454 22748 55582 7 FreeSans 300 180 0 0 cell_unit_42/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 55798 23081 55864 0 FreeSans 300 0 0 0 cell_unit_42/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 55454 22812 55470 3 FreeSans 300 90 0 0 cell_unit_42/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 55350 23081 55416 0 FreeSans 300 0 0 0 cell_unit_42/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 55454 23206 55470 3 FreeSans 300 90 0 0 cell_unit_42/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 53850 36800 53850 7 FreeSans 2400 0 0 0 cell_unit_43/ON
flabel metal1 36800 57210 36800 57210 7 FreeSans 2400 0 0 0 cell_unit_43/V_bias
flabel metal4 29550 59270 29550 59270 5 FreeSans 2400 0 0 0 cell_unit_43/OUT_P
flabel metal4 34810 59270 34810 59270 5 FreeSans 2400 0 0 0 cell_unit_43/OUT_N
flabel metal1 36800 51390 36800 51390 7 FreeSans 2400 0 0 0 cell_unit_43/GND
flabel metal2 31928 55632 31948 55760 7 FreeSans 300 180 0 0 cell_unit_43/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 55454 31948 55582 7 FreeSans 300 180 0 0 cell_unit_43/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 55798 32281 55864 0 FreeSans 300 0 0 0 cell_unit_43/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 55454 32012 55470 3 FreeSans 300 90 0 0 cell_unit_43/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 55350 32281 55416 0 FreeSans 300 0 0 0 cell_unit_43/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 55454 32406 55470 3 FreeSans 300 90 0 0 cell_unit_43/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 53850 55200 53850 7 FreeSans 2400 0 0 0 cell_unit_45/ON
flabel metal1 55200 57210 55200 57210 7 FreeSans 2400 0 0 0 cell_unit_45/V_bias
flabel metal4 47950 59270 47950 59270 5 FreeSans 2400 0 0 0 cell_unit_45/OUT_P
flabel metal4 53210 59270 53210 59270 5 FreeSans 2400 0 0 0 cell_unit_45/OUT_N
flabel metal1 55200 51390 55200 51390 7 FreeSans 2400 0 0 0 cell_unit_45/GND
flabel metal2 50328 55632 50348 55760 7 FreeSans 300 180 0 0 cell_unit_45/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 55454 50348 55582 7 FreeSans 300 180 0 0 cell_unit_45/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 55798 50681 55864 0 FreeSans 300 0 0 0 cell_unit_45/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 55454 50412 55470 3 FreeSans 300 90 0 0 cell_unit_45/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 55350 50681 55416 0 FreeSans 300 0 0 0 cell_unit_45/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 55454 50806 55470 3 FreeSans 300 90 0 0 cell_unit_45/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 53850 46000 53850 7 FreeSans 2400 0 0 0 cell_unit_44/ON
flabel metal1 46000 57210 46000 57210 7 FreeSans 2400 0 0 0 cell_unit_44/V_bias
flabel metal4 38750 59270 38750 59270 5 FreeSans 2400 0 0 0 cell_unit_44/OUT_P
flabel metal4 44010 59270 44010 59270 5 FreeSans 2400 0 0 0 cell_unit_44/OUT_N
flabel metal1 46000 51390 46000 51390 7 FreeSans 2400 0 0 0 cell_unit_44/GND
flabel metal2 41128 55632 41148 55760 7 FreeSans 300 180 0 0 cell_unit_44/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 55454 41148 55582 7 FreeSans 300 180 0 0 cell_unit_44/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 55798 41481 55864 0 FreeSans 300 0 0 0 cell_unit_44/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 55454 41212 55470 3 FreeSans 300 90 0 0 cell_unit_44/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 55350 41481 55416 0 FreeSans 300 0 0 0 cell_unit_44/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 55454 41606 55470 3 FreeSans 300 90 0 0 cell_unit_44/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 53850 64400 53850 7 FreeSans 2400 0 0 0 cell_unit_46/ON
flabel metal1 64400 57210 64400 57210 7 FreeSans 2400 0 0 0 cell_unit_46/V_bias
flabel metal4 57150 59270 57150 59270 5 FreeSans 2400 0 0 0 cell_unit_46/OUT_P
flabel metal4 62410 59270 62410 59270 5 FreeSans 2400 0 0 0 cell_unit_46/OUT_N
flabel metal1 64400 51390 64400 51390 7 FreeSans 2400 0 0 0 cell_unit_46/GND
flabel metal2 59528 55632 59548 55760 7 FreeSans 300 180 0 0 cell_unit_46/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 55454 59548 55582 7 FreeSans 300 180 0 0 cell_unit_46/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 55798 59881 55864 0 FreeSans 300 0 0 0 cell_unit_46/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 55454 59612 55470 3 FreeSans 300 90 0 0 cell_unit_46/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 55350 59881 55416 0 FreeSans 300 0 0 0 cell_unit_46/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 55454 60006 55470 3 FreeSans 300 90 0 0 cell_unit_46/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 53850 73600 53850 7 FreeSans 2400 0 0 0 cell_unit_47/ON
flabel metal1 73600 57210 73600 57210 7 FreeSans 2400 0 0 0 cell_unit_47/V_bias
flabel metal4 66350 59270 66350 59270 5 FreeSans 2400 0 0 0 cell_unit_47/OUT_P
flabel metal4 71610 59270 71610 59270 5 FreeSans 2400 0 0 0 cell_unit_47/OUT_N
flabel metal1 73600 51390 73600 51390 7 FreeSans 2400 0 0 0 cell_unit_47/GND
flabel metal2 68728 55632 68748 55760 7 FreeSans 300 180 0 0 cell_unit_47/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 55454 68748 55582 7 FreeSans 300 180 0 0 cell_unit_47/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 55798 69081 55864 0 FreeSans 300 0 0 0 cell_unit_47/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 55454 68812 55470 3 FreeSans 300 90 0 0 cell_unit_47/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 55350 69081 55416 0 FreeSans 300 0 0 0 cell_unit_47/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 55454 69206 55470 3 FreeSans 300 90 0 0 cell_unit_47/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 -610 65170 -610 65170 1 FreeSans 400 0 0 0 inv_1_2/OUT
flabel metal2 -110 65120 -110 65120 1 FreeSans 400 0 0 0 inv_1_2/ON
flabel metal2 -5820 69150 -5820 69150 5 FreeSans 2400 0 0 0 inv_1_2/VDD
flabel metal1 -2820 69150 -2820 69150 5 FreeSans 2400 0 0 0 inv_1_2/GND
flabel metal2 9200 63730 9200 63730 7 FreeSans 2400 0 0 0 cell_unit_48/ON
flabel metal1 9200 67090 9200 67090 7 FreeSans 2400 0 0 0 cell_unit_48/V_bias
flabel metal4 1950 69150 1950 69150 5 FreeSans 2400 0 0 0 cell_unit_48/OUT_P
flabel metal4 7210 69150 7210 69150 5 FreeSans 2400 0 0 0 cell_unit_48/OUT_N
flabel metal1 9200 61270 9200 61270 7 FreeSans 2400 0 0 0 cell_unit_48/GND
flabel metal2 4328 65512 4348 65640 7 FreeSans 300 180 0 0 cell_unit_48/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 65334 4348 65462 7 FreeSans 300 180 0 0 cell_unit_48/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 65678 4681 65744 0 FreeSans 300 0 0 0 cell_unit_48/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 65334 4412 65350 3 FreeSans 300 90 0 0 cell_unit_48/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 65230 4681 65296 0 FreeSans 300 0 0 0 cell_unit_48/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 65334 4806 65350 3 FreeSans 300 90 0 0 cell_unit_48/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 63730 18400 63730 7 FreeSans 2400 0 0 0 cell_unit_49/ON
flabel metal1 18400 67090 18400 67090 7 FreeSans 2400 0 0 0 cell_unit_49/V_bias
flabel metal4 11150 69150 11150 69150 5 FreeSans 2400 0 0 0 cell_unit_49/OUT_P
flabel metal4 16410 69150 16410 69150 5 FreeSans 2400 0 0 0 cell_unit_49/OUT_N
flabel metal1 18400 61270 18400 61270 7 FreeSans 2400 0 0 0 cell_unit_49/GND
flabel metal2 13528 65512 13548 65640 7 FreeSans 300 180 0 0 cell_unit_49/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 65334 13548 65462 7 FreeSans 300 180 0 0 cell_unit_49/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 65678 13881 65744 0 FreeSans 300 0 0 0 cell_unit_49/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 65334 13612 65350 3 FreeSans 300 90 0 0 cell_unit_49/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 65230 13881 65296 0 FreeSans 300 0 0 0 cell_unit_49/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 65334 14006 65350 3 FreeSans 300 90 0 0 cell_unit_49/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 63730 27600 63730 7 FreeSans 2400 0 0 0 cell_unit_50/ON
flabel metal1 27600 67090 27600 67090 7 FreeSans 2400 0 0 0 cell_unit_50/V_bias
flabel metal4 20350 69150 20350 69150 5 FreeSans 2400 0 0 0 cell_unit_50/OUT_P
flabel metal4 25610 69150 25610 69150 5 FreeSans 2400 0 0 0 cell_unit_50/OUT_N
flabel metal1 27600 61270 27600 61270 7 FreeSans 2400 0 0 0 cell_unit_50/GND
flabel metal2 22728 65512 22748 65640 7 FreeSans 300 180 0 0 cell_unit_50/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 65334 22748 65462 7 FreeSans 300 180 0 0 cell_unit_50/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 65678 23081 65744 0 FreeSans 300 0 0 0 cell_unit_50/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 65334 22812 65350 3 FreeSans 300 90 0 0 cell_unit_50/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 65230 23081 65296 0 FreeSans 300 0 0 0 cell_unit_50/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 65334 23206 65350 3 FreeSans 300 90 0 0 cell_unit_50/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 63730 36800 63730 7 FreeSans 2400 0 0 0 cell_unit_51/ON
flabel metal1 36800 67090 36800 67090 7 FreeSans 2400 0 0 0 cell_unit_51/V_bias
flabel metal4 29550 69150 29550 69150 5 FreeSans 2400 0 0 0 cell_unit_51/OUT_P
flabel metal4 34810 69150 34810 69150 5 FreeSans 2400 0 0 0 cell_unit_51/OUT_N
flabel metal1 36800 61270 36800 61270 7 FreeSans 2400 0 0 0 cell_unit_51/GND
flabel metal2 31928 65512 31948 65640 7 FreeSans 300 180 0 0 cell_unit_51/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 65334 31948 65462 7 FreeSans 300 180 0 0 cell_unit_51/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 65678 32281 65744 0 FreeSans 300 0 0 0 cell_unit_51/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 65334 32012 65350 3 FreeSans 300 90 0 0 cell_unit_51/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 65230 32281 65296 0 FreeSans 300 0 0 0 cell_unit_51/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 65334 32406 65350 3 FreeSans 300 90 0 0 cell_unit_51/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 55200 63730 55200 63730 7 FreeSans 2400 0 0 0 cell_unit_53/ON
flabel metal1 55200 67090 55200 67090 7 FreeSans 2400 0 0 0 cell_unit_53/V_bias
flabel metal4 47950 69150 47950 69150 5 FreeSans 2400 0 0 0 cell_unit_53/OUT_P
flabel metal4 53210 69150 53210 69150 5 FreeSans 2400 0 0 0 cell_unit_53/OUT_N
flabel metal1 55200 61270 55200 61270 7 FreeSans 2400 0 0 0 cell_unit_53/GND
flabel metal2 50328 65512 50348 65640 7 FreeSans 300 180 0 0 cell_unit_53/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 50328 65334 50348 65462 7 FreeSans 300 180 0 0 cell_unit_53/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 50479 65678 50681 65744 0 FreeSans 300 0 0 0 cell_unit_53/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50354 65334 50412 65350 3 FreeSans 300 90 0 0 cell_unit_53/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 50479 65230 50681 65296 0 FreeSans 300 0 0 0 cell_unit_53/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 50748 65334 50806 65350 3 FreeSans 300 90 0 0 cell_unit_53/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 46000 63730 46000 63730 7 FreeSans 2400 0 0 0 cell_unit_52/ON
flabel metal1 46000 67090 46000 67090 7 FreeSans 2400 0 0 0 cell_unit_52/V_bias
flabel metal4 38750 69150 38750 69150 5 FreeSans 2400 0 0 0 cell_unit_52/OUT_P
flabel metal4 44010 69150 44010 69150 5 FreeSans 2400 0 0 0 cell_unit_52/OUT_N
flabel metal1 46000 61270 46000 61270 7 FreeSans 2400 0 0 0 cell_unit_52/GND
flabel metal2 41128 65512 41148 65640 7 FreeSans 300 180 0 0 cell_unit_52/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 41128 65334 41148 65462 7 FreeSans 300 180 0 0 cell_unit_52/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 41279 65678 41481 65744 0 FreeSans 300 0 0 0 cell_unit_52/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41154 65334 41212 65350 3 FreeSans 300 90 0 0 cell_unit_52/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 41279 65230 41481 65296 0 FreeSans 300 0 0 0 cell_unit_52/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 41548 65334 41606 65350 3 FreeSans 300 90 0 0 cell_unit_52/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 64400 63730 64400 63730 7 FreeSans 2400 0 0 0 cell_unit_54/ON
flabel metal1 64400 67090 64400 67090 7 FreeSans 2400 0 0 0 cell_unit_54/V_bias
flabel metal4 57150 69150 57150 69150 5 FreeSans 2400 0 0 0 cell_unit_54/OUT_P
flabel metal4 62410 69150 62410 69150 5 FreeSans 2400 0 0 0 cell_unit_54/OUT_N
flabel metal1 64400 61270 64400 61270 7 FreeSans 2400 0 0 0 cell_unit_54/GND
flabel metal2 59528 65512 59548 65640 7 FreeSans 300 180 0 0 cell_unit_54/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 59528 65334 59548 65462 7 FreeSans 300 180 0 0 cell_unit_54/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 59679 65678 59881 65744 0 FreeSans 300 0 0 0 cell_unit_54/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59554 65334 59612 65350 3 FreeSans 300 90 0 0 cell_unit_54/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 59679 65230 59881 65296 0 FreeSans 300 0 0 0 cell_unit_54/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 59948 65334 60006 65350 3 FreeSans 300 90 0 0 cell_unit_54/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 73600 63730 73600 63730 7 FreeSans 2400 0 0 0 cell_unit_55/ON
flabel metal1 73600 67090 73600 67090 7 FreeSans 2400 0 0 0 cell_unit_55/V_bias
flabel metal4 66350 69150 66350 69150 5 FreeSans 2400 0 0 0 cell_unit_55/OUT_P
flabel metal4 71610 69150 71610 69150 5 FreeSans 2400 0 0 0 cell_unit_55/OUT_N
flabel metal1 73600 61270 73600 61270 7 FreeSans 2400 0 0 0 cell_unit_55/GND
flabel metal2 68728 65512 68748 65640 7 FreeSans 300 180 0 0 cell_unit_55/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 68728 65334 68748 65462 7 FreeSans 300 180 0 0 cell_unit_55/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 68879 65678 69081 65744 0 FreeSans 300 0 0 0 cell_unit_55/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 68754 65334 68812 65350 3 FreeSans 300 90 0 0 cell_unit_55/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 68879 65230 69081 65296 0 FreeSans 300 0 0 0 cell_unit_55/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 69148 65334 69206 65350 3 FreeSans 300 90 0 0 cell_unit_55/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 -610 75050 -610 75050 1 FreeSans 400 0 0 0 inv_1_3/OUT
flabel metal2 -110 75000 -110 75000 1 FreeSans 400 0 0 0 inv_1_3/ON
flabel metal2 -5820 79030 -5820 79030 5 FreeSans 2400 0 0 0 inv_1_3/VDD
flabel metal1 -2820 79030 -2820 79030 5 FreeSans 2400 0 0 0 inv_1_3/GND
flabel metal2 9200 73610 9200 73610 7 FreeSans 2400 0 0 0 cell_unit_56/ON
flabel metal1 9200 76970 9200 76970 7 FreeSans 2400 0 0 0 cell_unit_56/V_bias
flabel metal4 1950 79030 1950 79030 5 FreeSans 2400 0 0 0 cell_unit_56/OUT_P
flabel metal4 7210 79030 7210 79030 5 FreeSans 2400 0 0 0 cell_unit_56/OUT_N
flabel metal1 9200 71150 9200 71150 7 FreeSans 2400 0 0 0 cell_unit_56/GND
flabel metal2 4328 75392 4348 75520 7 FreeSans 300 180 0 0 cell_unit_56/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 75214 4348 75342 7 FreeSans 300 180 0 0 cell_unit_56/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 75558 4681 75624 0 FreeSans 300 0 0 0 cell_unit_56/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 75214 4412 75230 3 FreeSans 300 90 0 0 cell_unit_56/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 75110 4681 75176 0 FreeSans 300 0 0 0 cell_unit_56/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 75214 4806 75230 3 FreeSans 300 90 0 0 cell_unit_56/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 73610 18400 73610 7 FreeSans 2400 0 0 0 cell_unit_57/ON
flabel metal1 18400 76970 18400 76970 7 FreeSans 2400 0 0 0 cell_unit_57/V_bias
flabel metal4 11150 79030 11150 79030 5 FreeSans 2400 0 0 0 cell_unit_57/OUT_P
flabel metal4 16410 79030 16410 79030 5 FreeSans 2400 0 0 0 cell_unit_57/OUT_N
flabel metal1 18400 71150 18400 71150 7 FreeSans 2400 0 0 0 cell_unit_57/GND
flabel metal2 13528 75392 13548 75520 7 FreeSans 300 180 0 0 cell_unit_57/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 75214 13548 75342 7 FreeSans 300 180 0 0 cell_unit_57/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 75558 13881 75624 0 FreeSans 300 0 0 0 cell_unit_57/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 75214 13612 75230 3 FreeSans 300 90 0 0 cell_unit_57/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 75110 13881 75176 0 FreeSans 300 0 0 0 cell_unit_57/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 75214 14006 75230 3 FreeSans 300 90 0 0 cell_unit_57/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 27600 73610 27600 73610 7 FreeSans 2400 0 0 0 cell_unit_58/ON
flabel metal1 27600 76970 27600 76970 7 FreeSans 2400 0 0 0 cell_unit_58/V_bias
flabel metal4 20350 79030 20350 79030 5 FreeSans 2400 0 0 0 cell_unit_58/OUT_P
flabel metal4 25610 79030 25610 79030 5 FreeSans 2400 0 0 0 cell_unit_58/OUT_N
flabel metal1 27600 71150 27600 71150 7 FreeSans 2400 0 0 0 cell_unit_58/GND
flabel metal2 22728 75392 22748 75520 7 FreeSans 300 180 0 0 cell_unit_58/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 22728 75214 22748 75342 7 FreeSans 300 180 0 0 cell_unit_58/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 22879 75558 23081 75624 0 FreeSans 300 0 0 0 cell_unit_58/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 22754 75214 22812 75230 3 FreeSans 300 90 0 0 cell_unit_58/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 22879 75110 23081 75176 0 FreeSans 300 0 0 0 cell_unit_58/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 23148 75214 23206 75230 3 FreeSans 300 90 0 0 cell_unit_58/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 36800 73610 36800 73610 7 FreeSans 2400 0 0 0 cell_unit_59/ON
flabel metal1 36800 76970 36800 76970 7 FreeSans 2400 0 0 0 cell_unit_59/V_bias
flabel metal4 29550 79030 29550 79030 5 FreeSans 2400 0 0 0 cell_unit_59/OUT_P
flabel metal4 34810 79030 34810 79030 5 FreeSans 2400 0 0 0 cell_unit_59/OUT_N
flabel metal1 36800 71150 36800 71150 7 FreeSans 2400 0 0 0 cell_unit_59/GND
flabel metal2 31928 75392 31948 75520 7 FreeSans 300 180 0 0 cell_unit_59/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 31928 75214 31948 75342 7 FreeSans 300 180 0 0 cell_unit_59/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 32079 75558 32281 75624 0 FreeSans 300 0 0 0 cell_unit_59/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 31954 75214 32012 75230 3 FreeSans 300 90 0 0 cell_unit_59/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 32079 75110 32281 75176 0 FreeSans 300 0 0 0 cell_unit_59/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 32348 75214 32406 75230 3 FreeSans 300 90 0 0 cell_unit_59/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 -610 84930 -610 84930 1 FreeSans 400 0 0 0 inv_1_4/OUT
flabel metal2 -110 84880 -110 84880 1 FreeSans 400 0 0 0 inv_1_4/ON
flabel metal2 -5820 88910 -5820 88910 5 FreeSans 2400 0 0 0 inv_1_4/VDD
flabel metal1 -2820 88910 -2820 88910 5 FreeSans 2400 0 0 0 inv_1_4/GND
flabel metal2 9200 83490 9200 83490 7 FreeSans 2400 0 0 0 cell_unit_60/ON
flabel metal1 9200 86850 9200 86850 7 FreeSans 2400 0 0 0 cell_unit_60/V_bias
flabel metal4 1950 88910 1950 88910 5 FreeSans 2400 0 0 0 cell_unit_60/OUT_P
flabel metal4 7210 88910 7210 88910 5 FreeSans 2400 0 0 0 cell_unit_60/OUT_N
flabel metal1 9200 81030 9200 81030 7 FreeSans 2400 0 0 0 cell_unit_60/GND
flabel metal2 4328 85272 4348 85400 7 FreeSans 300 180 0 0 cell_unit_60/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 85094 4348 85222 7 FreeSans 300 180 0 0 cell_unit_60/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 85438 4681 85504 0 FreeSans 300 0 0 0 cell_unit_60/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 85094 4412 85110 3 FreeSans 300 90 0 0 cell_unit_60/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 84990 4681 85056 0 FreeSans 300 0 0 0 cell_unit_60/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 85094 4806 85110 3 FreeSans 300 90 0 0 cell_unit_60/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal2 18400 83490 18400 83490 7 FreeSans 2400 0 0 0 cell_unit_61/ON
flabel metal1 18400 86850 18400 86850 7 FreeSans 2400 0 0 0 cell_unit_61/V_bias
flabel metal4 11150 88910 11150 88910 5 FreeSans 2400 0 0 0 cell_unit_61/OUT_P
flabel metal4 16410 88910 16410 88910 5 FreeSans 2400 0 0 0 cell_unit_61/OUT_N
flabel metal1 18400 81030 18400 81030 7 FreeSans 2400 0 0 0 cell_unit_61/GND
flabel metal2 13528 85272 13548 85400 7 FreeSans 300 180 0 0 cell_unit_61/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 13528 85094 13548 85222 7 FreeSans 300 180 0 0 cell_unit_61/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 13679 85438 13881 85504 0 FreeSans 300 0 0 0 cell_unit_61/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13554 85094 13612 85110 3 FreeSans 300 90 0 0 cell_unit_61/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 13679 84990 13881 85056 0 FreeSans 300 0 0 0 cell_unit_61/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 13948 85094 14006 85110 3 FreeSans 300 90 0 0 cell_unit_61/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 -610 94810 -610 94810 1 FreeSans 400 0 0 0 inv_1_5/OUT
flabel metal2 -110 94760 -110 94760 1 FreeSans 400 0 0 0 inv_1_5/ON
flabel metal2 -5820 98790 -5820 98790 5 FreeSans 2400 0 0 0 inv_1_5/VDD
flabel metal1 -2820 98790 -2820 98790 5 FreeSans 2400 0 0 0 inv_1_5/GND
flabel metal2 9200 93370 9200 93370 7 FreeSans 2400 0 0 0 cell_unit_62/ON
flabel metal1 9200 96730 9200 96730 7 FreeSans 2400 0 0 0 cell_unit_62/V_bias
flabel metal4 1950 98790 1950 98790 5 FreeSans 2400 0 0 0 cell_unit_62/OUT_P
flabel metal4 7210 98790 7210 98790 5 FreeSans 2400 0 0 0 cell_unit_62/OUT_N
flabel metal1 9200 90910 9200 90910 7 FreeSans 2400 0 0 0 cell_unit_62/GND
flabel metal2 4328 95152 4348 95280 7 FreeSans 300 180 0 0 cell_unit_62/rf_nfet_01v8_aM02W1p65L0p15_0/DRAIN
flabel metal2 4328 94974 4348 95102 7 FreeSans 300 180 0 0 cell_unit_62/rf_nfet_01v8_aM02W1p65L0p15_0/SOURCE
flabel metal1 4479 95318 4681 95384 0 FreeSans 300 0 0 0 cell_unit_62/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4354 94974 4412 94990 3 FreeSans 300 90 0 0 cell_unit_62/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
flabel metal1 4479 94870 4681 94936 0 FreeSans 300 0 0 0 cell_unit_62/rf_nfet_01v8_aM02W1p65L0p15_0/GATE
flabel metal1 4748 94974 4806 94990 3 FreeSans 300 90 0 0 cell_unit_62/rf_nfet_01v8_aM02W1p65L0p15_0/SUBSTRATE
<< end >>
