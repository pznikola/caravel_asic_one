** sch_path: /home/nikolap/Desktop/ASIC/caravel_asic_one/xschem/inv_tb.sch
**.subckt inv_tb
X1 VIN VOUT VDD GND inv
V1 VDD GND 1.8
VIN VIN GND 0
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/nikolap/Desktop/ASIC/PDK/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/nikolap/Desktop/ASIC/PDK/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/nikolap/Desktop/ASIC/PDK/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/nikolap/Desktop/ASIC/PDK/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice



.dc VIN 0 1.8 0.1
.save all


**** end user architecture code
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/nikolap/Desktop/ASIC/caravel_asic_one/xschem/inv.sym
** sch_path: /home/nikolap/Desktop/ASIC/caravel_asic_one/xschem/inv.sch
.subckt inv  IN OUT VDD GND
*.ipin IN
*.opin OUT
*.iopin VDD
*.iopin GND
XM1 OUT IN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.end
