magic
tech sky130B
timestamp 1654635176
<< pwell >>
rect -184 541 -155 564
rect 13 541 42 564
rect 210 541 239 564
rect 407 541 436 564
rect 604 541 633 564
rect 801 541 830 564
rect 998 541 1027 564
rect 1195 541 1224 564
rect 1392 541 1421 564
rect 1589 541 1618 564
rect 0 -631 63 -100
rect 201 -631 252 -100
<< psubdiff >>
rect -184 634 1618 640
rect -184 617 -161 634
rect -144 617 -121 634
rect -104 617 -81 634
rect -64 617 -41 634
rect -24 617 -1 634
rect 16 617 39 634
rect 56 617 79 634
rect 96 617 119 634
rect 136 617 159 634
rect 176 617 199 634
rect 216 617 239 634
rect 256 617 279 634
rect 296 617 319 634
rect 336 617 359 634
rect 376 617 399 634
rect 416 617 439 634
rect 456 617 479 634
rect 496 617 519 634
rect 536 617 559 634
rect 576 617 599 634
rect 616 617 639 634
rect 656 617 679 634
rect 696 617 719 634
rect 736 617 759 634
rect 776 617 799 634
rect 816 617 839 634
rect 856 617 879 634
rect 896 617 919 634
rect 936 617 959 634
rect 976 617 999 634
rect 1016 617 1039 634
rect 1056 617 1079 634
rect 1096 617 1119 634
rect 1136 617 1159 634
rect 1176 617 1199 634
rect 1216 617 1239 634
rect 1256 617 1279 634
rect 1296 617 1319 634
rect 1336 617 1359 634
rect 1376 617 1399 634
rect 1416 617 1439 634
rect 1456 617 1479 634
rect 1496 617 1519 634
rect 1536 617 1559 634
rect 1576 617 1618 634
rect -184 611 1618 617
rect -184 581 -155 611
rect -184 564 -178 581
rect -161 564 -155 581
rect -184 541 -155 564
rect 13 581 42 611
rect 13 564 19 581
rect 36 564 42 581
rect 13 541 42 564
rect 210 581 239 611
rect 210 564 216 581
rect 233 564 239 581
rect 210 541 239 564
rect 407 581 436 611
rect 407 564 413 581
rect 430 564 436 581
rect 407 541 436 564
rect 604 581 633 611
rect 604 564 610 581
rect 627 564 633 581
rect 604 541 633 564
rect 801 581 830 611
rect 801 564 807 581
rect 824 564 830 581
rect 801 541 830 564
rect 998 581 1027 611
rect 998 564 1004 581
rect 1021 564 1027 581
rect 998 541 1027 564
rect 1195 581 1224 611
rect 1195 564 1201 581
rect 1218 564 1224 581
rect 1195 541 1224 564
rect 1392 581 1421 611
rect 1392 564 1398 581
rect 1415 564 1421 581
rect 1392 541 1421 564
rect 1589 581 1618 611
rect 1589 564 1595 581
rect 1612 564 1618 581
rect 1589 541 1618 564
rect -184 37 -155 63
rect -184 20 -178 37
rect -161 20 -155 37
rect -184 -3 -155 20
rect -184 -20 -178 -3
rect -161 -20 -155 -3
rect -184 -43 -155 -20
rect -184 -60 -178 -43
rect -161 -60 -155 -43
rect -184 -83 -155 -60
rect -184 -100 -178 -83
rect -161 -100 -155 -83
rect -184 -132 -155 -100
rect 13 37 42 63
rect 13 20 19 37
rect 36 20 42 37
rect 13 -3 42 20
rect 13 -20 19 -3
rect 36 -20 42 -3
rect 13 -43 42 -20
rect 13 -60 19 -43
rect 36 -60 42 -43
rect 13 -83 42 -60
rect 13 -100 19 -83
rect 36 -100 42 -83
rect 13 -136 42 -100
rect 13 -153 19 -136
rect 36 -153 42 -136
rect 13 -170 42 -153
rect 13 -187 19 -170
rect 36 -187 42 -170
rect 13 -204 42 -187
rect 13 -221 19 -204
rect 36 -221 42 -204
rect 13 -238 42 -221
rect 13 -255 19 -238
rect 36 -255 42 -238
rect 13 -272 42 -255
rect 13 -289 19 -272
rect 36 -289 42 -272
rect 13 -306 42 -289
rect 13 -323 19 -306
rect 36 -323 42 -306
rect 13 -340 42 -323
rect 13 -357 19 -340
rect 36 -357 42 -340
rect 13 -374 42 -357
rect 13 -391 19 -374
rect 36 -391 42 -374
rect 13 -408 42 -391
rect 13 -425 19 -408
rect 36 -425 42 -408
rect 13 -442 42 -425
rect 13 -459 19 -442
rect 36 -459 42 -442
rect 13 -476 42 -459
rect 13 -493 19 -476
rect 36 -493 42 -476
rect 13 -510 42 -493
rect 13 -527 19 -510
rect 36 -527 42 -510
rect 13 -544 42 -527
rect 13 -561 19 -544
rect 36 -561 42 -544
rect 13 -578 42 -561
rect 13 -595 19 -578
rect 36 -595 42 -578
rect -184 -631 -155 -613
rect -184 -648 -178 -631
rect -161 -648 -155 -631
rect -184 -678 -155 -648
rect 13 -631 42 -595
rect 13 -648 19 -631
rect 36 -648 42 -631
rect 13 -678 42 -648
rect 210 37 239 63
rect 210 20 216 37
rect 233 20 239 37
rect 210 -3 239 20
rect 210 -20 216 -3
rect 233 -20 239 -3
rect 210 -43 239 -20
rect 210 -60 216 -43
rect 233 -60 239 -43
rect 210 -83 239 -60
rect 210 -100 216 -83
rect 233 -100 239 -83
rect 210 -136 239 -100
rect 407 37 436 63
rect 407 20 413 37
rect 430 20 436 37
rect 407 -3 436 20
rect 407 -20 413 -3
rect 430 -20 436 -3
rect 407 -43 436 -20
rect 407 -60 413 -43
rect 430 -60 436 -43
rect 407 -83 436 -60
rect 407 -100 413 -83
rect 430 -100 436 -83
rect 407 -132 436 -100
rect 604 37 633 63
rect 604 20 610 37
rect 627 20 633 37
rect 604 -3 633 20
rect 604 -20 610 -3
rect 627 -20 633 -3
rect 604 -43 633 -20
rect 604 -60 610 -43
rect 627 -60 633 -43
rect 604 -83 633 -60
rect 604 -100 610 -83
rect 627 -100 633 -83
rect 604 -132 633 -100
rect 801 37 830 63
rect 801 20 807 37
rect 824 20 830 37
rect 801 -3 830 20
rect 801 -20 807 -3
rect 824 -20 830 -3
rect 801 -43 830 -20
rect 801 -60 807 -43
rect 824 -60 830 -43
rect 801 -83 830 -60
rect 801 -100 807 -83
rect 824 -100 830 -83
rect 801 -132 830 -100
rect 998 37 1027 63
rect 998 20 1004 37
rect 1021 20 1027 37
rect 998 -3 1027 20
rect 998 -20 1004 -3
rect 1021 -20 1027 -3
rect 998 -43 1027 -20
rect 998 -60 1004 -43
rect 1021 -60 1027 -43
rect 998 -83 1027 -60
rect 998 -100 1004 -83
rect 1021 -100 1027 -83
rect 998 -132 1027 -100
rect 1195 37 1224 63
rect 1195 20 1201 37
rect 1218 20 1224 37
rect 1195 -3 1224 20
rect 1195 -20 1201 -3
rect 1218 -20 1224 -3
rect 1195 -43 1224 -20
rect 1195 -60 1201 -43
rect 1218 -60 1224 -43
rect 1195 -83 1224 -60
rect 1195 -100 1201 -83
rect 1218 -100 1224 -83
rect 1195 -132 1224 -100
rect 1392 37 1421 63
rect 1392 20 1398 37
rect 1415 20 1421 37
rect 1392 -3 1421 20
rect 1392 -20 1398 -3
rect 1415 -20 1421 -3
rect 1392 -43 1421 -20
rect 1392 -60 1398 -43
rect 1415 -60 1421 -43
rect 1392 -83 1421 -60
rect 1392 -100 1398 -83
rect 1415 -100 1421 -83
rect 1392 -132 1421 -100
rect 1589 37 1618 63
rect 1589 20 1595 37
rect 1612 20 1618 37
rect 1589 -3 1618 20
rect 1589 -20 1595 -3
rect 1612 -20 1618 -3
rect 1589 -43 1618 -20
rect 1589 -60 1595 -43
rect 1612 -60 1618 -43
rect 1589 -83 1618 -60
rect 1589 -100 1595 -83
rect 1612 -100 1618 -83
rect 1589 -132 1618 -100
rect 210 -153 216 -136
rect 233 -153 239 -136
rect 210 -170 239 -153
rect 210 -187 216 -170
rect 233 -187 239 -170
rect 210 -204 239 -187
rect 210 -221 216 -204
rect 233 -221 239 -204
rect 210 -238 239 -221
rect 210 -255 216 -238
rect 233 -255 239 -238
rect 210 -272 239 -255
rect 210 -289 216 -272
rect 233 -289 239 -272
rect 210 -306 239 -289
rect 210 -323 216 -306
rect 233 -323 239 -306
rect 210 -340 239 -323
rect 210 -357 216 -340
rect 233 -357 239 -340
rect 210 -374 239 -357
rect 210 -391 216 -374
rect 233 -391 239 -374
rect 210 -408 239 -391
rect 210 -425 216 -408
rect 233 -425 239 -408
rect 210 -442 239 -425
rect 210 -459 216 -442
rect 233 -459 239 -442
rect 210 -476 239 -459
rect 210 -493 216 -476
rect 233 -493 239 -476
rect 210 -510 239 -493
rect 210 -527 216 -510
rect 233 -527 239 -510
rect 210 -544 239 -527
rect 210 -561 216 -544
rect 233 -561 239 -544
rect 210 -578 239 -561
rect 210 -595 216 -578
rect 233 -595 239 -578
rect 210 -631 239 -595
rect 210 -648 216 -631
rect 233 -648 239 -631
rect 210 -678 239 -648
rect 407 -631 436 -613
rect 407 -648 413 -631
rect 430 -648 436 -631
rect 407 -678 436 -648
rect 604 -631 633 -613
rect 604 -648 610 -631
rect 627 -648 633 -631
rect 604 -678 633 -648
rect 801 -631 830 -613
rect 801 -648 807 -631
rect 824 -648 830 -631
rect 801 -678 830 -648
rect 998 -631 1027 -613
rect 998 -648 1004 -631
rect 1021 -648 1027 -631
rect 998 -678 1027 -648
rect 1195 -631 1224 -613
rect 1195 -648 1201 -631
rect 1218 -648 1224 -631
rect 1195 -678 1224 -648
rect 1392 -631 1421 -613
rect 1392 -648 1398 -631
rect 1415 -648 1421 -631
rect 1392 -678 1421 -648
rect 1589 -631 1618 -613
rect 1589 -648 1595 -631
rect 1612 -648 1618 -631
rect 1589 -678 1618 -648
rect -184 -684 1618 -678
rect -184 -701 -161 -684
rect -144 -701 -121 -684
rect -104 -701 -81 -684
rect -64 -701 -41 -684
rect -24 -701 -1 -684
rect 16 -701 39 -684
rect 56 -701 79 -684
rect 96 -701 119 -684
rect 136 -701 159 -684
rect 176 -701 199 -684
rect 216 -701 239 -684
rect 256 -701 279 -684
rect 296 -701 319 -684
rect 336 -701 359 -684
rect 376 -701 399 -684
rect 416 -701 439 -684
rect 456 -701 479 -684
rect 496 -701 519 -684
rect 536 -701 559 -684
rect 576 -701 599 -684
rect 616 -701 639 -684
rect 656 -701 679 -684
rect 696 -701 719 -684
rect 736 -701 759 -684
rect 776 -701 799 -684
rect 816 -701 839 -684
rect 856 -701 879 -684
rect 896 -701 919 -684
rect 936 -701 959 -684
rect 976 -701 999 -684
rect 1016 -701 1039 -684
rect 1056 -701 1079 -684
rect 1096 -701 1119 -684
rect 1136 -701 1159 -684
rect 1176 -701 1199 -684
rect 1216 -701 1239 -684
rect 1256 -701 1279 -684
rect 1296 -701 1319 -684
rect 1336 -701 1359 -684
rect 1376 -701 1399 -684
rect 1416 -701 1439 -684
rect 1456 -701 1479 -684
rect 1496 -701 1519 -684
rect 1536 -701 1559 -684
rect 1576 -701 1618 -684
rect -184 -707 1618 -701
<< psubdiffcont >>
rect -161 617 -144 634
rect -121 617 -104 634
rect -81 617 -64 634
rect -41 617 -24 634
rect -1 617 16 634
rect 39 617 56 634
rect 79 617 96 634
rect 119 617 136 634
rect 159 617 176 634
rect 199 617 216 634
rect 239 617 256 634
rect 279 617 296 634
rect 319 617 336 634
rect 359 617 376 634
rect 399 617 416 634
rect 439 617 456 634
rect 479 617 496 634
rect 519 617 536 634
rect 559 617 576 634
rect 599 617 616 634
rect 639 617 656 634
rect 679 617 696 634
rect 719 617 736 634
rect 759 617 776 634
rect 799 617 816 634
rect 839 617 856 634
rect 879 617 896 634
rect 919 617 936 634
rect 959 617 976 634
rect 999 617 1016 634
rect 1039 617 1056 634
rect 1079 617 1096 634
rect 1119 617 1136 634
rect 1159 617 1176 634
rect 1199 617 1216 634
rect 1239 617 1256 634
rect 1279 617 1296 634
rect 1319 617 1336 634
rect 1359 617 1376 634
rect 1399 617 1416 634
rect 1439 617 1456 634
rect 1479 617 1496 634
rect 1519 617 1536 634
rect 1559 617 1576 634
rect -178 564 -161 581
rect 19 564 36 581
rect 216 564 233 581
rect 413 564 430 581
rect 610 564 627 581
rect 807 564 824 581
rect 1004 564 1021 581
rect 1201 564 1218 581
rect 1398 564 1415 581
rect 1595 564 1612 581
rect -178 20 -161 37
rect -178 -20 -161 -3
rect -178 -60 -161 -43
rect -178 -100 -161 -83
rect 19 20 36 37
rect 19 -20 36 -3
rect 19 -60 36 -43
rect 19 -100 36 -83
rect 19 -153 36 -136
rect 19 -187 36 -170
rect 19 -221 36 -204
rect 19 -255 36 -238
rect 19 -289 36 -272
rect 19 -323 36 -306
rect 19 -357 36 -340
rect 19 -391 36 -374
rect 19 -425 36 -408
rect 19 -459 36 -442
rect 19 -493 36 -476
rect 19 -527 36 -510
rect 19 -561 36 -544
rect 19 -595 36 -578
rect -178 -648 -161 -631
rect 19 -648 36 -631
rect 216 20 233 37
rect 216 -20 233 -3
rect 216 -60 233 -43
rect 216 -100 233 -83
rect 413 20 430 37
rect 413 -20 430 -3
rect 413 -60 430 -43
rect 413 -100 430 -83
rect 610 20 627 37
rect 610 -20 627 -3
rect 610 -60 627 -43
rect 610 -100 627 -83
rect 807 20 824 37
rect 807 -20 824 -3
rect 807 -60 824 -43
rect 807 -100 824 -83
rect 1004 20 1021 37
rect 1004 -20 1021 -3
rect 1004 -60 1021 -43
rect 1004 -100 1021 -83
rect 1201 20 1218 37
rect 1201 -20 1218 -3
rect 1201 -60 1218 -43
rect 1201 -100 1218 -83
rect 1398 20 1415 37
rect 1398 -20 1415 -3
rect 1398 -60 1415 -43
rect 1398 -100 1415 -83
rect 1595 20 1612 37
rect 1595 -20 1612 -3
rect 1595 -60 1612 -43
rect 1595 -100 1612 -83
rect 216 -153 233 -136
rect 216 -187 233 -170
rect 216 -221 233 -204
rect 216 -255 233 -238
rect 216 -289 233 -272
rect 216 -323 233 -306
rect 216 -357 233 -340
rect 216 -391 233 -374
rect 216 -425 233 -408
rect 216 -459 233 -442
rect 216 -493 233 -476
rect 216 -527 233 -510
rect 216 -561 233 -544
rect 216 -595 233 -578
rect 216 -648 233 -631
rect 413 -648 430 -631
rect 610 -648 627 -631
rect 807 -648 824 -631
rect 1004 -648 1021 -631
rect 1201 -648 1218 -631
rect 1398 -648 1415 -631
rect 1595 -648 1612 -631
rect -161 -701 -144 -684
rect -121 -701 -104 -684
rect -81 -701 -64 -684
rect -41 -701 -24 -684
rect -1 -701 16 -684
rect 39 -701 56 -684
rect 79 -701 96 -684
rect 119 -701 136 -684
rect 159 -701 176 -684
rect 199 -701 216 -684
rect 239 -701 256 -684
rect 279 -701 296 -684
rect 319 -701 336 -684
rect 359 -701 376 -684
rect 399 -701 416 -684
rect 439 -701 456 -684
rect 479 -701 496 -684
rect 519 -701 536 -684
rect 559 -701 576 -684
rect 599 -701 616 -684
rect 639 -701 656 -684
rect 679 -701 696 -684
rect 719 -701 736 -684
rect 759 -701 776 -684
rect 799 -701 816 -684
rect 839 -701 856 -684
rect 879 -701 896 -684
rect 919 -701 936 -684
rect 959 -701 976 -684
rect 999 -701 1016 -684
rect 1039 -701 1056 -684
rect 1079 -701 1096 -684
rect 1119 -701 1136 -684
rect 1159 -701 1176 -684
rect 1199 -701 1216 -684
rect 1239 -701 1256 -684
rect 1279 -701 1296 -684
rect 1319 -701 1336 -684
rect 1359 -701 1376 -684
rect 1399 -701 1416 -684
rect 1439 -701 1456 -684
rect 1479 -701 1496 -684
rect 1519 -701 1536 -684
rect 1559 -701 1576 -684
<< locali >>
rect -178 581 -161 634
rect -144 617 -121 634
rect -104 617 -81 634
rect -64 617 -41 634
rect -24 617 -1 634
rect 16 617 39 634
rect 56 617 79 634
rect 96 617 119 634
rect 136 617 159 634
rect 176 617 199 634
rect 216 617 239 634
rect 256 617 279 634
rect 296 617 319 634
rect 336 617 359 634
rect 376 617 399 634
rect 416 617 439 634
rect 456 617 479 634
rect 496 617 519 634
rect 536 617 559 634
rect 576 617 599 634
rect 616 617 639 634
rect 656 617 679 634
rect 696 617 719 634
rect 736 617 759 634
rect 776 617 799 634
rect 816 617 839 634
rect 856 617 879 634
rect 896 617 919 634
rect 936 617 959 634
rect 976 617 999 634
rect 1016 617 1039 634
rect 1056 617 1079 634
rect 1096 617 1119 634
rect 1136 617 1159 634
rect 1176 617 1199 634
rect 1216 617 1239 634
rect 1256 617 1279 634
rect 1296 617 1319 634
rect 1336 617 1359 634
rect 1376 617 1399 634
rect 1416 617 1439 634
rect 1456 617 1479 634
rect 1496 617 1519 634
rect 1536 617 1559 634
rect 1576 617 1612 634
rect -178 541 -161 564
rect 19 581 36 617
rect 19 541 36 564
rect 216 581 233 617
rect 216 541 233 564
rect 413 581 430 617
rect 413 541 430 564
rect 610 581 627 617
rect 610 541 627 564
rect 807 581 824 617
rect 807 541 824 564
rect 1004 581 1021 617
rect 1004 541 1021 564
rect 1201 581 1218 617
rect 1201 541 1218 564
rect 1398 581 1415 617
rect 1398 541 1415 564
rect 1595 581 1612 617
rect 1595 541 1612 564
rect -178 37 -161 66
rect -178 -3 -161 20
rect -178 -43 -161 -20
rect -178 -83 -161 -60
rect -178 -126 -161 -100
rect 19 37 36 66
rect 19 -3 36 20
rect 19 -43 36 -20
rect 19 -83 36 -60
rect 19 -123 36 -100
rect 19 -159 36 -153
rect 19 -195 36 -187
rect 19 -231 36 -221
rect 19 -267 36 -255
rect 19 -303 36 -289
rect 19 -339 36 -323
rect 19 -374 36 -357
rect 19 -408 36 -392
rect 19 -442 36 -428
rect 19 -476 36 -464
rect 19 -510 36 -500
rect 19 -544 36 -536
rect 19 -578 36 -572
rect -178 -631 -161 -608
rect -178 -701 -161 -648
rect 19 -631 36 -608
rect 19 -684 36 -648
rect 216 37 233 66
rect 216 -3 233 20
rect 216 -43 233 -20
rect 216 -83 233 -60
rect 216 -123 233 -100
rect 413 37 430 66
rect 413 -3 430 20
rect 413 -43 430 -20
rect 413 -83 430 -60
rect 413 -126 430 -100
rect 610 37 627 66
rect 610 -3 627 20
rect 610 -43 627 -20
rect 610 -83 627 -60
rect 610 -126 627 -100
rect 807 37 824 66
rect 807 -3 824 20
rect 807 -43 824 -20
rect 807 -83 824 -60
rect 807 -126 824 -100
rect 1004 37 1021 66
rect 1004 -3 1021 20
rect 1004 -43 1021 -20
rect 1004 -83 1021 -60
rect 1004 -126 1021 -100
rect 1201 37 1218 66
rect 1201 -3 1218 20
rect 1201 -43 1218 -20
rect 1201 -83 1218 -60
rect 1201 -126 1218 -100
rect 1398 37 1415 66
rect 1398 -3 1415 20
rect 1398 -43 1415 -20
rect 1398 -83 1415 -60
rect 1398 -126 1415 -100
rect 1595 37 1612 66
rect 1595 -3 1612 20
rect 1595 -43 1612 -20
rect 1595 -83 1612 -60
rect 1595 -126 1612 -100
rect 216 -159 233 -153
rect 216 -195 233 -187
rect 216 -231 233 -221
rect 216 -267 233 -255
rect 216 -303 233 -289
rect 216 -339 233 -323
rect 216 -374 233 -357
rect 216 -408 233 -392
rect 216 -442 233 -428
rect 216 -476 233 -464
rect 216 -510 233 -500
rect 216 -544 233 -536
rect 216 -578 233 -572
rect 216 -631 233 -608
rect 216 -684 233 -648
rect 413 -631 430 -608
rect 413 -684 430 -648
rect 610 -631 627 -608
rect 610 -684 627 -648
rect 807 -631 824 -608
rect 807 -684 824 -648
rect 1004 -631 1021 -608
rect 1004 -684 1021 -648
rect 1201 -631 1218 -608
rect 1201 -684 1218 -648
rect 1398 -631 1415 -608
rect 1398 -684 1415 -648
rect 1595 -631 1612 -608
rect 1595 -684 1612 -648
rect -144 -701 -121 -684
rect -104 -701 -81 -684
rect -64 -701 -41 -684
rect -24 -701 -1 -684
rect 16 -701 39 -684
rect 56 -701 79 -684
rect 96 -701 119 -684
rect 136 -701 159 -684
rect 176 -701 199 -684
rect 216 -701 239 -684
rect 256 -701 279 -684
rect 296 -701 319 -684
rect 336 -701 359 -684
rect 376 -701 399 -684
rect 416 -701 439 -684
rect 456 -701 479 -684
rect 496 -701 519 -684
rect 536 -701 559 -684
rect 576 -701 599 -684
rect 616 -701 639 -684
rect 656 -701 679 -684
rect 696 -701 719 -684
rect 736 -701 759 -684
rect 776 -701 799 -684
rect 816 -701 839 -684
rect 856 -701 879 -684
rect 896 -701 919 -684
rect 936 -701 959 -684
rect 976 -701 999 -684
rect 1016 -701 1039 -684
rect 1056 -701 1079 -684
rect 1096 -701 1119 -684
rect 1136 -701 1159 -684
rect 1176 -701 1199 -684
rect 1216 -701 1239 -684
rect 1256 -701 1279 -684
rect 1296 -701 1319 -684
rect 1336 -701 1359 -684
rect 1376 -701 1399 -684
rect 1416 -701 1439 -684
rect 1456 -701 1479 -684
rect 1496 -701 1519 -684
rect 1536 -701 1559 -684
rect 1576 -701 1612 -684
<< viali >>
rect -161 617 -144 634
rect -121 617 -104 634
rect -81 617 -64 634
rect -41 617 -24 634
rect -1 617 16 634
rect 39 617 56 634
rect 79 617 96 634
rect 119 617 136 634
rect 159 617 176 634
rect 199 617 216 634
rect 239 617 256 634
rect 279 617 296 634
rect 319 617 336 634
rect 359 617 376 634
rect 399 617 416 634
rect 439 617 456 634
rect 479 617 496 634
rect 519 617 536 634
rect 559 617 576 634
rect 599 617 616 634
rect 639 617 656 634
rect 679 617 696 634
rect 719 617 736 634
rect 759 617 776 634
rect 799 617 816 634
rect 839 617 856 634
rect 879 617 896 634
rect 919 617 936 634
rect 959 617 976 634
rect 999 617 1016 634
rect 1039 617 1056 634
rect 1079 617 1096 634
rect 1119 617 1136 634
rect 1159 617 1176 634
rect 1199 617 1216 634
rect 1239 617 1256 634
rect 1279 617 1296 634
rect 1319 617 1336 634
rect 1359 617 1376 634
rect 1399 617 1416 634
rect 1439 617 1456 634
rect 1479 617 1496 634
rect 1519 617 1536 634
rect 1559 617 1576 634
rect -178 564 -161 581
rect 19 564 36 581
rect 216 564 233 581
rect 413 564 430 581
rect 610 564 627 581
rect 807 564 824 581
rect 1004 564 1021 581
rect 1201 564 1218 581
rect 1398 564 1415 581
rect 1595 564 1612 581
rect -178 20 -161 37
rect -178 -20 -161 -3
rect -178 -60 -161 -43
rect -178 -100 -161 -83
rect 19 20 36 37
rect 19 -20 36 -3
rect 19 -60 36 -43
rect 19 -100 36 -83
rect 19 -136 36 -123
rect 19 -140 36 -136
rect 19 -170 36 -159
rect 19 -176 36 -170
rect 19 -204 36 -195
rect 19 -212 36 -204
rect 19 -238 36 -231
rect 19 -248 36 -238
rect 19 -272 36 -267
rect 19 -284 36 -272
rect 19 -306 36 -303
rect 19 -320 36 -306
rect 19 -340 36 -339
rect 19 -356 36 -340
rect 19 -391 36 -375
rect 19 -392 36 -391
rect 19 -425 36 -411
rect 19 -428 36 -425
rect 19 -459 36 -447
rect 19 -464 36 -459
rect 19 -493 36 -483
rect 19 -500 36 -493
rect 19 -527 36 -519
rect 19 -536 36 -527
rect 19 -561 36 -555
rect 19 -572 36 -561
rect 19 -595 36 -591
rect 19 -608 36 -595
rect -178 -648 -161 -631
rect 19 -648 36 -631
rect 216 20 233 37
rect 216 -20 233 -3
rect 216 -60 233 -43
rect 216 -100 233 -83
rect 216 -136 233 -123
rect 413 20 430 37
rect 413 -20 430 -3
rect 413 -60 430 -43
rect 413 -100 430 -83
rect 610 20 627 37
rect 610 -20 627 -3
rect 610 -60 627 -43
rect 610 -100 627 -83
rect 807 20 824 37
rect 807 -20 824 -3
rect 807 -60 824 -43
rect 807 -100 824 -83
rect 1004 20 1021 37
rect 1004 -20 1021 -3
rect 1004 -60 1021 -43
rect 1004 -100 1021 -83
rect 1201 20 1218 37
rect 1201 -20 1218 -3
rect 1201 -60 1218 -43
rect 1201 -100 1218 -83
rect 1398 20 1415 37
rect 1398 -20 1415 -3
rect 1398 -60 1415 -43
rect 1398 -100 1415 -83
rect 1595 20 1612 37
rect 1595 -20 1612 -3
rect 1595 -60 1612 -43
rect 1595 -100 1612 -83
rect 216 -140 233 -136
rect 216 -170 233 -159
rect 216 -176 233 -170
rect 216 -204 233 -195
rect 216 -212 233 -204
rect 216 -238 233 -231
rect 216 -248 233 -238
rect 216 -272 233 -267
rect 216 -284 233 -272
rect 216 -306 233 -303
rect 216 -320 233 -306
rect 216 -340 233 -339
rect 216 -356 233 -340
rect 216 -391 233 -375
rect 216 -392 233 -391
rect 216 -425 233 -411
rect 216 -428 233 -425
rect 216 -459 233 -447
rect 216 -464 233 -459
rect 216 -493 233 -483
rect 216 -500 233 -493
rect 216 -527 233 -519
rect 216 -536 233 -527
rect 216 -561 233 -555
rect 216 -572 233 -561
rect 216 -595 233 -591
rect 216 -608 233 -595
rect 1595 -608 1612 -591
rect 216 -648 233 -631
rect 413 -648 430 -631
rect 610 -648 627 -631
rect 807 -648 824 -631
rect 1004 -648 1021 -631
rect 1201 -648 1218 -631
rect 1398 -648 1415 -631
rect 1595 -648 1612 -631
rect -161 -701 -144 -684
rect -121 -701 -104 -684
rect -81 -701 -64 -684
rect -41 -701 -24 -684
rect -1 -701 16 -684
rect 39 -701 56 -684
rect 79 -701 96 -684
rect 119 -701 136 -684
rect 159 -701 176 -684
rect 199 -701 216 -684
rect 239 -701 256 -684
rect 279 -701 296 -684
rect 319 -701 336 -684
rect 359 -701 376 -684
rect 399 -701 416 -684
rect 439 -701 456 -684
rect 479 -701 496 -684
rect 519 -701 536 -684
rect 559 -701 576 -684
rect 599 -701 616 -684
rect 639 -701 656 -684
rect 679 -701 696 -684
rect 719 -701 736 -684
rect 759 -701 776 -684
rect 799 -701 816 -684
rect 839 -701 856 -684
rect 879 -701 896 -684
rect 919 -701 936 -684
rect 959 -701 976 -684
rect 999 -701 1016 -684
rect 1039 -701 1056 -684
rect 1079 -701 1096 -684
rect 1119 -701 1136 -684
rect 1159 -701 1176 -684
rect 1199 -701 1216 -684
rect 1239 -701 1256 -684
rect 1279 -701 1296 -684
rect 1319 -701 1336 -684
rect 1359 -701 1376 -684
rect 1399 -701 1416 -684
rect 1439 -701 1456 -684
rect 1479 -701 1496 -684
rect 1519 -701 1536 -684
rect 1559 -701 1576 -684
<< metal1 >>
rect -184 634 1618 640
rect -184 617 -161 634
rect -144 617 -121 634
rect -104 617 -81 634
rect -64 617 -41 634
rect -24 617 -1 634
rect 16 617 39 634
rect 56 617 79 634
rect 96 617 119 634
rect 136 617 159 634
rect 176 617 199 634
rect 216 617 239 634
rect 256 617 279 634
rect 296 617 319 634
rect 336 617 359 634
rect 376 617 399 634
rect 416 617 439 634
rect 456 617 479 634
rect 496 617 519 634
rect 536 617 559 634
rect 576 617 599 634
rect 616 617 639 634
rect 656 617 679 634
rect 696 617 719 634
rect 736 617 759 634
rect 776 617 799 634
rect 816 617 839 634
rect 856 617 879 634
rect 896 617 919 634
rect 936 617 959 634
rect 976 617 999 634
rect 1016 617 1039 634
rect 1056 617 1079 634
rect 1096 617 1119 634
rect 1136 617 1159 634
rect 1176 617 1199 634
rect 1216 617 1239 634
rect 1256 617 1279 634
rect 1296 617 1319 634
rect 1336 617 1359 634
rect 1376 617 1399 634
rect 1416 617 1439 634
rect 1456 617 1479 634
rect 1496 617 1519 634
rect 1536 617 1559 634
rect 1576 617 1618 634
rect -184 611 1618 617
rect -184 581 42 611
rect -184 564 -178 581
rect -161 564 19 581
rect 36 564 42 581
rect -184 522 -155 564
rect -127 522 -101 564
rect -84 522 -58 564
rect -41 522 -15 564
rect 13 522 42 564
rect 210 581 239 611
rect 210 564 216 581
rect 233 564 239 581
rect 210 541 239 564
rect 407 581 436 611
rect 407 564 413 581
rect 430 564 436 581
rect 407 541 436 564
rect 604 581 633 611
rect 604 564 610 581
rect 627 564 633 581
rect 604 541 633 564
rect 801 581 830 611
rect 801 564 807 581
rect 824 564 830 581
rect 801 541 830 564
rect 998 581 1027 611
rect 998 564 1004 581
rect 1021 564 1027 581
rect 998 541 1027 564
rect 1195 581 1224 611
rect 1195 564 1201 581
rect 1218 564 1224 581
rect 1195 541 1224 564
rect 1392 581 1618 611
rect 1392 564 1398 581
rect 1415 564 1595 581
rect 1612 564 1618 581
rect 1392 522 1421 564
rect 1449 522 1475 564
rect 1492 522 1518 564
rect 1535 522 1561 564
rect 1589 522 1618 564
rect -184 37 -155 75
rect -184 20 -178 37
rect -161 33 -155 37
rect -127 33 -101 75
rect -84 33 -58 75
rect -41 33 -15 75
rect 13 37 42 75
rect 13 33 19 37
rect -161 20 19 33
rect 36 20 42 37
rect -184 0 42 20
rect -184 -3 -155 0
rect -184 -20 -178 -3
rect -161 -20 -155 -3
rect -184 -43 -155 -20
rect -184 -60 -178 -43
rect -161 -60 -155 -43
rect -184 -67 -155 -60
rect 13 -3 42 0
rect 13 -20 19 -3
rect 36 -20 42 -3
rect 13 -43 42 -20
rect 13 -60 19 -43
rect 36 -60 42 -43
rect 13 -67 42 -60
rect -184 -83 42 -67
rect -184 -100 -178 -83
rect -161 -100 19 -83
rect 36 -100 42 -83
rect -184 -142 -155 -100
rect -127 -142 -101 -100
rect -84 -142 -58 -100
rect -41 -142 -15 -100
rect 13 -123 42 -100
rect 13 -140 19 -123
rect 36 -140 42 -123
rect 13 -159 42 -140
rect 13 -176 19 -159
rect 36 -176 42 -159
rect 13 -195 42 -176
rect 13 -212 19 -195
rect 36 -212 42 -195
rect 13 -231 42 -212
rect 13 -248 19 -231
rect 36 -248 42 -231
rect 13 -267 42 -248
rect 13 -284 19 -267
rect 36 -284 42 -267
rect 13 -303 42 -284
rect 13 -320 19 -303
rect 36 -320 42 -303
rect 13 -339 42 -320
rect 13 -356 19 -339
rect 36 -356 42 -339
rect 13 -375 42 -356
rect 13 -392 19 -375
rect 36 -392 42 -375
rect 13 -411 42 -392
rect 13 -428 19 -411
rect 36 -428 42 -411
rect 13 -447 42 -428
rect 13 -464 19 -447
rect 36 -464 42 -447
rect 13 -483 42 -464
rect 13 -500 19 -483
rect 36 -500 42 -483
rect 13 -519 42 -500
rect 13 -536 19 -519
rect 36 -536 42 -519
rect 13 -555 42 -536
rect 13 -572 19 -555
rect 36 -572 42 -555
rect -184 -631 -155 -589
rect -127 -631 -101 -589
rect -84 -631 -58 -589
rect -41 -631 -15 -589
rect 13 -591 42 -572
rect 13 -608 19 -591
rect 36 -608 42 -591
rect 13 -631 42 -608
rect -184 -648 -178 -631
rect -161 -648 19 -631
rect 36 -648 42 -631
rect -184 -678 42 -648
rect 210 37 239 63
rect 210 20 216 37
rect 233 20 239 37
rect 210 -3 239 20
rect 210 -20 216 -3
rect 233 -20 239 -3
rect 210 -43 239 -20
rect 210 -60 216 -43
rect 233 -60 239 -43
rect 210 -83 239 -60
rect 210 -100 216 -83
rect 233 -100 239 -83
rect 210 -123 239 -100
rect 210 -140 216 -123
rect 233 -140 239 -123
rect 407 37 436 63
rect 407 20 413 37
rect 430 20 436 37
rect 407 -3 436 20
rect 407 -20 413 -3
rect 430 -20 436 -3
rect 407 -43 436 -20
rect 407 -60 413 -43
rect 430 -60 436 -43
rect 407 -83 436 -60
rect 407 -100 413 -83
rect 430 -100 436 -83
rect 407 -132 436 -100
rect 604 37 633 63
rect 604 20 610 37
rect 627 20 633 37
rect 604 -3 633 20
rect 604 -20 610 -3
rect 627 -20 633 -3
rect 604 -43 633 -20
rect 604 -60 610 -43
rect 627 -60 633 -43
rect 604 -83 633 -60
rect 604 -100 610 -83
rect 627 -100 633 -83
rect 604 -132 633 -100
rect 801 37 830 63
rect 801 20 807 37
rect 824 20 830 37
rect 801 -3 830 20
rect 801 -20 807 -3
rect 824 -20 830 -3
rect 801 -43 830 -20
rect 801 -60 807 -43
rect 824 -60 830 -43
rect 801 -83 830 -60
rect 801 -100 807 -83
rect 824 -100 830 -83
rect 801 -132 830 -100
rect 998 37 1027 63
rect 998 20 1004 37
rect 1021 20 1027 37
rect 998 -3 1027 20
rect 998 -20 1004 -3
rect 1021 -20 1027 -3
rect 998 -43 1027 -20
rect 998 -60 1004 -43
rect 1021 -60 1027 -43
rect 998 -83 1027 -60
rect 998 -100 1004 -83
rect 1021 -100 1027 -83
rect 998 -132 1027 -100
rect 1195 37 1224 63
rect 1195 20 1201 37
rect 1218 20 1224 37
rect 1195 -3 1224 20
rect 1195 -20 1201 -3
rect 1218 -20 1224 -3
rect 1195 -43 1224 -20
rect 1195 -60 1201 -43
rect 1218 -60 1224 -43
rect 1195 -83 1224 -60
rect 1195 -100 1201 -83
rect 1218 -100 1224 -83
rect 1195 -132 1224 -100
rect 1392 37 1421 75
rect 1392 20 1398 37
rect 1415 33 1421 37
rect 1449 33 1475 75
rect 1492 33 1518 75
rect 1535 33 1561 75
rect 1589 37 1618 75
rect 1589 33 1595 37
rect 1415 20 1595 33
rect 1612 20 1618 37
rect 1392 0 1618 20
rect 1392 -3 1421 0
rect 1392 -20 1398 -3
rect 1415 -20 1421 -3
rect 1392 -43 1421 -20
rect 1392 -60 1398 -43
rect 1415 -60 1421 -43
rect 1392 -67 1421 -60
rect 1589 -3 1618 0
rect 1589 -20 1595 -3
rect 1612 -20 1618 -3
rect 1589 -43 1618 -20
rect 1589 -60 1595 -43
rect 1612 -60 1618 -43
rect 1589 -67 1618 -60
rect 1392 -83 1618 -67
rect 1392 -100 1398 -83
rect 1415 -100 1595 -83
rect 1612 -100 1618 -83
rect 210 -159 239 -140
rect 1392 -142 1421 -100
rect 1449 -142 1475 -100
rect 1492 -142 1518 -100
rect 1535 -142 1561 -100
rect 1589 -142 1618 -100
rect 210 -176 216 -159
rect 233 -176 239 -159
rect 210 -195 239 -176
rect 210 -212 216 -195
rect 233 -212 239 -195
rect 210 -231 239 -212
rect 210 -248 216 -231
rect 233 -248 239 -231
rect 210 -267 239 -248
rect 210 -284 216 -267
rect 233 -284 239 -267
rect 210 -303 239 -284
rect 210 -320 216 -303
rect 233 -320 239 -303
rect 210 -339 239 -320
rect 210 -356 216 -339
rect 233 -356 239 -339
rect 210 -375 239 -356
rect 210 -392 216 -375
rect 233 -392 239 -375
rect 210 -411 239 -392
rect 210 -428 216 -411
rect 233 -428 239 -411
rect 210 -447 239 -428
rect 210 -464 216 -447
rect 233 -464 239 -447
rect 210 -483 239 -464
rect 210 -500 216 -483
rect 233 -500 239 -483
rect 210 -519 239 -500
rect 210 -536 216 -519
rect 233 -536 239 -519
rect 210 -555 239 -536
rect 210 -572 216 -555
rect 233 -572 239 -555
rect 210 -591 239 -572
rect 210 -608 216 -591
rect 233 -608 239 -591
rect 210 -631 239 -608
rect 210 -648 216 -631
rect 233 -648 239 -631
rect 210 -678 239 -648
rect 407 -631 436 -613
rect 407 -648 413 -631
rect 430 -648 436 -631
rect 407 -678 436 -648
rect 604 -631 633 -613
rect 604 -648 610 -631
rect 627 -648 633 -631
rect 604 -678 633 -648
rect 801 -631 830 -613
rect 801 -648 807 -631
rect 824 -648 830 -631
rect 801 -678 830 -648
rect 998 -631 1027 -613
rect 998 -648 1004 -631
rect 1021 -648 1027 -631
rect 998 -678 1027 -648
rect 1195 -631 1224 -613
rect 1195 -648 1201 -631
rect 1218 -648 1224 -631
rect 1195 -678 1224 -648
rect 1392 -631 1421 -589
rect 1449 -631 1475 -589
rect 1492 -631 1518 -589
rect 1535 -631 1561 -589
rect 1589 -591 1618 -589
rect 1589 -608 1595 -591
rect 1612 -608 1618 -591
rect 1589 -631 1618 -608
rect 1392 -648 1398 -631
rect 1415 -648 1595 -631
rect 1612 -648 1618 -631
rect 1392 -678 1618 -648
rect -184 -684 1618 -678
rect -184 -701 -161 -684
rect -144 -701 -121 -684
rect -104 -701 -81 -684
rect -64 -701 -41 -684
rect -24 -701 -1 -684
rect 16 -701 39 -684
rect 56 -701 79 -684
rect 96 -701 119 -684
rect 136 -701 159 -684
rect 176 -701 199 -684
rect 216 -701 239 -684
rect 256 -701 279 -684
rect 296 -701 319 -684
rect 336 -701 359 -684
rect 376 -701 399 -684
rect 416 -701 439 -684
rect 456 -701 479 -684
rect 496 -701 519 -684
rect 536 -701 559 -684
rect 576 -701 599 -684
rect 616 -701 639 -684
rect 656 -701 679 -684
rect 696 -701 719 -684
rect 736 -701 759 -684
rect 776 -701 799 -684
rect 816 -701 839 -684
rect 856 -701 879 -684
rect 896 -701 919 -684
rect 936 -701 959 -684
rect 976 -701 999 -684
rect 1016 -701 1039 -684
rect 1056 -701 1079 -684
rect 1096 -701 1119 -684
rect 1136 -701 1159 -684
rect 1176 -701 1199 -684
rect 1216 -701 1239 -684
rect 1256 -701 1279 -684
rect 1296 -701 1319 -684
rect 1336 -701 1359 -684
rect 1376 -701 1399 -684
rect 1416 -701 1439 -684
rect 1456 -701 1479 -684
rect 1496 -701 1519 -684
rect 1536 -701 1559 -684
rect 1576 -701 1618 -684
rect -184 -707 1618 -701
use rf_nfet_01v8_aM02W5p00L0p15  rf_nfet_01v8_aM02W5p00L0p15_0
timestamp 1654634331
transform 1 0 -5 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1654628751
transform -1 0 257 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_1
timestamp 1654628751
transform 1 0 192 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_2
timestamp 1654628751
transform 1 0 389 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_3
timestamp 1654628751
transform 1 0 586 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_4
timestamp 1654628751
transform 1 0 783 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_5
timestamp 1654628751
transform 1 0 980 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_6
timestamp 1654628751
transform 1 0 1177 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_7
timestamp 1654628751
transform 1 0 1177 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_8
timestamp 1654628751
transform 1 0 980 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_9
timestamp 1654628751
transform 1 0 783 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_10
timestamp 1654628751
transform 1 0 586 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_11
timestamp 1654628751
transform 1 0 389 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_12
timestamp 1654628751
transform 1 0 192 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_13
timestamp 1654628751
transform -1 0 60 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_14
timestamp 1654628751
transform -1 0 1636 0 -1 602
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_15
timestamp 1654628751
transform -1 0 1636 0 1 -669
box 5 5 257 602
use sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W5p00L0p15_16
timestamp 1654628751
transform -1 0 60 0 1 -669
box 5 5 257 602
<< labels >>
flabel metal1 s 210 -614 239 -606 7 FreeSans 150 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 13 -614 42 -606 7 FreeSans 150 90 0 0 SUBSTRATE
port 4 nsew
<< end >>
