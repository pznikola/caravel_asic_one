magic
tech sky130B
magscale 1 2
timestamp 1654082934
<< pwell >>
rect -96 -34 814 1130
<< metal1 >>
rect -44 920 764 1080
rect -54 16 -44 448
rect 26 16 36 448
rect 146 -106 180 172
rect 259 0 461 20
rect 259 -60 273 0
rect 447 -60 461 0
rect 540 -106 574 172
rect 684 16 694 448
rect 764 16 774 448
rect 146 -140 574 -106
<< via1 >>
rect -44 16 26 448
rect 273 -60 447 0
rect 694 16 764 448
<< metal2 >>
rect -44 448 26 458
rect -50 282 -44 410
rect 694 448 764 458
rect 26 282 30 410
rect 612 104 694 232
rect -44 10 26 16
rect 764 104 770 232
rect 694 10 764 16
rect -50 -240 30 10
rect -60 -260 30 -240
rect -60 -330 -50 -260
rect 20 -330 30 -260
rect -60 -340 30 -330
rect 270 0 450 10
rect 270 -60 273 0
rect 447 -60 450 0
rect 270 -350 450 -60
rect 690 -240 770 10
rect 690 -260 780 -240
rect 690 -330 700 -260
rect 770 -330 780 -260
rect 690 -340 780 -330
<< via2 >>
rect -50 -330 20 -260
rect 700 -330 770 -260
<< metal3 >>
rect -320 -240 -230 90
rect 950 -240 1040 90
rect -320 -260 40 -240
rect -320 -330 -50 -260
rect 20 -330 40 -260
rect -320 -350 40 -330
rect 680 -260 1040 -240
rect 680 -330 700 -260
rect 770 -330 1040 -260
rect 1610 -270 1760 180
rect 680 -350 1040 -330
<< metal4 >>
rect -990 -260 -840 180
rect 1610 -270 1760 180
use rf_nfet_01v8_aM02W1p65L0p15  rf_nfet_01v8_aM02W1p65L0p15_0
timestamp 1648127584
transform 1 0 98 0 1 -10
box 10 10 514 524
use sky130_fd_pr__cap_mim_m3_1_V3VADT  sky130_fd_pr__cap_mim_m3_1_V3VADT_0
timestamp 1654038913
transform 1 0 -655 0 1 430
box -480 -430 479 430
use sky130_fd_pr__cap_mim_m3_1_V3VADT  sky130_fd_pr__cap_mim_m3_1_V3VADT_1
timestamp 1654038913
transform -1 0 1423 0 1 430
box -480 -430 479 430
use sky130_fd_pr__res_xhigh_po_0p35_WX6KG8  sky130_fd_pr__res_xhigh_po_0p35_WX6KG8_0
timestamp 1654038913
transform 1 0 -9 0 1 548
box -37 -532 37 532
use sky130_fd_pr__res_xhigh_po_0p35_WX6KG8  sky130_fd_pr__res_xhigh_po_0p35_WX6KG8_1
timestamp 1654038913
transform 1 0 729 0 1 548
box -37 -532 37 532
<< labels >>
flabel metal1 194 -140 194 -140 0 FreeSans 320 0 0 0 GND
port 3 nsew
flabel metal2 360 -350 360 -350 1 FreeSans 400 0 0 0 ON
port 2 n
flabel metal1 360 1080 360 1080 1 FreeSans 400 0 0 0 V_bias
port 1 n
flabel metal4 -930 -260 -930 -260 1 FreeSans 400 0 0 0 OUT_P
port 4 n
flabel metal4 1690 -270 1690 -270 1 FreeSans 400 0 0 0 OUT_N
port 5 n
<< end >>
