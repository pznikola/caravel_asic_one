magic
tech sky130B
timestamp 1654380865
<< nwell >>
rect -24 2852 121 3273
<< pwell >>
rect -23 2595 121 2829
<< nmos >>
rect 41 2668 56 2818
<< pmos >>
rect 41 2883 56 3183
<< ndiff >>
rect 12 2812 41 2818
rect 12 2674 18 2812
rect 35 2674 41 2812
rect 12 2668 41 2674
rect 56 2812 85 2818
rect 56 2674 62 2812
rect 79 2674 85 2812
rect 56 2668 85 2674
<< pdiff >>
rect 12 3177 41 3183
rect 12 2889 18 3177
rect 35 2889 41 3177
rect 12 2883 41 2889
rect 56 3177 85 3183
rect 56 2889 62 3177
rect 79 2889 85 3177
rect 56 2883 85 2889
<< ndiffc >>
rect 18 2674 35 2812
rect 62 2674 79 2812
<< pdiffc >>
rect 18 2889 35 3177
rect 62 2889 79 3177
<< psubdiff >>
rect 1 2623 100 2624
rect 1 2605 13 2623
rect 31 2605 61 2623
rect 80 2605 100 2623
rect 1 2604 100 2605
<< nsubdiff >>
rect -2 3251 103 3255
rect -2 3232 10 3251
rect 34 3232 67 3251
rect 91 3232 103 3251
rect -2 3228 103 3232
<< psubdiffcont >>
rect 13 2605 31 2623
rect 61 2605 80 2623
<< nsubdiffcont >>
rect 10 3232 34 3251
rect 67 3232 91 3251
<< poly >>
rect 41 3183 56 3196
rect 41 2861 56 2883
rect 110 2861 150 2865
rect 41 2855 150 2861
rect 41 2835 120 2855
rect 140 2835 150 2855
rect 41 2830 150 2835
rect 41 2818 56 2830
rect 110 2825 150 2830
rect 41 2655 56 2668
<< polycont >>
rect 120 2835 140 2855
<< locali >>
rect -23 3251 121 3265
rect -23 3250 10 3251
rect 34 3250 67 3251
rect 91 3250 121 3251
rect -23 3230 -10 3250
rect 50 3232 67 3250
rect 10 3230 30 3232
rect 50 3230 75 3232
rect 95 3230 121 3250
rect -23 3214 121 3230
rect 18 3177 35 3185
rect -75 2865 -45 2870
rect -75 2845 -70 2865
rect -50 2860 -45 2865
rect 18 2861 35 2889
rect 62 3177 79 3214
rect 62 2881 79 2889
rect -24 2860 35 2861
rect -50 2845 35 2860
rect -75 2841 35 2845
rect -75 2840 -15 2841
rect 18 2812 35 2841
rect 110 2855 150 2865
rect 110 2835 120 2855
rect 140 2835 150 2855
rect 110 2825 150 2835
rect 18 2666 35 2674
rect 62 2812 79 2820
rect 62 2634 79 2674
rect -23 2630 121 2634
rect -23 2605 10 2630
rect 35 2623 65 2630
rect 35 2605 61 2623
rect 90 2605 121 2630
rect -23 2595 121 2605
<< viali >>
rect -10 3230 10 3250
rect 30 3232 34 3250
rect 34 3232 50 3250
rect 75 3232 91 3250
rect 91 3232 95 3250
rect 30 3230 50 3232
rect 75 3230 95 3232
rect 18 2889 35 3177
rect -70 2845 -50 2865
rect 62 2889 79 3177
rect 120 2835 140 2855
rect 18 2674 35 2812
rect 62 2674 79 2812
rect 10 2623 35 2630
rect 65 2623 90 2630
rect 10 2605 13 2623
rect 13 2605 31 2623
rect 31 2605 35 2623
rect 65 2605 80 2623
rect 80 2605 90 2623
<< metal1 >>
rect -1710 2635 -705 4880
rect -75 3380 230 4380
rect -75 2865 -45 3380
rect -25 3255 120 3265
rect -25 3225 -15 3255
rect 110 3225 120 3255
rect -25 3215 120 3225
rect 15 3177 38 3183
rect 15 2889 18 3177
rect 35 2889 38 3177
rect 15 2883 38 2889
rect 59 3177 82 3183
rect 59 2889 62 3177
rect 79 2889 82 3177
rect 59 2883 82 2889
rect -75 2845 -70 2865
rect -50 2860 -45 2865
rect 110 2860 150 2865
rect -50 2845 15 2860
rect -75 2840 15 2845
rect -75 2835 -45 2840
rect 110 2830 115 2860
rect 145 2830 150 2860
rect 110 2825 150 2830
rect 15 2812 38 2818
rect 15 2674 18 2812
rect 35 2674 38 2812
rect 15 2668 38 2674
rect 59 2812 82 2818
rect 59 2674 62 2812
rect 79 2674 82 2812
rect 59 2668 82 2674
rect -1710 2630 230 2635
rect -1710 2605 10 2630
rect 35 2605 65 2630
rect 90 2605 230 2630
rect -1710 2595 230 2605
rect -1710 1440 -705 2595
rect -1710 440 230 1440
rect -1710 -60 -705 440
<< via1 >>
rect -15 3250 110 3255
rect -15 3230 -10 3250
rect -10 3230 10 3250
rect 10 3230 30 3250
rect 30 3230 50 3250
rect 50 3230 75 3250
rect 75 3230 95 3250
rect 95 3230 110 3250
rect -15 3225 110 3230
rect 115 2855 145 2860
rect 115 2835 120 2855
rect 120 2835 140 2855
rect 140 2835 145 2855
rect 115 2830 145 2835
<< metal2 >>
rect -3210 3265 -2205 4880
rect -3210 3255 120 3265
rect -3210 3225 -15 3255
rect 110 3225 120 3255
rect -3210 3215 120 3225
rect -3210 -60 -2205 3215
rect 110 2860 230 2865
rect 110 2830 115 2860
rect 145 2830 230 2860
rect 110 2825 230 2830
rect 150 1690 230 2825
<< labels >>
flabel metal1 -75 2890 -75 2890 1 FreeSans 200 0 0 0 OUT
port 2 n
flabel metal2 175 2865 175 2865 1 FreeSans 200 0 0 0 ON
port 1 n
flabel metal2 -2680 4880 -2680 4880 5 FreeSans 1200 0 0 0 VDD
port 3 s
flabel metal1 -1180 4880 -1180 4880 5 FreeSans 1200 0 0 0 GND
port 4 s
<< end >>
